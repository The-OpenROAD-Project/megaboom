// Standard header to adapt well known macros for prints and assertions.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module TLROM(
  input         clock,
                reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
                auto_in_a_bits_param,
  input  [1:0]  auto_in_a_bits_size,
  input  [10:0] auto_in_a_bits_source,
  input  [16:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_a_bits_corrupt,
                auto_in_d_ready,
  output        auto_in_d_valid,
  output [1:0]  auto_in_d_bits_size,
  output [10:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data
);

  reg [63:0] casez_tmp;
  always @(*) begin
    casez (auto_in_a_bits_address[12:3])
      10'b0000000000:
        casez_tmp = 64'h405051300000517;
      10'b0000000001:
        casez_tmp = 64'h301022F330551073;
      10'b0000000010:
        casez_tmp = 64'h12F2934122D293;
      10'b0000000011:
        casez_tmp = 64'h3030107300028463;
      10'b0000000100:
        casez_tmp = 64'h3045107300800513;
      10'b0000000101:
        casez_tmp = 64'h1050007330052073;
      10'b0000000110:
        casez_tmp = 64'hFFDFF06F;
      10'b0000000111:
        casez_tmp = 64'h0;
      10'b0000001000:
        casez_tmp = 64'hF1402573020005B7;
      10'b0000001001:
        casez_tmp = 64'h380006F00050463;
      10'b0000001010:
        casez_tmp = 64'h10069300458613;
      10'b0000001011:
        casez_tmp = 64'h46061300D62023;
      10'b0000001100:
        casez_tmp = 64'hFE069AE3FFC62683;
      10'b0000001101:
        casez_tmp = 64'h2C0006F;
      10'b0000001110:
        casez_tmp = 64'h0;
      10'b0000001111:
        casez_tmp = 64'h0;
      10'b0000010000:
        casez_tmp = 64'h5A283F81FF06F;
      10'b0000010001:
        casez_tmp = 64'h251513FE029EE3;
      10'b0000010010:
        casez_tmp = 64'h5A02300B505B3;
      10'b0000010011:
        casez_tmp = 64'h5350300001537;
      10'b0000010100:
        casez_tmp = 64'hF140257334151073;
      10'b0000010101:
        casez_tmp = 64'h185859300000597;
      10'b0000010110:
        casez_tmp = 64'h3006307308000613;
      10'b0000010111:
        casez_tmp = 64'h1330200073;
      10'b0000011000:
        casez_tmp = 64'hA40F0000EDFE0DD0;
      10'b0000011001:
        casez_tmp = 64'h440D000038000000;
      10'b0000011010:
        casez_tmp = 64'h1100000028000000;
      10'b0000011011:
        casez_tmp = 64'h10000000;
      10'b0000011100:
        casez_tmp = 64'hC0D000060020000;
      10'b0000011101:
        casez_tmp = 64'h0;
      10'b0000011110:
        casez_tmp = 64'h0;
      10'b0000011111:
        casez_tmp = 64'h1000000;
      10'b0000100000:
        casez_tmp = 64'h400000003000000;
      10'b0000100001:
        casez_tmp = 64'h200000000000000;
      10'b0000100010:
        casez_tmp = 64'h400000003000000;
      10'b0000100011:
        casez_tmp = 64'h20000000F000000;
      10'b0000100100:
        casez_tmp = 64'h1500000003000000;
      10'b0000100101:
        casez_tmp = 64'h2D6263751B000000;
      10'b0000100110:
        casez_tmp = 64'h706968632C726162;
      10'b0000100111:
        casez_tmp = 64'h7665642D64726179;
      10'b0000101000:
        casez_tmp = 64'h300000000000000;
      10'b0000101001:
        casez_tmp = 64'h2600000011000000;
      10'b0000101010:
        casez_tmp = 64'h2C7261622D626375;
      10'b0000101011:
        casez_tmp = 64'h6472617970696863;
      10'b0000101100:
        casez_tmp = 64'h100000000000000;
      10'b0000101101:
        casez_tmp = 64'h73657361696C61;
      10'b0000101110:
        casez_tmp = 64'h1500000003000000;
      10'b0000101111:
        casez_tmp = 64'h636F732F2C000000;
      10'b0000110000:
        casez_tmp = 64'h406C61697265732F;
      10'b0000110001:
        casez_tmp = 64'h3030303032303031;
      10'b0000110010:
        casez_tmp = 64'h200000000000000;
      10'b0000110011:
        casez_tmp = 64'h736F686301000000;
      10'b0000110100:
        casez_tmp = 64'h300000000006E65;
      10'b0000110101:
        casez_tmp = 64'h3400000015000000;
      10'b0000110110:
        casez_tmp = 64'h7265732F636F732F;
      10'b0000110111:
        casez_tmp = 64'h32303031406C6169;
      10'b0000111000:
        casez_tmp = 64'h30303030;
      10'b0000111001:
        casez_tmp = 64'h100000002000000;
      10'b0000111010:
        casez_tmp = 64'h73757063;
      10'b0000111011:
        casez_tmp = 64'h400000003000000;
      10'b0000111100:
        casez_tmp = 64'h100000000000000;
      10'b0000111101:
        casez_tmp = 64'h400000003000000;
      10'b0000111110:
        casez_tmp = 64'hF000000;
      10'b0000111111:
        casez_tmp = 64'h400000003000000;
      10'b0001000000:
        casez_tmp = 64'h40420F0040000000;
      10'b0001000001:
        casez_tmp = 64'h4075706301000000;
      10'b0001000010:
        casez_tmp = 64'h300000000000030;
      10'b0001000011:
        casez_tmp = 64'h5300000004000000;
      10'b0001000100:
        casez_tmp = 64'h300000000000000;
      10'b0001000101:
        casez_tmp = 64'h1B00000014000000;
      10'b0001000110:
        casez_tmp = 64'h2C7261622D626375;
      10'b0001000111:
        casez_tmp = 64'h697200306D6F6F62;
      10'b0001001000:
        casez_tmp = 64'h300000000766373;
      10'b0001001001:
        casez_tmp = 64'h6300000004000000;
      10'b0001001010:
        casez_tmp = 64'h300000040000000;
      10'b0001001011:
        casez_tmp = 64'h7600000004000000;
      10'b0001001100:
        casez_tmp = 64'h300000040000000;
      10'b0001001101:
        casez_tmp = 64'h8300000004000000;
      10'b0001001110:
        casez_tmp = 64'h300000000800000;
      10'b0001001111:
        casez_tmp = 64'h9000000004000000;
      10'b0001010000:
        casez_tmp = 64'h300000001000000;
      10'b0001010001:
        casez_tmp = 64'h9B00000004000000;
      10'b0001010010:
        casez_tmp = 64'h300000020000000;
      10'b0001010011:
        casez_tmp = 64'hA600000004000000;
      10'b0001010100:
        casez_tmp = 64'h300000000757063;
      10'b0001010101:
        casez_tmp = 64'hB200000004000000;
      10'b0001010110:
        casez_tmp = 64'h300000000000000;
      10'b0001010111:
        casez_tmp = 64'hD100000004000000;
      10'b0001011000:
        casez_tmp = 64'h300000040000000;
      10'b0001011001:
        casez_tmp = 64'hE400000004000000;
      10'b0001011010:
        casez_tmp = 64'h300000040000000;
      10'b0001011011:
        casez_tmp = 64'hF100000004000000;
      10'b0001011100:
        casez_tmp = 64'h300000000800000;
      10'b0001011101:
        casez_tmp = 64'hFE00000004000000;
      10'b0001011110:
        casez_tmp = 64'h300000001000000;
      10'b0001011111:
        casez_tmp = 64'h901000004000000;
      10'b0001100000:
        casez_tmp = 64'h300000020000000;
      10'b0001100001:
        casez_tmp = 64'h140100000B000000;
      10'b0001100010:
        casez_tmp = 64'h76732C7663736972;
      10'b0001100011:
        casez_tmp = 64'h300000000003933;
      10'b0001100100:
        casez_tmp = 64'h1D01000004000000;
      10'b0001100101:
        casez_tmp = 64'h300000001000000;
      10'b0001100110:
        casez_tmp = 64'h2E01000004000000;
      10'b0001100111:
        casez_tmp = 64'h300000000000000;
      10'b0001101000:
        casez_tmp = 64'h320100001F000000;
      10'b0001101001:
        casez_tmp = 64'h66616D6934367672;
      10'b0001101010:
        casez_tmp = 64'h5F727363697A6364;
      10'b0001101011:
        casez_tmp = 64'h6965636E6566697A;
      10'b0001101100:
        casez_tmp = 64'h6D7068697A5F;
      10'b0001101101:
        casez_tmp = 64'h400000003000000;
      10'b0001101110:
        casez_tmp = 64'h40000003C010000;
      10'b0001101111:
        casez_tmp = 64'h400000003000000;
      10'b0001110000:
        casez_tmp = 64'h800000051010000;
      10'b0001110001:
        casez_tmp = 64'h500000003000000;
      10'b0001110010:
        casez_tmp = 64'h79616B6F62010000;
      10'b0001110011:
        casez_tmp = 64'h300000000000000;
      10'b0001110100:
        casez_tmp = 64'h4000000004000000;
      10'b0001110101:
        casez_tmp = 64'h300000040420F00;
      10'b0001110110:
        casez_tmp = 64'h6901000000000000;
      10'b0001110111:
        casez_tmp = 64'h65746E6901000000;
      10'b0001111000:
        casez_tmp = 64'h6F632D7470757272;
      10'b0001111001:
        casez_tmp = 64'h72656C6C6F72746E;
      10'b0001111010:
        casez_tmp = 64'h300000000000000;
      10'b0001111011:
        casez_tmp = 64'h7301000004000000;
      10'b0001111100:
        casez_tmp = 64'h300000001000000;
      10'b0001111101:
        casez_tmp = 64'h1B0000000F000000;
      10'b0001111110:
        casez_tmp = 64'h70632C7663736972;
      10'b0001111111:
        casez_tmp = 64'h63746E692D75;
      10'b0010000000:
        casez_tmp = 64'h3000000;
      10'b0010000001:
        casez_tmp = 64'h300000084010000;
      10'b0010000010:
        casez_tmp = 64'h9901000004000000;
      10'b0010000011:
        casez_tmp = 64'h200000004000000;
      10'b0010000100:
        casez_tmp = 64'h200000002000000;
      10'b0010000101:
        casez_tmp = 64'h6669746801000000;
      10'b0010000110:
        casez_tmp = 64'h300000000000000;
      10'b0010000111:
        casez_tmp = 64'h1B0000000A000000;
      10'b0010001000:
        casez_tmp = 64'h666974682C626375;
      10'b0010001001:
        casez_tmp = 64'h200000000000030;
      10'b0010001010:
        casez_tmp = 64'h6F6D656D01000000;
      10'b0010001011:
        casez_tmp = 64'h3030303038407972;
      10'b0010001100:
        casez_tmp = 64'h300000000003030;
      10'b0010001101:
        casez_tmp = 64'hA600000007000000;
      10'b0010001110:
        casez_tmp = 64'h79726F6D656D;
      10'b0010001111:
        casez_tmp = 64'h1000000003000000;
      10'b0010010000:
        casez_tmp = 64'h2E010000;
      10'b0010010001:
        casez_tmp = 64'h8;
      10'b0010010010:
        casez_tmp = 64'h300000000000100;
      10'b0010010011:
        casez_tmp = 64'h9901000004000000;
      10'b0010010100:
        casez_tmp = 64'h200000003000000;
      10'b0010010101:
        casez_tmp = 64'h6F6D656D01000000;
      10'b0010010110:
        casez_tmp = 64'h3030303038407972;
      10'b0010010111:
        casez_tmp = 64'h300000000303030;
      10'b0010011000:
        casez_tmp = 64'hA600000007000000;
      10'b0010011001:
        casez_tmp = 64'h79726F6D656D;
      10'b0010011010:
        casez_tmp = 64'h1000000003000000;
      10'b0010011011:
        casez_tmp = 64'h2E010000;
      10'b0010011100:
        casez_tmp = 64'h100000000000080;
      10'b0010011101:
        casez_tmp = 64'h300000000000000;
      10'b0010011110:
        casez_tmp = 64'h9901000004000000;
      10'b0010011111:
        casez_tmp = 64'h200000002000000;
      10'b0010100000:
        casez_tmp = 64'h636F7301000000;
      10'b0010100001:
        casez_tmp = 64'h400000003000000;
      10'b0010100010:
        casez_tmp = 64'h200000000000000;
      10'b0010100011:
        casez_tmp = 64'h400000003000000;
      10'b0010100100:
        casez_tmp = 64'h20000000F000000;
      10'b0010100101:
        casez_tmp = 64'h2000000003000000;
      10'b0010100110:
        casez_tmp = 64'h2D6263751B000000;
      10'b0010100111:
        casez_tmp = 64'h706968632C726162;
      10'b0010101000:
        casez_tmp = 64'h636F732D64726179;
      10'b0010101001:
        casez_tmp = 64'h2D656C706D697300;
      10'b0010101010:
        casez_tmp = 64'h300000000737562;
      10'b0010101011:
        casez_tmp = 64'hA101000000000000;
      10'b0010101100:
        casez_tmp = 64'h746F6F6201000000;
      10'b0010101101:
        casez_tmp = 64'h737365726464612D;
      10'b0010101110:
        casez_tmp = 64'h303031406765722D;
      10'b0010101111:
        casez_tmp = 64'h300000000000030;
      10'b0010110000:
        casez_tmp = 64'h2E01000010000000;
      10'b0010110001:
        casez_tmp = 64'h10000000000000;
      10'b0010110010:
        casez_tmp = 64'h10000000000000;
      10'b0010110011:
        casez_tmp = 64'h800000003000000;
      10'b0010110100:
        casez_tmp = 64'h746E6F63A8010000;
      10'b0010110101:
        casez_tmp = 64'h2000000006C6F72;
      10'b0010110110:
        casez_tmp = 64'h6863616301000000;
      10'b0010110111:
        casez_tmp = 64'h6F72746E6F632D65;
      10'b0010111000:
        casez_tmp = 64'h3130324072656C6C;
      10'b0010111001:
        casez_tmp = 64'h30303030;
      10'b0010111010:
        casez_tmp = 64'h400000003000000;
      10'b0010111011:
        casez_tmp = 64'h4000000065000000;
      10'b0010111100:
        casez_tmp = 64'h400000003000000;
      10'b0010111101:
        casez_tmp = 64'h2000000B2010000;
      10'b0010111110:
        casez_tmp = 64'h400000003000000;
      10'b0010111111:
        casez_tmp = 64'h4000078000000;
      10'b0011000000:
        casez_tmp = 64'h400000003000000;
      10'b0011000001:
        casez_tmp = 64'h80085000000;
      10'b0011000010:
        casez_tmp = 64'h3000000;
      10'b0011000011:
        casez_tmp = 64'h3000000BE010000;
      10'b0011000100:
        casez_tmp = 64'h1B0000001D000000;
      10'b0011000101:
        casez_tmp = 64'h692C657669666973;
      10'b0011000110:
        casez_tmp = 64'h65766973756C636E;
      10'b0011000111:
        casez_tmp = 64'h6300306568636163;
      10'b0011001000:
        casez_tmp = 64'h65686361;
      10'b0011001001:
        casez_tmp = 64'h800000003000000;
      10'b0011001010:
        casez_tmp = 64'h20000001D010000;
      10'b0011001011:
        casez_tmp = 64'h300000003000000;
      10'b0011001100:
        casez_tmp = 64'h2E01000010000000;
      10'b0011001101:
        casez_tmp = 64'h10200000000;
      10'b0011001110:
        casez_tmp = 64'h10000000000000;
      10'b0011001111:
        casez_tmp = 64'h800000003000000;
      10'b0011010000:
        casez_tmp = 64'h746E6F63A8010000;
      10'b0011010001:
        casez_tmp = 64'h3000000006C6F72;
      10'b0011010010:
        casez_tmp = 64'hCC01000004000000;
      10'b0011010011:
        casez_tmp = 64'h300000007000000;
      10'b0011010100:
        casez_tmp = 64'h9901000004000000;
      10'b0011010101:
        casez_tmp = 64'h200000001000000;
      10'b0011010110:
        casez_tmp = 64'h6E696C6301000000;
      10'b0011010111:
        casez_tmp = 64'h3030303030324074;
      10'b0011011000:
        casez_tmp = 64'h300000000000030;
      10'b0011011001:
        casez_tmp = 64'h1B0000000D000000;
      10'b0011011010:
        casez_tmp = 64'h6C632C7663736972;
      10'b0011011011:
        casez_tmp = 64'h30746E69;
      10'b0011011100:
        casez_tmp = 64'h1000000003000000;
      10'b0011011101:
        casez_tmp = 64'h4000000DE010000;
      10'b0011011110:
        casez_tmp = 64'h400000003000000;
      10'b0011011111:
        casez_tmp = 64'h300000007000000;
      10'b0011100000:
        casez_tmp = 64'h2E01000010000000;
      10'b0011100001:
        casez_tmp = 64'h200000000;
      10'b0011100010:
        casez_tmp = 64'h10000000000;
      10'b0011100011:
        casez_tmp = 64'h800000003000000;
      10'b0011100100:
        casez_tmp = 64'h746E6F63A8010000;
      10'b0011100101:
        casez_tmp = 64'h2000000006C6F72;
      10'b0011100110:
        casez_tmp = 64'h636F6C6301000000;
      10'b0011100111:
        casez_tmp = 64'h4072657461672D6B;
      10'b0011101000:
        casez_tmp = 64'h303030303031;
      10'b0011101001:
        casez_tmp = 64'h1000000003000000;
      10'b0011101010:
        casez_tmp = 64'h2E010000;
      10'b0011101011:
        casez_tmp = 64'h1000;
      10'b0011101100:
        casez_tmp = 64'h300000000100000;
      10'b0011101101:
        casez_tmp = 64'hA801000008000000;
      10'b0011101110:
        casez_tmp = 64'h6C6F72746E6F63;
      10'b0011101111:
        casez_tmp = 64'h100000002000000;
      10'b0011110000:
        casez_tmp = 64'h6F632D6775626564;
      10'b0011110001:
        casez_tmp = 64'h72656C6C6F72746E;
      10'b0011110010:
        casez_tmp = 64'h300000000003040;
      10'b0011110011:
        casez_tmp = 64'h1B00000021000000;
      10'b0011110100:
        casez_tmp = 64'h642C657669666973;
      10'b0011110101:
        casez_tmp = 64'h3331302D67756265;
      10'b0011110110:
        casez_tmp = 64'h642C766373697200;
      10'b0011110111:
        casez_tmp = 64'h3331302D67756265;
      10'b0011111000:
        casez_tmp = 64'h300000000000000;
      10'b0011111001:
        casez_tmp = 64'hF201000005000000;
      10'b0011111010:
        casez_tmp = 64'h6761746A;
      10'b0011111011:
        casez_tmp = 64'h800000003000000;
      10'b0011111100:
        casez_tmp = 64'h4000000DE010000;
      10'b0011111101:
        casez_tmp = 64'h3000000FFFF0000;
      10'b0011111110:
        casez_tmp = 64'h2E01000010000000;
      10'b0011111111:
        casez_tmp = 64'h0;
      10'b0100000000:
        casez_tmp = 64'h10000000000000;
      10'b0100000001:
        casez_tmp = 64'h800000003000000;
      10'b0100000010:
        casez_tmp = 64'h746E6F63A8010000;
      10'b0100000011:
        casez_tmp = 64'h2000000006C6F72;
      10'b0100000100:
        casez_tmp = 64'h6F72726501000000;
      10'b0100000101:
        casez_tmp = 64'h6563697665642D72;
      10'b0100000110:
        casez_tmp = 64'h3030303340;
      10'b0100000111:
        casez_tmp = 64'hE00000003000000;
      10'b0100001000:
        casez_tmp = 64'h696669731B000000;
      10'b0100001001:
        casez_tmp = 64'h726F7272652C6576;
      10'b0100001010:
        casez_tmp = 64'h300000000000030;
      10'b0100001011:
        casez_tmp = 64'h2E01000010000000;
      10'b0100001100:
        casez_tmp = 64'h30000000000000;
      10'b0100001101:
        casez_tmp = 64'h10000000000000;
      10'b0100001110:
        casez_tmp = 64'h100000002000000;
      10'b0100001111:
        casez_tmp = 64'h7075727265746E69;
      10'b0100010000:
        casez_tmp = 64'h6F72746E6F632D74;
      10'b0100010001:
        casez_tmp = 64'h3030634072656C6C;
      10'b0100010010:
        casez_tmp = 64'h30303030;
      10'b0100010011:
        casez_tmp = 64'h400000003000000;
      10'b0100010100:
        casez_tmp = 64'h100000073010000;
      10'b0100010101:
        casez_tmp = 64'hC00000003000000;
      10'b0100010110:
        casez_tmp = 64'h637369721B000000;
      10'b0100010111:
        casez_tmp = 64'h3063696C702C76;
      10'b0100011000:
        casez_tmp = 64'h3000000;
      10'b0100011001:
        casez_tmp = 64'h300000084010000;
      10'b0100011010:
        casez_tmp = 64'hDE01000010000000;
      10'b0100011011:
        casez_tmp = 64'hB00000004000000;
      10'b0100011100:
        casez_tmp = 64'h900000004000000;
      10'b0100011101:
        casez_tmp = 64'h1000000003000000;
      10'b0100011110:
        casez_tmp = 64'h2E010000;
      10'b0100011111:
        casez_tmp = 64'hC;
      10'b0100100000:
        casez_tmp = 64'h300000000000004;
      10'b0100100001:
        casez_tmp = 64'hA801000008000000;
      10'b0100100010:
        casez_tmp = 64'h6C6F72746E6F63;
      10'b0100100011:
        casez_tmp = 64'h400000003000000;
      10'b0100100100:
        casez_tmp = 64'h1000000FF010000;
      10'b0100100101:
        casez_tmp = 64'h400000003000000;
      10'b0100100110:
        casez_tmp = 64'h100000012020000;
      10'b0100100111:
        casez_tmp = 64'h400000003000000;
      10'b0100101000:
        casez_tmp = 64'h600000099010000;
      10'b0100101001:
        casez_tmp = 64'h100000002000000;
      10'b0100101010:
        casez_tmp = 64'h30303031406D6F72;
      10'b0100101011:
        casez_tmp = 64'h300000000000030;
      10'b0100101100:
        casez_tmp = 64'h1B0000000C000000;
      10'b0100101101:
        casez_tmp = 64'h722C657669666973;
      10'b0100101110:
        casez_tmp = 64'h300000000306D6F;
      10'b0100101111:
        casez_tmp = 64'h2E01000010000000;
      10'b0100110000:
        casez_tmp = 64'h10000000000;
      10'b0100110001:
        casez_tmp = 64'h10000000000;
      10'b0100110010:
        casez_tmp = 64'h400000003000000;
      10'b0100110011:
        casez_tmp = 64'h6D656DA8010000;
      10'b0100110100:
        casez_tmp = 64'h100000002000000;
      10'b0100110101:
        casez_tmp = 64'h31406C6169726573;
      10'b0100110110:
        casez_tmp = 64'h30303030323030;
      10'b0100110111:
        casez_tmp = 64'h400000003000000;
      10'b0100111000:
        casez_tmp = 64'h50000001D020000;
      10'b0100111001:
        casez_tmp = 64'hD00000003000000;
      10'b0100111010:
        casez_tmp = 64'h696669731B000000;
      10'b0100111011:
        casez_tmp = 64'h30747261752C6576;
      10'b0100111100:
        casez_tmp = 64'h300000000000000;
      10'b0100111101:
        casez_tmp = 64'h2402000004000000;
      10'b0100111110:
        casez_tmp = 64'h300000006000000;
      10'b0100111111:
        casez_tmp = 64'h3502000004000000;
      10'b0101000000:
        casez_tmp = 64'h300000001000000;
      10'b0101000001:
        casez_tmp = 64'h2E01000010000000;
      10'b0101000010:
        casez_tmp = 64'h21000000000;
      10'b0101000011:
        casez_tmp = 64'h10000000000000;
      10'b0101000100:
        casez_tmp = 64'h800000003000000;
      10'b0101000101:
        casez_tmp = 64'h746E6F63A8010000;
      10'b0101000110:
        casez_tmp = 64'h2000000006C6F72;
      10'b0101000111:
        casez_tmp = 64'h7362757301000000;
      10'b0101001000:
        casez_tmp = 64'h62635F6D65747379;
      10'b0101001001:
        casez_tmp = 64'h6B636F6C635F7375;
      10'b0101001010:
        casez_tmp = 64'h300000000000000;
      10'b0101001011:
        casez_tmp = 64'h4002000004000000;
      10'b0101001100:
        casez_tmp = 64'h300000000000000;
      10'b0101001101:
        casez_tmp = 64'h5300000004000000;
      10'b0101001110:
        casez_tmp = 64'h30000000065CD1D;
      10'b0101001111:
        casez_tmp = 64'h4D02000015000000;
      10'b0101010000:
        casez_tmp = 64'h6574737973627573;
      10'b0101010001:
        casez_tmp = 64'h635F737562635F6D;
      10'b0101010010:
        casez_tmp = 64'h6B636F6C;
      10'b0101010011:
        casez_tmp = 64'hC00000003000000;
      10'b0101010100:
        casez_tmp = 64'h657869661B000000;
      10'b0101010101:
        casez_tmp = 64'h6B636F6C632D64;
      10'b0101010110:
        casez_tmp = 64'h100000002000000;
      10'b0101010111:
        casez_tmp = 64'h6574737973627573;
      10'b0101011000:
        casez_tmp = 64'h635F737562665F6D;
      10'b0101011001:
        casez_tmp = 64'h6B636F6C;
      10'b0101011010:
        casez_tmp = 64'h400000003000000;
      10'b0101011011:
        casez_tmp = 64'h40020000;
      10'b0101011100:
        casez_tmp = 64'h400000003000000;
      10'b0101011101:
        casez_tmp = 64'h65CD1D53000000;
      10'b0101011110:
        casez_tmp = 64'h1500000003000000;
      10'b0101011111:
        casez_tmp = 64'h736275734D020000;
      10'b0101100000:
        casez_tmp = 64'h62665F6D65747379;
      10'b0101100001:
        casez_tmp = 64'h6B636F6C635F7375;
      10'b0101100010:
        casez_tmp = 64'h300000000000000;
      10'b0101100011:
        casez_tmp = 64'h1B0000000C000000;
      10'b0101100100:
        casez_tmp = 64'h6C632D6465786966;
      10'b0101100101:
        casez_tmp = 64'h2000000006B636F;
      10'b0101100110:
        casez_tmp = 64'h7362757301000000;
      10'b0101100111:
        casez_tmp = 64'h326C5F6D65747379;
      10'b0101101000:
        casez_tmp = 64'h6B636F6C635F;
      10'b0101101001:
        casez_tmp = 64'h400000003000000;
      10'b0101101010:
        casez_tmp = 64'h40020000;
      10'b0101101011:
        casez_tmp = 64'h400000003000000;
      10'b0101101100:
        casez_tmp = 64'h65CD1D53000000;
      10'b0101101101:
        casez_tmp = 64'h1300000003000000;
      10'b0101101110:
        casez_tmp = 64'h736275734D020000;
      10'b0101101111:
        casez_tmp = 64'h326C5F6D65747379;
      10'b0101110000:
        casez_tmp = 64'h6B636F6C635F;
      10'b0101110001:
        casez_tmp = 64'hC00000003000000;
      10'b0101110010:
        casez_tmp = 64'h657869661B000000;
      10'b0101110011:
        casez_tmp = 64'h6B636F6C632D64;
      10'b0101110100:
        casez_tmp = 64'h100000002000000;
      10'b0101110101:
        casez_tmp = 64'h6574737973627573;
      10'b0101110110:
        casez_tmp = 64'h635F7375626D5F6D;
      10'b0101110111:
        casez_tmp = 64'h6B636F6C;
      10'b0101111000:
        casez_tmp = 64'h400000003000000;
      10'b0101111001:
        casez_tmp = 64'h40020000;
      10'b0101111010:
        casez_tmp = 64'h400000003000000;
      10'b0101111011:
        casez_tmp = 64'h65CD1D53000000;
      10'b0101111100:
        casez_tmp = 64'h1500000003000000;
      10'b0101111101:
        casez_tmp = 64'h736275734D020000;
      10'b0101111110:
        casez_tmp = 64'h626D5F6D65747379;
      10'b0101111111:
        casez_tmp = 64'h6B636F6C635F7375;
      10'b0110000000:
        casez_tmp = 64'h300000000000000;
      10'b0110000001:
        casez_tmp = 64'h1B0000000C000000;
      10'b0110000010:
        casez_tmp = 64'h6C632D6465786966;
      10'b0110000011:
        casez_tmp = 64'h2000000006B636F;
      10'b0110000100:
        casez_tmp = 64'h7362757301000000;
      10'b0110000101:
        casez_tmp = 64'h626F5F6D65747379;
      10'b0110000110:
        casez_tmp = 64'h6B636F6C635F7375;
      10'b0110000111:
        casez_tmp = 64'h300000000000000;
      10'b0110001000:
        casez_tmp = 64'h4002000004000000;
      10'b0110001001:
        casez_tmp = 64'h300000000000000;
      10'b0110001010:
        casez_tmp = 64'h5300000004000000;
      10'b0110001011:
        casez_tmp = 64'h30000000065CD1D;
      10'b0110001100:
        casez_tmp = 64'h4D02000015000000;
      10'b0110001101:
        casez_tmp = 64'h6574737973627573;
      10'b0110001110:
        casez_tmp = 64'h635F7375626F5F6D;
      10'b0110001111:
        casez_tmp = 64'h6B636F6C;
      10'b0110010000:
        casez_tmp = 64'hC00000003000000;
      10'b0110010001:
        casez_tmp = 64'h657869661B000000;
      10'b0110010010:
        casez_tmp = 64'h6B636F6C632D64;
      10'b0110010011:
        casez_tmp = 64'h100000002000000;
      10'b0110010100:
        casez_tmp = 64'h6574737973627573;
      10'b0110010101:
        casez_tmp = 64'h635F737562705F6D;
      10'b0110010110:
        casez_tmp = 64'h6B636F6C;
      10'b0110010111:
        casez_tmp = 64'h400000003000000;
      10'b0110011000:
        casez_tmp = 64'h40020000;
      10'b0110011001:
        casez_tmp = 64'h400000003000000;
      10'b0110011010:
        casez_tmp = 64'h65CD1D53000000;
      10'b0110011011:
        casez_tmp = 64'h1500000003000000;
      10'b0110011100:
        casez_tmp = 64'h736275734D020000;
      10'b0110011101:
        casez_tmp = 64'h62705F6D65747379;
      10'b0110011110:
        casez_tmp = 64'h6B636F6C635F7375;
      10'b0110011111:
        casez_tmp = 64'h300000000000000;
      10'b0110100000:
        casez_tmp = 64'h1B0000000C000000;
      10'b0110100001:
        casez_tmp = 64'h6C632D6465786966;
      10'b0110100010:
        casez_tmp = 64'h3000000006B636F;
      10'b0110100011:
        casez_tmp = 64'h9901000004000000;
      10'b0110100100:
        casez_tmp = 64'h200000005000000;
      10'b0110100101:
        casez_tmp = 64'h7362757301000000;
      10'b0110100110:
        casez_tmp = 64'h62735F6D65747379;
      10'b0110100111:
        casez_tmp = 64'h6B636F6C635F7375;
      10'b0110101000:
        casez_tmp = 64'h300000000000000;
      10'b0110101001:
        casez_tmp = 64'h4002000004000000;
      10'b0110101010:
        casez_tmp = 64'h300000000000000;
      10'b0110101011:
        casez_tmp = 64'h5300000004000000;
      10'b0110101100:
        casez_tmp = 64'h30000000065CD1D;
      10'b0110101101:
        casez_tmp = 64'h4D02000015000000;
      10'b0110101110:
        casez_tmp = 64'h6574737973627573;
      10'b0110101111:
        casez_tmp = 64'h635F737562735F6D;
      10'b0110110000:
        casez_tmp = 64'h6B636F6C;
      10'b0110110001:
        casez_tmp = 64'hC00000003000000;
      10'b0110110010:
        casez_tmp = 64'h657869661B000000;
      10'b0110110011:
        casez_tmp = 64'h6B636F6C632D64;
      10'b0110110100:
        casez_tmp = 64'h100000002000000;
      10'b0110110101:
        casez_tmp = 64'h7365722D656C6974;
      10'b0110110110:
        casez_tmp = 64'h65747465732D7465;
      10'b0110110111:
        casez_tmp = 64'h3030303031314072;
      10'b0110111000:
        casez_tmp = 64'h300000000000000;
      10'b0110111001:
        casez_tmp = 64'h2E01000010000000;
      10'b0110111010:
        casez_tmp = 64'h110000000000;
      10'b0110111011:
        casez_tmp = 64'h10000000000000;
      10'b0110111100:
        casez_tmp = 64'h800000003000000;
      10'b0110111101:
        casez_tmp = 64'h746E6F63A8010000;
      10'b0110111110:
        casez_tmp = 64'h2000000006C6F72;
      10'b0110111111:
        casez_tmp = 64'h200000002000000;
      10'b0111000000:
        casez_tmp = 64'h6464612309000000;
      10'b0111000001:
        casez_tmp = 64'h6C65632D73736572;
      10'b0111000010:
        casez_tmp = 64'h657A69732300736C;
      10'b0111000011:
        casez_tmp = 64'h6300736C6C65632D;
      10'b0111000100:
        casez_tmp = 64'h6C62697461706D6F;
      10'b0111000101:
        casez_tmp = 64'h6C65646F6D0065;
      10'b0111000110:
        casez_tmp = 64'h306C6169726573;
      10'b0111000111:
        casez_tmp = 64'h702D74756F647473;
      10'b0111001000:
        casez_tmp = 64'h656D697400687461;
      10'b0111001001:
        casez_tmp = 64'h6572662D65736162;
      10'b0111001010:
        casez_tmp = 64'h630079636E657571;
      10'b0111001011:
        casez_tmp = 64'h6572662D6B636F6C;
      10'b0111001100:
        casez_tmp = 64'h640079636E657571;
      10'b0111001101:
        casez_tmp = 64'h622D65686361632D;
      10'b0111001110:
        casez_tmp = 64'h7A69732D6B636F6C;
      10'b0111001111:
        casez_tmp = 64'h686361632D640065;
      10'b0111010000:
        casez_tmp = 64'h6400737465732D65;
      10'b0111010001:
        casez_tmp = 64'h732D65686361632D;
      10'b0111010010:
        casez_tmp = 64'h6C742D6400657A69;
      10'b0111010011:
        casez_tmp = 64'h6400737465732D62;
      10'b0111010100:
        casez_tmp = 64'h7A69732D626C742D;
      10'b0111010101:
        casez_tmp = 64'h6563697665640065;
      10'b0111010110:
        casez_tmp = 64'h616800657079745F;
      10'b0111010111:
        casez_tmp = 64'h652D657261776472;
      10'b0111011000:
        casez_tmp = 64'h616572622D636578;
      10'b0111011001:
        casez_tmp = 64'h632D746E696F706B;
      10'b0111011010:
        casez_tmp = 64'h632D6900746E756F;
      10'b0111011011:
        casez_tmp = 64'h6F6C622D65686361;
      10'b0111011100:
        casez_tmp = 64'h657A69732D6B63;
      10'b0111011101:
        casez_tmp = 64'h2D65686361632D69;
      10'b0111011110:
        casez_tmp = 64'h632D690073746573;
      10'b0111011111:
        casez_tmp = 64'h7A69732D65686361;
      10'b0111100000:
        casez_tmp = 64'h2D626C742D690065;
      10'b0111100001:
        casez_tmp = 64'h742D690073746573;
      10'b0111100010:
        casez_tmp = 64'h657A69732D626C;
      10'b0111100011:
        casez_tmp = 64'h657079742D756D6D;
      10'b0111100100:
        casez_tmp = 64'h656C2D7478656E00;
      10'b0111100101:
        casez_tmp = 64'h686361632D6C6576;
      10'b0111100110:
        casez_tmp = 64'h6972006765720065;
      10'b0111100111:
        casez_tmp = 64'h6173692C766373;
      10'b0111101000:
        casez_tmp = 64'h6D702C7663736972;
      10'b0111101001:
        casez_tmp = 64'h616C756E61726770;
      10'b0111101010:
        casez_tmp = 64'h7369720079746972;
      10'b0111101011:
        casez_tmp = 64'h6572706D702C7663;
      10'b0111101100:
        casez_tmp = 64'h747300736E6F6967;
      10'b0111101101:
        casez_tmp = 64'h626C740073757461;
      10'b0111101110:
        casez_tmp = 64'h230074696C70732D;
      10'b0111101111:
        casez_tmp = 64'h7075727265746E69;
      10'b0111110000:
        casez_tmp = 64'h736C6C65632D74;
      10'b0111110001:
        casez_tmp = 64'h7075727265746E69;
      10'b0111110010:
        casez_tmp = 64'h6F72746E6F632D74;
      10'b0111110011:
        casez_tmp = 64'h6168700072656C6C;
      10'b0111110100:
        casez_tmp = 64'h6E617200656C646E;
      10'b0111110101:
        casez_tmp = 64'h2D67657200736567;
      10'b0111110110:
        casez_tmp = 64'h61630073656D616E;
      10'b0111110111:
        casez_tmp = 64'h6576656C2D656863;
      10'b0111111000:
        casez_tmp = 64'h2D6568636163006C;
      10'b0111111001:
        casez_tmp = 64'h64656966696E75;
      10'b0111111010:
        casez_tmp = 64'h6D2C657669666973;
      10'b0111111011:
        casez_tmp = 64'h6E756F632D726873;
      10'b0111111100:
        casez_tmp = 64'h727265746E690074;
      10'b0111111101:
        casez_tmp = 64'h7478652D73747075;
      10'b0111111110:
        casez_tmp = 64'h6564006465646E65;
      10'b0111111111:
        casez_tmp = 64'h617474612D677562;
      10'b1000000000:
        casez_tmp = 64'h7663736972006863;
      10'b1000000001:
        casez_tmp = 64'h6972702D78616D2C;
      10'b1000000010:
        casez_tmp = 64'h697200797469726F;
      10'b1000000011:
        casez_tmp = 64'h7665646E2C766373;
      10'b1000000100:
        casez_tmp = 64'h736B636F6C6300;
      10'b1000000101:
        casez_tmp = 64'h7075727265746E69;
      10'b1000000110:
        casez_tmp = 64'h746E657261702D74;
      10'b1000000111:
        casez_tmp = 64'h75727265746E6900;
      10'b1000001000:
        casez_tmp = 64'h6F6C632300737470;
      10'b1000001001:
        casez_tmp = 64'h736C6C65632D6B63;
      10'b1000001010:
        casez_tmp = 64'h6F2D6B636F6C6300;
      10'b1000001011:
        casez_tmp = 64'h616E2D7475707475;
      10'b1000001100:
        casez_tmp = 64'h73656D;
      10'b1000001101:
        casez_tmp = 64'h0;
      10'b1000001110:
        casez_tmp = 64'h0;
      10'b1000001111:
        casez_tmp = 64'h0;
      10'b1000010000:
        casez_tmp = 64'h0;
      10'b1000010001:
        casez_tmp = 64'h0;
      10'b1000010010:
        casez_tmp = 64'h0;
      10'b1000010011:
        casez_tmp = 64'h0;
      10'b1000010100:
        casez_tmp = 64'h0;
      10'b1000010101:
        casez_tmp = 64'h0;
      10'b1000010110:
        casez_tmp = 64'h0;
      10'b1000010111:
        casez_tmp = 64'h0;
      10'b1000011000:
        casez_tmp = 64'h0;
      10'b1000011001:
        casez_tmp = 64'h0;
      10'b1000011010:
        casez_tmp = 64'h0;
      10'b1000011011:
        casez_tmp = 64'h0;
      10'b1000011100:
        casez_tmp = 64'h0;
      10'b1000011101:
        casez_tmp = 64'h0;
      10'b1000011110:
        casez_tmp = 64'h0;
      10'b1000011111:
        casez_tmp = 64'h0;
      10'b1000100000:
        casez_tmp = 64'h0;
      10'b1000100001:
        casez_tmp = 64'h0;
      10'b1000100010:
        casez_tmp = 64'h0;
      10'b1000100011:
        casez_tmp = 64'h0;
      10'b1000100100:
        casez_tmp = 64'h0;
      10'b1000100101:
        casez_tmp = 64'h0;
      10'b1000100110:
        casez_tmp = 64'h0;
      10'b1000100111:
        casez_tmp = 64'h0;
      10'b1000101000:
        casez_tmp = 64'h0;
      10'b1000101001:
        casez_tmp = 64'h0;
      10'b1000101010:
        casez_tmp = 64'h0;
      10'b1000101011:
        casez_tmp = 64'h0;
      10'b1000101100:
        casez_tmp = 64'h0;
      10'b1000101101:
        casez_tmp = 64'h0;
      10'b1000101110:
        casez_tmp = 64'h0;
      10'b1000101111:
        casez_tmp = 64'h0;
      10'b1000110000:
        casez_tmp = 64'h0;
      10'b1000110001:
        casez_tmp = 64'h0;
      10'b1000110010:
        casez_tmp = 64'h0;
      10'b1000110011:
        casez_tmp = 64'h0;
      10'b1000110100:
        casez_tmp = 64'h0;
      10'b1000110101:
        casez_tmp = 64'h0;
      10'b1000110110:
        casez_tmp = 64'h0;
      10'b1000110111:
        casez_tmp = 64'h0;
      10'b1000111000:
        casez_tmp = 64'h0;
      10'b1000111001:
        casez_tmp = 64'h0;
      10'b1000111010:
        casez_tmp = 64'h0;
      10'b1000111011:
        casez_tmp = 64'h0;
      10'b1000111100:
        casez_tmp = 64'h0;
      10'b1000111101:
        casez_tmp = 64'h0;
      10'b1000111110:
        casez_tmp = 64'h0;
      10'b1000111111:
        casez_tmp = 64'h0;
      10'b1001000000:
        casez_tmp = 64'h0;
      10'b1001000001:
        casez_tmp = 64'h0;
      10'b1001000010:
        casez_tmp = 64'h0;
      10'b1001000011:
        casez_tmp = 64'h0;
      10'b1001000100:
        casez_tmp = 64'h0;
      10'b1001000101:
        casez_tmp = 64'h0;
      10'b1001000110:
        casez_tmp = 64'h0;
      10'b1001000111:
        casez_tmp = 64'h0;
      10'b1001001000:
        casez_tmp = 64'h0;
      10'b1001001001:
        casez_tmp = 64'h0;
      10'b1001001010:
        casez_tmp = 64'h0;
      10'b1001001011:
        casez_tmp = 64'h0;
      10'b1001001100:
        casez_tmp = 64'h0;
      10'b1001001101:
        casez_tmp = 64'h0;
      10'b1001001110:
        casez_tmp = 64'h0;
      10'b1001001111:
        casez_tmp = 64'h0;
      10'b1001010000:
        casez_tmp = 64'h0;
      10'b1001010001:
        casez_tmp = 64'h0;
      10'b1001010010:
        casez_tmp = 64'h0;
      10'b1001010011:
        casez_tmp = 64'h0;
      10'b1001010100:
        casez_tmp = 64'h0;
      10'b1001010101:
        casez_tmp = 64'h0;
      10'b1001010110:
        casez_tmp = 64'h0;
      10'b1001010111:
        casez_tmp = 64'h0;
      10'b1001011000:
        casez_tmp = 64'h0;
      10'b1001011001:
        casez_tmp = 64'h0;
      10'b1001011010:
        casez_tmp = 64'h0;
      10'b1001011011:
        casez_tmp = 64'h0;
      10'b1001011100:
        casez_tmp = 64'h0;
      10'b1001011101:
        casez_tmp = 64'h0;
      10'b1001011110:
        casez_tmp = 64'h0;
      10'b1001011111:
        casez_tmp = 64'h0;
      10'b1001100000:
        casez_tmp = 64'h0;
      10'b1001100001:
        casez_tmp = 64'h0;
      10'b1001100010:
        casez_tmp = 64'h0;
      10'b1001100011:
        casez_tmp = 64'h0;
      10'b1001100100:
        casez_tmp = 64'h0;
      10'b1001100101:
        casez_tmp = 64'h0;
      10'b1001100110:
        casez_tmp = 64'h0;
      10'b1001100111:
        casez_tmp = 64'h0;
      10'b1001101000:
        casez_tmp = 64'h0;
      10'b1001101001:
        casez_tmp = 64'h0;
      10'b1001101010:
        casez_tmp = 64'h0;
      10'b1001101011:
        casez_tmp = 64'h0;
      10'b1001101100:
        casez_tmp = 64'h0;
      10'b1001101101:
        casez_tmp = 64'h0;
      10'b1001101110:
        casez_tmp = 64'h0;
      10'b1001101111:
        casez_tmp = 64'h0;
      10'b1001110000:
        casez_tmp = 64'h0;
      10'b1001110001:
        casez_tmp = 64'h0;
      10'b1001110010:
        casez_tmp = 64'h0;
      10'b1001110011:
        casez_tmp = 64'h0;
      10'b1001110100:
        casez_tmp = 64'h0;
      10'b1001110101:
        casez_tmp = 64'h0;
      10'b1001110110:
        casez_tmp = 64'h0;
      10'b1001110111:
        casez_tmp = 64'h0;
      10'b1001111000:
        casez_tmp = 64'h0;
      10'b1001111001:
        casez_tmp = 64'h0;
      10'b1001111010:
        casez_tmp = 64'h0;
      10'b1001111011:
        casez_tmp = 64'h0;
      10'b1001111100:
        casez_tmp = 64'h0;
      10'b1001111101:
        casez_tmp = 64'h0;
      10'b1001111110:
        casez_tmp = 64'h0;
      10'b1001111111:
        casez_tmp = 64'h0;
      10'b1010000000:
        casez_tmp = 64'h0;
      10'b1010000001:
        casez_tmp = 64'h0;
      10'b1010000010:
        casez_tmp = 64'h0;
      10'b1010000011:
        casez_tmp = 64'h0;
      10'b1010000100:
        casez_tmp = 64'h0;
      10'b1010000101:
        casez_tmp = 64'h0;
      10'b1010000110:
        casez_tmp = 64'h0;
      10'b1010000111:
        casez_tmp = 64'h0;
      10'b1010001000:
        casez_tmp = 64'h0;
      10'b1010001001:
        casez_tmp = 64'h0;
      10'b1010001010:
        casez_tmp = 64'h0;
      10'b1010001011:
        casez_tmp = 64'h0;
      10'b1010001100:
        casez_tmp = 64'h0;
      10'b1010001101:
        casez_tmp = 64'h0;
      10'b1010001110:
        casez_tmp = 64'h0;
      10'b1010001111:
        casez_tmp = 64'h0;
      10'b1010010000:
        casez_tmp = 64'h0;
      10'b1010010001:
        casez_tmp = 64'h0;
      10'b1010010010:
        casez_tmp = 64'h0;
      10'b1010010011:
        casez_tmp = 64'h0;
      10'b1010010100:
        casez_tmp = 64'h0;
      10'b1010010101:
        casez_tmp = 64'h0;
      10'b1010010110:
        casez_tmp = 64'h0;
      10'b1010010111:
        casez_tmp = 64'h0;
      10'b1010011000:
        casez_tmp = 64'h0;
      10'b1010011001:
        casez_tmp = 64'h0;
      10'b1010011010:
        casez_tmp = 64'h0;
      10'b1010011011:
        casez_tmp = 64'h0;
      10'b1010011100:
        casez_tmp = 64'h0;
      10'b1010011101:
        casez_tmp = 64'h0;
      10'b1010011110:
        casez_tmp = 64'h0;
      10'b1010011111:
        casez_tmp = 64'h0;
      10'b1010100000:
        casez_tmp = 64'h0;
      10'b1010100001:
        casez_tmp = 64'h0;
      10'b1010100010:
        casez_tmp = 64'h0;
      10'b1010100011:
        casez_tmp = 64'h0;
      10'b1010100100:
        casez_tmp = 64'h0;
      10'b1010100101:
        casez_tmp = 64'h0;
      10'b1010100110:
        casez_tmp = 64'h0;
      10'b1010100111:
        casez_tmp = 64'h0;
      10'b1010101000:
        casez_tmp = 64'h0;
      10'b1010101001:
        casez_tmp = 64'h0;
      10'b1010101010:
        casez_tmp = 64'h0;
      10'b1010101011:
        casez_tmp = 64'h0;
      10'b1010101100:
        casez_tmp = 64'h0;
      10'b1010101101:
        casez_tmp = 64'h0;
      10'b1010101110:
        casez_tmp = 64'h0;
      10'b1010101111:
        casez_tmp = 64'h0;
      10'b1010110000:
        casez_tmp = 64'h0;
      10'b1010110001:
        casez_tmp = 64'h0;
      10'b1010110010:
        casez_tmp = 64'h0;
      10'b1010110011:
        casez_tmp = 64'h0;
      10'b1010110100:
        casez_tmp = 64'h0;
      10'b1010110101:
        casez_tmp = 64'h0;
      10'b1010110110:
        casez_tmp = 64'h0;
      10'b1010110111:
        casez_tmp = 64'h0;
      10'b1010111000:
        casez_tmp = 64'h0;
      10'b1010111001:
        casez_tmp = 64'h0;
      10'b1010111010:
        casez_tmp = 64'h0;
      10'b1010111011:
        casez_tmp = 64'h0;
      10'b1010111100:
        casez_tmp = 64'h0;
      10'b1010111101:
        casez_tmp = 64'h0;
      10'b1010111110:
        casez_tmp = 64'h0;
      10'b1010111111:
        casez_tmp = 64'h0;
      10'b1011000000:
        casez_tmp = 64'h0;
      10'b1011000001:
        casez_tmp = 64'h0;
      10'b1011000010:
        casez_tmp = 64'h0;
      10'b1011000011:
        casez_tmp = 64'h0;
      10'b1011000100:
        casez_tmp = 64'h0;
      10'b1011000101:
        casez_tmp = 64'h0;
      10'b1011000110:
        casez_tmp = 64'h0;
      10'b1011000111:
        casez_tmp = 64'h0;
      10'b1011001000:
        casez_tmp = 64'h0;
      10'b1011001001:
        casez_tmp = 64'h0;
      10'b1011001010:
        casez_tmp = 64'h0;
      10'b1011001011:
        casez_tmp = 64'h0;
      10'b1011001100:
        casez_tmp = 64'h0;
      10'b1011001101:
        casez_tmp = 64'h0;
      10'b1011001110:
        casez_tmp = 64'h0;
      10'b1011001111:
        casez_tmp = 64'h0;
      10'b1011010000:
        casez_tmp = 64'h0;
      10'b1011010001:
        casez_tmp = 64'h0;
      10'b1011010010:
        casez_tmp = 64'h0;
      10'b1011010011:
        casez_tmp = 64'h0;
      10'b1011010100:
        casez_tmp = 64'h0;
      10'b1011010101:
        casez_tmp = 64'h0;
      10'b1011010110:
        casez_tmp = 64'h0;
      10'b1011010111:
        casez_tmp = 64'h0;
      10'b1011011000:
        casez_tmp = 64'h0;
      10'b1011011001:
        casez_tmp = 64'h0;
      10'b1011011010:
        casez_tmp = 64'h0;
      10'b1011011011:
        casez_tmp = 64'h0;
      10'b1011011100:
        casez_tmp = 64'h0;
      10'b1011011101:
        casez_tmp = 64'h0;
      10'b1011011110:
        casez_tmp = 64'h0;
      10'b1011011111:
        casez_tmp = 64'h0;
      10'b1011100000:
        casez_tmp = 64'h0;
      10'b1011100001:
        casez_tmp = 64'h0;
      10'b1011100010:
        casez_tmp = 64'h0;
      10'b1011100011:
        casez_tmp = 64'h0;
      10'b1011100100:
        casez_tmp = 64'h0;
      10'b1011100101:
        casez_tmp = 64'h0;
      10'b1011100110:
        casez_tmp = 64'h0;
      10'b1011100111:
        casez_tmp = 64'h0;
      10'b1011101000:
        casez_tmp = 64'h0;
      10'b1011101001:
        casez_tmp = 64'h0;
      10'b1011101010:
        casez_tmp = 64'h0;
      10'b1011101011:
        casez_tmp = 64'h0;
      10'b1011101100:
        casez_tmp = 64'h0;
      10'b1011101101:
        casez_tmp = 64'h0;
      10'b1011101110:
        casez_tmp = 64'h0;
      10'b1011101111:
        casez_tmp = 64'h0;
      10'b1011110000:
        casez_tmp = 64'h0;
      10'b1011110001:
        casez_tmp = 64'h0;
      10'b1011110010:
        casez_tmp = 64'h0;
      10'b1011110011:
        casez_tmp = 64'h0;
      10'b1011110100:
        casez_tmp = 64'h0;
      10'b1011110101:
        casez_tmp = 64'h0;
      10'b1011110110:
        casez_tmp = 64'h0;
      10'b1011110111:
        casez_tmp = 64'h0;
      10'b1011111000:
        casez_tmp = 64'h0;
      10'b1011111001:
        casez_tmp = 64'h0;
      10'b1011111010:
        casez_tmp = 64'h0;
      10'b1011111011:
        casez_tmp = 64'h0;
      10'b1011111100:
        casez_tmp = 64'h0;
      10'b1011111101:
        casez_tmp = 64'h0;
      10'b1011111110:
        casez_tmp = 64'h0;
      10'b1011111111:
        casez_tmp = 64'h0;
      10'b1100000000:
        casez_tmp = 64'h0;
      10'b1100000001:
        casez_tmp = 64'h0;
      10'b1100000010:
        casez_tmp = 64'h0;
      10'b1100000011:
        casez_tmp = 64'h0;
      10'b1100000100:
        casez_tmp = 64'h0;
      10'b1100000101:
        casez_tmp = 64'h0;
      10'b1100000110:
        casez_tmp = 64'h0;
      10'b1100000111:
        casez_tmp = 64'h0;
      10'b1100001000:
        casez_tmp = 64'h0;
      10'b1100001001:
        casez_tmp = 64'h0;
      10'b1100001010:
        casez_tmp = 64'h0;
      10'b1100001011:
        casez_tmp = 64'h0;
      10'b1100001100:
        casez_tmp = 64'h0;
      10'b1100001101:
        casez_tmp = 64'h0;
      10'b1100001110:
        casez_tmp = 64'h0;
      10'b1100001111:
        casez_tmp = 64'h0;
      10'b1100010000:
        casez_tmp = 64'h0;
      10'b1100010001:
        casez_tmp = 64'h0;
      10'b1100010010:
        casez_tmp = 64'h0;
      10'b1100010011:
        casez_tmp = 64'h0;
      10'b1100010100:
        casez_tmp = 64'h0;
      10'b1100010101:
        casez_tmp = 64'h0;
      10'b1100010110:
        casez_tmp = 64'h0;
      10'b1100010111:
        casez_tmp = 64'h0;
      10'b1100011000:
        casez_tmp = 64'h0;
      10'b1100011001:
        casez_tmp = 64'h0;
      10'b1100011010:
        casez_tmp = 64'h0;
      10'b1100011011:
        casez_tmp = 64'h0;
      10'b1100011100:
        casez_tmp = 64'h0;
      10'b1100011101:
        casez_tmp = 64'h0;
      10'b1100011110:
        casez_tmp = 64'h0;
      10'b1100011111:
        casez_tmp = 64'h0;
      10'b1100100000:
        casez_tmp = 64'h0;
      10'b1100100001:
        casez_tmp = 64'h0;
      10'b1100100010:
        casez_tmp = 64'h0;
      10'b1100100011:
        casez_tmp = 64'h0;
      10'b1100100100:
        casez_tmp = 64'h0;
      10'b1100100101:
        casez_tmp = 64'h0;
      10'b1100100110:
        casez_tmp = 64'h0;
      10'b1100100111:
        casez_tmp = 64'h0;
      10'b1100101000:
        casez_tmp = 64'h0;
      10'b1100101001:
        casez_tmp = 64'h0;
      10'b1100101010:
        casez_tmp = 64'h0;
      10'b1100101011:
        casez_tmp = 64'h0;
      10'b1100101100:
        casez_tmp = 64'h0;
      10'b1100101101:
        casez_tmp = 64'h0;
      10'b1100101110:
        casez_tmp = 64'h0;
      10'b1100101111:
        casez_tmp = 64'h0;
      10'b1100110000:
        casez_tmp = 64'h0;
      10'b1100110001:
        casez_tmp = 64'h0;
      10'b1100110010:
        casez_tmp = 64'h0;
      10'b1100110011:
        casez_tmp = 64'h0;
      10'b1100110100:
        casez_tmp = 64'h0;
      10'b1100110101:
        casez_tmp = 64'h0;
      10'b1100110110:
        casez_tmp = 64'h0;
      10'b1100110111:
        casez_tmp = 64'h0;
      10'b1100111000:
        casez_tmp = 64'h0;
      10'b1100111001:
        casez_tmp = 64'h0;
      10'b1100111010:
        casez_tmp = 64'h0;
      10'b1100111011:
        casez_tmp = 64'h0;
      10'b1100111100:
        casez_tmp = 64'h0;
      10'b1100111101:
        casez_tmp = 64'h0;
      10'b1100111110:
        casez_tmp = 64'h0;
      10'b1100111111:
        casez_tmp = 64'h0;
      10'b1101000000:
        casez_tmp = 64'h0;
      10'b1101000001:
        casez_tmp = 64'h0;
      10'b1101000010:
        casez_tmp = 64'h0;
      10'b1101000011:
        casez_tmp = 64'h0;
      10'b1101000100:
        casez_tmp = 64'h0;
      10'b1101000101:
        casez_tmp = 64'h0;
      10'b1101000110:
        casez_tmp = 64'h0;
      10'b1101000111:
        casez_tmp = 64'h0;
      10'b1101001000:
        casez_tmp = 64'h0;
      10'b1101001001:
        casez_tmp = 64'h0;
      10'b1101001010:
        casez_tmp = 64'h0;
      10'b1101001011:
        casez_tmp = 64'h0;
      10'b1101001100:
        casez_tmp = 64'h0;
      10'b1101001101:
        casez_tmp = 64'h0;
      10'b1101001110:
        casez_tmp = 64'h0;
      10'b1101001111:
        casez_tmp = 64'h0;
      10'b1101010000:
        casez_tmp = 64'h0;
      10'b1101010001:
        casez_tmp = 64'h0;
      10'b1101010010:
        casez_tmp = 64'h0;
      10'b1101010011:
        casez_tmp = 64'h0;
      10'b1101010100:
        casez_tmp = 64'h0;
      10'b1101010101:
        casez_tmp = 64'h0;
      10'b1101010110:
        casez_tmp = 64'h0;
      10'b1101010111:
        casez_tmp = 64'h0;
      10'b1101011000:
        casez_tmp = 64'h0;
      10'b1101011001:
        casez_tmp = 64'h0;
      10'b1101011010:
        casez_tmp = 64'h0;
      10'b1101011011:
        casez_tmp = 64'h0;
      10'b1101011100:
        casez_tmp = 64'h0;
      10'b1101011101:
        casez_tmp = 64'h0;
      10'b1101011110:
        casez_tmp = 64'h0;
      10'b1101011111:
        casez_tmp = 64'h0;
      10'b1101100000:
        casez_tmp = 64'h0;
      10'b1101100001:
        casez_tmp = 64'h0;
      10'b1101100010:
        casez_tmp = 64'h0;
      10'b1101100011:
        casez_tmp = 64'h0;
      10'b1101100100:
        casez_tmp = 64'h0;
      10'b1101100101:
        casez_tmp = 64'h0;
      10'b1101100110:
        casez_tmp = 64'h0;
      10'b1101100111:
        casez_tmp = 64'h0;
      10'b1101101000:
        casez_tmp = 64'h0;
      10'b1101101001:
        casez_tmp = 64'h0;
      10'b1101101010:
        casez_tmp = 64'h0;
      10'b1101101011:
        casez_tmp = 64'h0;
      10'b1101101100:
        casez_tmp = 64'h0;
      10'b1101101101:
        casez_tmp = 64'h0;
      10'b1101101110:
        casez_tmp = 64'h0;
      10'b1101101111:
        casez_tmp = 64'h0;
      10'b1101110000:
        casez_tmp = 64'h0;
      10'b1101110001:
        casez_tmp = 64'h0;
      10'b1101110010:
        casez_tmp = 64'h0;
      10'b1101110011:
        casez_tmp = 64'h0;
      10'b1101110100:
        casez_tmp = 64'h0;
      10'b1101110101:
        casez_tmp = 64'h0;
      10'b1101110110:
        casez_tmp = 64'h0;
      10'b1101110111:
        casez_tmp = 64'h0;
      10'b1101111000:
        casez_tmp = 64'h0;
      10'b1101111001:
        casez_tmp = 64'h0;
      10'b1101111010:
        casez_tmp = 64'h0;
      10'b1101111011:
        casez_tmp = 64'h0;
      10'b1101111100:
        casez_tmp = 64'h0;
      10'b1101111101:
        casez_tmp = 64'h0;
      10'b1101111110:
        casez_tmp = 64'h0;
      10'b1101111111:
        casez_tmp = 64'h0;
      10'b1110000000:
        casez_tmp = 64'h0;
      10'b1110000001:
        casez_tmp = 64'h0;
      10'b1110000010:
        casez_tmp = 64'h0;
      10'b1110000011:
        casez_tmp = 64'h0;
      10'b1110000100:
        casez_tmp = 64'h0;
      10'b1110000101:
        casez_tmp = 64'h0;
      10'b1110000110:
        casez_tmp = 64'h0;
      10'b1110000111:
        casez_tmp = 64'h0;
      10'b1110001000:
        casez_tmp = 64'h0;
      10'b1110001001:
        casez_tmp = 64'h0;
      10'b1110001010:
        casez_tmp = 64'h0;
      10'b1110001011:
        casez_tmp = 64'h0;
      10'b1110001100:
        casez_tmp = 64'h0;
      10'b1110001101:
        casez_tmp = 64'h0;
      10'b1110001110:
        casez_tmp = 64'h0;
      10'b1110001111:
        casez_tmp = 64'h0;
      10'b1110010000:
        casez_tmp = 64'h0;
      10'b1110010001:
        casez_tmp = 64'h0;
      10'b1110010010:
        casez_tmp = 64'h0;
      10'b1110010011:
        casez_tmp = 64'h0;
      10'b1110010100:
        casez_tmp = 64'h0;
      10'b1110010101:
        casez_tmp = 64'h0;
      10'b1110010110:
        casez_tmp = 64'h0;
      10'b1110010111:
        casez_tmp = 64'h0;
      10'b1110011000:
        casez_tmp = 64'h0;
      10'b1110011001:
        casez_tmp = 64'h0;
      10'b1110011010:
        casez_tmp = 64'h0;
      10'b1110011011:
        casez_tmp = 64'h0;
      10'b1110011100:
        casez_tmp = 64'h0;
      10'b1110011101:
        casez_tmp = 64'h0;
      10'b1110011110:
        casez_tmp = 64'h0;
      10'b1110011111:
        casez_tmp = 64'h0;
      10'b1110100000:
        casez_tmp = 64'h0;
      10'b1110100001:
        casez_tmp = 64'h0;
      10'b1110100010:
        casez_tmp = 64'h0;
      10'b1110100011:
        casez_tmp = 64'h0;
      10'b1110100100:
        casez_tmp = 64'h0;
      10'b1110100101:
        casez_tmp = 64'h0;
      10'b1110100110:
        casez_tmp = 64'h0;
      10'b1110100111:
        casez_tmp = 64'h0;
      10'b1110101000:
        casez_tmp = 64'h0;
      10'b1110101001:
        casez_tmp = 64'h0;
      10'b1110101010:
        casez_tmp = 64'h0;
      10'b1110101011:
        casez_tmp = 64'h0;
      10'b1110101100:
        casez_tmp = 64'h0;
      10'b1110101101:
        casez_tmp = 64'h0;
      10'b1110101110:
        casez_tmp = 64'h0;
      10'b1110101111:
        casez_tmp = 64'h0;
      10'b1110110000:
        casez_tmp = 64'h0;
      10'b1110110001:
        casez_tmp = 64'h0;
      10'b1110110010:
        casez_tmp = 64'h0;
      10'b1110110011:
        casez_tmp = 64'h0;
      10'b1110110100:
        casez_tmp = 64'h0;
      10'b1110110101:
        casez_tmp = 64'h0;
      10'b1110110110:
        casez_tmp = 64'h0;
      10'b1110110111:
        casez_tmp = 64'h0;
      10'b1110111000:
        casez_tmp = 64'h0;
      10'b1110111001:
        casez_tmp = 64'h0;
      10'b1110111010:
        casez_tmp = 64'h0;
      10'b1110111011:
        casez_tmp = 64'h0;
      10'b1110111100:
        casez_tmp = 64'h0;
      10'b1110111101:
        casez_tmp = 64'h0;
      10'b1110111110:
        casez_tmp = 64'h0;
      10'b1110111111:
        casez_tmp = 64'h0;
      10'b1111000000:
        casez_tmp = 64'h0;
      10'b1111000001:
        casez_tmp = 64'h0;
      10'b1111000010:
        casez_tmp = 64'h0;
      10'b1111000011:
        casez_tmp = 64'h0;
      10'b1111000100:
        casez_tmp = 64'h0;
      10'b1111000101:
        casez_tmp = 64'h0;
      10'b1111000110:
        casez_tmp = 64'h0;
      10'b1111000111:
        casez_tmp = 64'h0;
      10'b1111001000:
        casez_tmp = 64'h0;
      10'b1111001001:
        casez_tmp = 64'h0;
      10'b1111001010:
        casez_tmp = 64'h0;
      10'b1111001011:
        casez_tmp = 64'h0;
      10'b1111001100:
        casez_tmp = 64'h0;
      10'b1111001101:
        casez_tmp = 64'h0;
      10'b1111001110:
        casez_tmp = 64'h0;
      10'b1111001111:
        casez_tmp = 64'h0;
      10'b1111010000:
        casez_tmp = 64'h0;
      10'b1111010001:
        casez_tmp = 64'h0;
      10'b1111010010:
        casez_tmp = 64'h0;
      10'b1111010011:
        casez_tmp = 64'h0;
      10'b1111010100:
        casez_tmp = 64'h0;
      10'b1111010101:
        casez_tmp = 64'h0;
      10'b1111010110:
        casez_tmp = 64'h0;
      10'b1111010111:
        casez_tmp = 64'h0;
      10'b1111011000:
        casez_tmp = 64'h0;
      10'b1111011001:
        casez_tmp = 64'h0;
      10'b1111011010:
        casez_tmp = 64'h0;
      10'b1111011011:
        casez_tmp = 64'h0;
      10'b1111011100:
        casez_tmp = 64'h0;
      10'b1111011101:
        casez_tmp = 64'h0;
      10'b1111011110:
        casez_tmp = 64'h0;
      10'b1111011111:
        casez_tmp = 64'h0;
      10'b1111100000:
        casez_tmp = 64'h0;
      10'b1111100001:
        casez_tmp = 64'h0;
      10'b1111100010:
        casez_tmp = 64'h0;
      10'b1111100011:
        casez_tmp = 64'h0;
      10'b1111100100:
        casez_tmp = 64'h0;
      10'b1111100101:
        casez_tmp = 64'h0;
      10'b1111100110:
        casez_tmp = 64'h0;
      10'b1111100111:
        casez_tmp = 64'h0;
      10'b1111101000:
        casez_tmp = 64'h0;
      10'b1111101001:
        casez_tmp = 64'h0;
      10'b1111101010:
        casez_tmp = 64'h0;
      10'b1111101011:
        casez_tmp = 64'h0;
      10'b1111101100:
        casez_tmp = 64'h0;
      10'b1111101101:
        casez_tmp = 64'h0;
      10'b1111101110:
        casez_tmp = 64'h0;
      10'b1111101111:
        casez_tmp = 64'h0;
      10'b1111110000:
        casez_tmp = 64'h0;
      10'b1111110001:
        casez_tmp = 64'h0;
      10'b1111110010:
        casez_tmp = 64'h0;
      10'b1111110011:
        casez_tmp = 64'h0;
      10'b1111110100:
        casez_tmp = 64'h0;
      10'b1111110101:
        casez_tmp = 64'h0;
      10'b1111110110:
        casez_tmp = 64'h0;
      10'b1111110111:
        casez_tmp = 64'h0;
      10'b1111111000:
        casez_tmp = 64'h0;
      10'b1111111001:
        casez_tmp = 64'h0;
      10'b1111111010:
        casez_tmp = 64'h0;
      10'b1111111011:
        casez_tmp = 64'h0;
      10'b1111111100:
        casez_tmp = 64'h0;
      10'b1111111101:
        casez_tmp = 64'h0;
      10'b1111111110:
        casez_tmp = 64'h0;
      default:
        casez_tmp = 64'h0;
    endcase
  end // always @(*)
  TLMonitor_54 monitor (
    .clock                (clock),
    .reset                (reset),
    .io_in_a_ready        (auto_in_d_ready),
    .io_in_a_valid        (auto_in_a_valid),
    .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
    .io_in_a_bits_param   (auto_in_a_bits_param),
    .io_in_a_bits_size    (auto_in_a_bits_size),
    .io_in_a_bits_source  (auto_in_a_bits_source),
    .io_in_a_bits_address (auto_in_a_bits_address),
    .io_in_a_bits_mask    (auto_in_a_bits_mask),
    .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
    .io_in_d_ready        (auto_in_d_ready),
    .io_in_d_valid        (auto_in_a_valid),
    .io_in_d_bits_size    (auto_in_a_bits_size),
    .io_in_d_bits_source  (auto_in_a_bits_source)
  );
  assign auto_in_a_ready = auto_in_d_ready;
  assign auto_in_d_valid = auto_in_a_valid;
  assign auto_in_d_bits_size = auto_in_a_bits_size;
  assign auto_in_d_bits_source = auto_in_a_bits_source;
  assign auto_in_d_bits_data = (|(auto_in_a_bits_address[15:13])) ? 64'h0 : casez_tmp;
endmodule

