// Standard header to adapt well known macros for prints and assertions.

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module IntSyncCrossingSource_5(
  input  clock,
         reset,
         auto_in_0,
         auto_in_1,
  output auto_out_sync_0,
         auto_out_sync_1
);

  wire [1:0] _reg_io_q;
  AsyncResetRegVec_w2_i0 reg_0 (
    .clock (clock),
    .reset (reset),
    .io_d  ({auto_in_1, auto_in_0}),
    .io_q  (_reg_io_q)
  );
  assign auto_out_sync_0 = _reg_io_q[0];
  assign auto_out_sync_1 = _reg_io_q[1];
endmodule

