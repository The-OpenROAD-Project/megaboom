// Standard header to adapt well known macros for prints and assertions.

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module ResetCatchAndSync_d3(
  input  clock,
         reset,
  output io_sync_reset
);

  wire _io_sync_reset_chain_io_q;
  AsyncResetSynchronizerShiftReg_w1_d3_i0 io_sync_reset_chain (
    .clock (clock),
    .reset (reset),
    .io_d  (1'h1),
    .io_q  (_io_sync_reset_chain_io_q)
  );
  assign io_sync_reset = ~_io_sync_reset_chain_io_q;
endmodule

