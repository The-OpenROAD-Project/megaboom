// Standard header to adapt well known macros for prints and assertions.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module Arbiter_5(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [6:0]  io_in_0_bits_uop_uopc,
  input  [31:0] io_in_0_bits_uop_inst,
                io_in_0_bits_uop_debug_inst,
  input         io_in_0_bits_uop_is_rvc,
  input  [39:0] io_in_0_bits_uop_debug_pc,
  input  [2:0]  io_in_0_bits_uop_iq_type,
  input  [9:0]  io_in_0_bits_uop_fu_code,
  input  [3:0]  io_in_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_0_bits_uop_ctrl_op2_sel,
                io_in_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_0_bits_uop_ctrl_op_fcn,
  input         io_in_0_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_0_bits_uop_ctrl_csr_cmd,
  input         io_in_0_bits_uop_ctrl_is_load,
                io_in_0_bits_uop_ctrl_is_sta,
                io_in_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_0_bits_uop_iw_state,
  input         io_in_0_bits_uop_iw_p1_poisoned,
                io_in_0_bits_uop_iw_p2_poisoned,
                io_in_0_bits_uop_is_br,
                io_in_0_bits_uop_is_jalr,
                io_in_0_bits_uop_is_jal,
                io_in_0_bits_uop_is_sfb,
  input  [19:0] io_in_0_bits_uop_br_mask,
  input  [4:0]  io_in_0_bits_uop_br_tag,
  input  [5:0]  io_in_0_bits_uop_ftq_idx,
  input         io_in_0_bits_uop_edge_inst,
  input  [5:0]  io_in_0_bits_uop_pc_lob,
  input         io_in_0_bits_uop_taken,
  input  [19:0] io_in_0_bits_uop_imm_packed,
  input  [11:0] io_in_0_bits_uop_csr_addr,
  input  [6:0]  io_in_0_bits_uop_rob_idx,
  input  [4:0]  io_in_0_bits_uop_ldq_idx,
                io_in_0_bits_uop_stq_idx,
  input  [1:0]  io_in_0_bits_uop_rxq_idx,
  input  [6:0]  io_in_0_bits_uop_pdst,
                io_in_0_bits_uop_prs1,
                io_in_0_bits_uop_prs2,
                io_in_0_bits_uop_prs3,
  input  [5:0]  io_in_0_bits_uop_ppred,
  input         io_in_0_bits_uop_prs1_busy,
                io_in_0_bits_uop_prs2_busy,
                io_in_0_bits_uop_prs3_busy,
                io_in_0_bits_uop_ppred_busy,
  input  [6:0]  io_in_0_bits_uop_stale_pdst,
  input         io_in_0_bits_uop_exception,
  input  [63:0] io_in_0_bits_uop_exc_cause,
  input         io_in_0_bits_uop_bypassable,
  input  [4:0]  io_in_0_bits_uop_mem_cmd,
  input  [1:0]  io_in_0_bits_uop_mem_size,
  input         io_in_0_bits_uop_mem_signed,
                io_in_0_bits_uop_is_fence,
                io_in_0_bits_uop_is_fencei,
                io_in_0_bits_uop_is_amo,
                io_in_0_bits_uop_uses_ldq,
                io_in_0_bits_uop_uses_stq,
                io_in_0_bits_uop_is_sys_pc2epc,
                io_in_0_bits_uop_is_unique,
                io_in_0_bits_uop_flush_on_commit,
                io_in_0_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_0_bits_uop_ldst,
                io_in_0_bits_uop_lrs1,
                io_in_0_bits_uop_lrs2,
                io_in_0_bits_uop_lrs3,
  input         io_in_0_bits_uop_ldst_val,
  input  [1:0]  io_in_0_bits_uop_dst_rtype,
                io_in_0_bits_uop_lrs1_rtype,
                io_in_0_bits_uop_lrs2_rtype,
  input         io_in_0_bits_uop_frs3_en,
                io_in_0_bits_uop_fp_val,
                io_in_0_bits_uop_fp_single,
                io_in_0_bits_uop_xcpt_pf_if,
                io_in_0_bits_uop_xcpt_ae_if,
                io_in_0_bits_uop_xcpt_ma_if,
                io_in_0_bits_uop_bp_debug_if,
                io_in_0_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_0_bits_uop_debug_fsrc,
                io_in_0_bits_uop_debug_tsrc,
  input  [39:0] io_in_0_bits_addr,
  input         io_in_0_bits_is_hella,
  input  [7:0]  io_in_0_bits_way_en,
  input  [4:0]  io_in_0_bits_sdq_id,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [6:0]  io_in_1_bits_uop_uopc,
  input  [31:0] io_in_1_bits_uop_inst,
                io_in_1_bits_uop_debug_inst,
  input         io_in_1_bits_uop_is_rvc,
  input  [39:0] io_in_1_bits_uop_debug_pc,
  input  [2:0]  io_in_1_bits_uop_iq_type,
  input  [9:0]  io_in_1_bits_uop_fu_code,
  input  [3:0]  io_in_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_1_bits_uop_ctrl_op2_sel,
                io_in_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_1_bits_uop_ctrl_op_fcn,
  input         io_in_1_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_1_bits_uop_ctrl_csr_cmd,
  input         io_in_1_bits_uop_ctrl_is_load,
                io_in_1_bits_uop_ctrl_is_sta,
                io_in_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_1_bits_uop_iw_state,
  input         io_in_1_bits_uop_iw_p1_poisoned,
                io_in_1_bits_uop_iw_p2_poisoned,
                io_in_1_bits_uop_is_br,
                io_in_1_bits_uop_is_jalr,
                io_in_1_bits_uop_is_jal,
                io_in_1_bits_uop_is_sfb,
  input  [19:0] io_in_1_bits_uop_br_mask,
  input  [4:0]  io_in_1_bits_uop_br_tag,
  input  [5:0]  io_in_1_bits_uop_ftq_idx,
  input         io_in_1_bits_uop_edge_inst,
  input  [5:0]  io_in_1_bits_uop_pc_lob,
  input         io_in_1_bits_uop_taken,
  input  [19:0] io_in_1_bits_uop_imm_packed,
  input  [11:0] io_in_1_bits_uop_csr_addr,
  input  [6:0]  io_in_1_bits_uop_rob_idx,
  input  [4:0]  io_in_1_bits_uop_ldq_idx,
                io_in_1_bits_uop_stq_idx,
  input  [1:0]  io_in_1_bits_uop_rxq_idx,
  input  [6:0]  io_in_1_bits_uop_pdst,
                io_in_1_bits_uop_prs1,
                io_in_1_bits_uop_prs2,
                io_in_1_bits_uop_prs3,
  input  [5:0]  io_in_1_bits_uop_ppred,
  input         io_in_1_bits_uop_prs1_busy,
                io_in_1_bits_uop_prs2_busy,
                io_in_1_bits_uop_prs3_busy,
                io_in_1_bits_uop_ppred_busy,
  input  [6:0]  io_in_1_bits_uop_stale_pdst,
  input         io_in_1_bits_uop_exception,
  input  [63:0] io_in_1_bits_uop_exc_cause,
  input         io_in_1_bits_uop_bypassable,
  input  [4:0]  io_in_1_bits_uop_mem_cmd,
  input  [1:0]  io_in_1_bits_uop_mem_size,
  input         io_in_1_bits_uop_mem_signed,
                io_in_1_bits_uop_is_fence,
                io_in_1_bits_uop_is_fencei,
                io_in_1_bits_uop_is_amo,
                io_in_1_bits_uop_uses_ldq,
                io_in_1_bits_uop_uses_stq,
                io_in_1_bits_uop_is_sys_pc2epc,
                io_in_1_bits_uop_is_unique,
                io_in_1_bits_uop_flush_on_commit,
                io_in_1_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_1_bits_uop_ldst,
                io_in_1_bits_uop_lrs1,
                io_in_1_bits_uop_lrs2,
                io_in_1_bits_uop_lrs3,
  input         io_in_1_bits_uop_ldst_val,
  input  [1:0]  io_in_1_bits_uop_dst_rtype,
                io_in_1_bits_uop_lrs1_rtype,
                io_in_1_bits_uop_lrs2_rtype,
  input         io_in_1_bits_uop_frs3_en,
                io_in_1_bits_uop_fp_val,
                io_in_1_bits_uop_fp_single,
                io_in_1_bits_uop_xcpt_pf_if,
                io_in_1_bits_uop_xcpt_ae_if,
                io_in_1_bits_uop_xcpt_ma_if,
                io_in_1_bits_uop_bp_debug_if,
                io_in_1_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_1_bits_uop_debug_fsrc,
                io_in_1_bits_uop_debug_tsrc,
  input  [39:0] io_in_1_bits_addr,
  input         io_in_1_bits_is_hella,
  input  [7:0]  io_in_1_bits_way_en,
  input  [4:0]  io_in_1_bits_sdq_id,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [6:0]  io_in_2_bits_uop_uopc,
  input  [31:0] io_in_2_bits_uop_inst,
                io_in_2_bits_uop_debug_inst,
  input         io_in_2_bits_uop_is_rvc,
  input  [39:0] io_in_2_bits_uop_debug_pc,
  input  [2:0]  io_in_2_bits_uop_iq_type,
  input  [9:0]  io_in_2_bits_uop_fu_code,
  input  [3:0]  io_in_2_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_2_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_2_bits_uop_ctrl_op2_sel,
                io_in_2_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_2_bits_uop_ctrl_op_fcn,
  input         io_in_2_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_2_bits_uop_ctrl_csr_cmd,
  input         io_in_2_bits_uop_ctrl_is_load,
                io_in_2_bits_uop_ctrl_is_sta,
                io_in_2_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_2_bits_uop_iw_state,
  input         io_in_2_bits_uop_iw_p1_poisoned,
                io_in_2_bits_uop_iw_p2_poisoned,
                io_in_2_bits_uop_is_br,
                io_in_2_bits_uop_is_jalr,
                io_in_2_bits_uop_is_jal,
                io_in_2_bits_uop_is_sfb,
  input  [19:0] io_in_2_bits_uop_br_mask,
  input  [4:0]  io_in_2_bits_uop_br_tag,
  input  [5:0]  io_in_2_bits_uop_ftq_idx,
  input         io_in_2_bits_uop_edge_inst,
  input  [5:0]  io_in_2_bits_uop_pc_lob,
  input         io_in_2_bits_uop_taken,
  input  [19:0] io_in_2_bits_uop_imm_packed,
  input  [11:0] io_in_2_bits_uop_csr_addr,
  input  [6:0]  io_in_2_bits_uop_rob_idx,
  input  [4:0]  io_in_2_bits_uop_ldq_idx,
                io_in_2_bits_uop_stq_idx,
  input  [1:0]  io_in_2_bits_uop_rxq_idx,
  input  [6:0]  io_in_2_bits_uop_pdst,
                io_in_2_bits_uop_prs1,
                io_in_2_bits_uop_prs2,
                io_in_2_bits_uop_prs3,
  input  [5:0]  io_in_2_bits_uop_ppred,
  input         io_in_2_bits_uop_prs1_busy,
                io_in_2_bits_uop_prs2_busy,
                io_in_2_bits_uop_prs3_busy,
                io_in_2_bits_uop_ppred_busy,
  input  [6:0]  io_in_2_bits_uop_stale_pdst,
  input         io_in_2_bits_uop_exception,
  input  [63:0] io_in_2_bits_uop_exc_cause,
  input         io_in_2_bits_uop_bypassable,
  input  [4:0]  io_in_2_bits_uop_mem_cmd,
  input  [1:0]  io_in_2_bits_uop_mem_size,
  input         io_in_2_bits_uop_mem_signed,
                io_in_2_bits_uop_is_fence,
                io_in_2_bits_uop_is_fencei,
                io_in_2_bits_uop_is_amo,
                io_in_2_bits_uop_uses_ldq,
                io_in_2_bits_uop_uses_stq,
                io_in_2_bits_uop_is_sys_pc2epc,
                io_in_2_bits_uop_is_unique,
                io_in_2_bits_uop_flush_on_commit,
                io_in_2_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_2_bits_uop_ldst,
                io_in_2_bits_uop_lrs1,
                io_in_2_bits_uop_lrs2,
                io_in_2_bits_uop_lrs3,
  input         io_in_2_bits_uop_ldst_val,
  input  [1:0]  io_in_2_bits_uop_dst_rtype,
                io_in_2_bits_uop_lrs1_rtype,
                io_in_2_bits_uop_lrs2_rtype,
  input         io_in_2_bits_uop_frs3_en,
                io_in_2_bits_uop_fp_val,
                io_in_2_bits_uop_fp_single,
                io_in_2_bits_uop_xcpt_pf_if,
                io_in_2_bits_uop_xcpt_ae_if,
                io_in_2_bits_uop_xcpt_ma_if,
                io_in_2_bits_uop_bp_debug_if,
                io_in_2_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_2_bits_uop_debug_fsrc,
                io_in_2_bits_uop_debug_tsrc,
  input  [39:0] io_in_2_bits_addr,
  input         io_in_2_bits_is_hella,
  input  [7:0]  io_in_2_bits_way_en,
  input  [4:0]  io_in_2_bits_sdq_id,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [6:0]  io_in_3_bits_uop_uopc,
  input  [31:0] io_in_3_bits_uop_inst,
                io_in_3_bits_uop_debug_inst,
  input         io_in_3_bits_uop_is_rvc,
  input  [39:0] io_in_3_bits_uop_debug_pc,
  input  [2:0]  io_in_3_bits_uop_iq_type,
  input  [9:0]  io_in_3_bits_uop_fu_code,
  input  [3:0]  io_in_3_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_3_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_3_bits_uop_ctrl_op2_sel,
                io_in_3_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_3_bits_uop_ctrl_op_fcn,
  input         io_in_3_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_3_bits_uop_ctrl_csr_cmd,
  input         io_in_3_bits_uop_ctrl_is_load,
                io_in_3_bits_uop_ctrl_is_sta,
                io_in_3_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_3_bits_uop_iw_state,
  input         io_in_3_bits_uop_iw_p1_poisoned,
                io_in_3_bits_uop_iw_p2_poisoned,
                io_in_3_bits_uop_is_br,
                io_in_3_bits_uop_is_jalr,
                io_in_3_bits_uop_is_jal,
                io_in_3_bits_uop_is_sfb,
  input  [19:0] io_in_3_bits_uop_br_mask,
  input  [4:0]  io_in_3_bits_uop_br_tag,
  input  [5:0]  io_in_3_bits_uop_ftq_idx,
  input         io_in_3_bits_uop_edge_inst,
  input  [5:0]  io_in_3_bits_uop_pc_lob,
  input         io_in_3_bits_uop_taken,
  input  [19:0] io_in_3_bits_uop_imm_packed,
  input  [11:0] io_in_3_bits_uop_csr_addr,
  input  [6:0]  io_in_3_bits_uop_rob_idx,
  input  [4:0]  io_in_3_bits_uop_ldq_idx,
                io_in_3_bits_uop_stq_idx,
  input  [1:0]  io_in_3_bits_uop_rxq_idx,
  input  [6:0]  io_in_3_bits_uop_pdst,
                io_in_3_bits_uop_prs1,
                io_in_3_bits_uop_prs2,
                io_in_3_bits_uop_prs3,
  input  [5:0]  io_in_3_bits_uop_ppred,
  input         io_in_3_bits_uop_prs1_busy,
                io_in_3_bits_uop_prs2_busy,
                io_in_3_bits_uop_prs3_busy,
                io_in_3_bits_uop_ppred_busy,
  input  [6:0]  io_in_3_bits_uop_stale_pdst,
  input         io_in_3_bits_uop_exception,
  input  [63:0] io_in_3_bits_uop_exc_cause,
  input         io_in_3_bits_uop_bypassable,
  input  [4:0]  io_in_3_bits_uop_mem_cmd,
  input  [1:0]  io_in_3_bits_uop_mem_size,
  input         io_in_3_bits_uop_mem_signed,
                io_in_3_bits_uop_is_fence,
                io_in_3_bits_uop_is_fencei,
                io_in_3_bits_uop_is_amo,
                io_in_3_bits_uop_uses_ldq,
                io_in_3_bits_uop_uses_stq,
                io_in_3_bits_uop_is_sys_pc2epc,
                io_in_3_bits_uop_is_unique,
                io_in_3_bits_uop_flush_on_commit,
                io_in_3_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_3_bits_uop_ldst,
                io_in_3_bits_uop_lrs1,
                io_in_3_bits_uop_lrs2,
                io_in_3_bits_uop_lrs3,
  input         io_in_3_bits_uop_ldst_val,
  input  [1:0]  io_in_3_bits_uop_dst_rtype,
                io_in_3_bits_uop_lrs1_rtype,
                io_in_3_bits_uop_lrs2_rtype,
  input         io_in_3_bits_uop_frs3_en,
                io_in_3_bits_uop_fp_val,
                io_in_3_bits_uop_fp_single,
                io_in_3_bits_uop_xcpt_pf_if,
                io_in_3_bits_uop_xcpt_ae_if,
                io_in_3_bits_uop_xcpt_ma_if,
                io_in_3_bits_uop_bp_debug_if,
                io_in_3_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_3_bits_uop_debug_fsrc,
                io_in_3_bits_uop_debug_tsrc,
  input  [39:0] io_in_3_bits_addr,
  input         io_in_3_bits_is_hella,
  input  [7:0]  io_in_3_bits_way_en,
  input  [4:0]  io_in_3_bits_sdq_id,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [6:0]  io_in_4_bits_uop_uopc,
  input  [31:0] io_in_4_bits_uop_inst,
                io_in_4_bits_uop_debug_inst,
  input         io_in_4_bits_uop_is_rvc,
  input  [39:0] io_in_4_bits_uop_debug_pc,
  input  [2:0]  io_in_4_bits_uop_iq_type,
  input  [9:0]  io_in_4_bits_uop_fu_code,
  input  [3:0]  io_in_4_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_4_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_4_bits_uop_ctrl_op2_sel,
                io_in_4_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_4_bits_uop_ctrl_op_fcn,
  input         io_in_4_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_4_bits_uop_ctrl_csr_cmd,
  input         io_in_4_bits_uop_ctrl_is_load,
                io_in_4_bits_uop_ctrl_is_sta,
                io_in_4_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_4_bits_uop_iw_state,
  input         io_in_4_bits_uop_iw_p1_poisoned,
                io_in_4_bits_uop_iw_p2_poisoned,
                io_in_4_bits_uop_is_br,
                io_in_4_bits_uop_is_jalr,
                io_in_4_bits_uop_is_jal,
                io_in_4_bits_uop_is_sfb,
  input  [19:0] io_in_4_bits_uop_br_mask,
  input  [4:0]  io_in_4_bits_uop_br_tag,
  input  [5:0]  io_in_4_bits_uop_ftq_idx,
  input         io_in_4_bits_uop_edge_inst,
  input  [5:0]  io_in_4_bits_uop_pc_lob,
  input         io_in_4_bits_uop_taken,
  input  [19:0] io_in_4_bits_uop_imm_packed,
  input  [11:0] io_in_4_bits_uop_csr_addr,
  input  [6:0]  io_in_4_bits_uop_rob_idx,
  input  [4:0]  io_in_4_bits_uop_ldq_idx,
                io_in_4_bits_uop_stq_idx,
  input  [1:0]  io_in_4_bits_uop_rxq_idx,
  input  [6:0]  io_in_4_bits_uop_pdst,
                io_in_4_bits_uop_prs1,
                io_in_4_bits_uop_prs2,
                io_in_4_bits_uop_prs3,
  input  [5:0]  io_in_4_bits_uop_ppred,
  input         io_in_4_bits_uop_prs1_busy,
                io_in_4_bits_uop_prs2_busy,
                io_in_4_bits_uop_prs3_busy,
                io_in_4_bits_uop_ppred_busy,
  input  [6:0]  io_in_4_bits_uop_stale_pdst,
  input         io_in_4_bits_uop_exception,
  input  [63:0] io_in_4_bits_uop_exc_cause,
  input         io_in_4_bits_uop_bypassable,
  input  [4:0]  io_in_4_bits_uop_mem_cmd,
  input  [1:0]  io_in_4_bits_uop_mem_size,
  input         io_in_4_bits_uop_mem_signed,
                io_in_4_bits_uop_is_fence,
                io_in_4_bits_uop_is_fencei,
                io_in_4_bits_uop_is_amo,
                io_in_4_bits_uop_uses_ldq,
                io_in_4_bits_uop_uses_stq,
                io_in_4_bits_uop_is_sys_pc2epc,
                io_in_4_bits_uop_is_unique,
                io_in_4_bits_uop_flush_on_commit,
                io_in_4_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_4_bits_uop_ldst,
                io_in_4_bits_uop_lrs1,
                io_in_4_bits_uop_lrs2,
                io_in_4_bits_uop_lrs3,
  input         io_in_4_bits_uop_ldst_val,
  input  [1:0]  io_in_4_bits_uop_dst_rtype,
                io_in_4_bits_uop_lrs1_rtype,
                io_in_4_bits_uop_lrs2_rtype,
  input         io_in_4_bits_uop_frs3_en,
                io_in_4_bits_uop_fp_val,
                io_in_4_bits_uop_fp_single,
                io_in_4_bits_uop_xcpt_pf_if,
                io_in_4_bits_uop_xcpt_ae_if,
                io_in_4_bits_uop_xcpt_ma_if,
                io_in_4_bits_uop_bp_debug_if,
                io_in_4_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_4_bits_uop_debug_fsrc,
                io_in_4_bits_uop_debug_tsrc,
  input  [39:0] io_in_4_bits_addr,
  input         io_in_4_bits_is_hella,
  input  [7:0]  io_in_4_bits_way_en,
  input  [4:0]  io_in_4_bits_sdq_id,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [6:0]  io_in_5_bits_uop_uopc,
  input  [31:0] io_in_5_bits_uop_inst,
                io_in_5_bits_uop_debug_inst,
  input         io_in_5_bits_uop_is_rvc,
  input  [39:0] io_in_5_bits_uop_debug_pc,
  input  [2:0]  io_in_5_bits_uop_iq_type,
  input  [9:0]  io_in_5_bits_uop_fu_code,
  input  [3:0]  io_in_5_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_5_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_5_bits_uop_ctrl_op2_sel,
                io_in_5_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_5_bits_uop_ctrl_op_fcn,
  input         io_in_5_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_5_bits_uop_ctrl_csr_cmd,
  input         io_in_5_bits_uop_ctrl_is_load,
                io_in_5_bits_uop_ctrl_is_sta,
                io_in_5_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_5_bits_uop_iw_state,
  input         io_in_5_bits_uop_iw_p1_poisoned,
                io_in_5_bits_uop_iw_p2_poisoned,
                io_in_5_bits_uop_is_br,
                io_in_5_bits_uop_is_jalr,
                io_in_5_bits_uop_is_jal,
                io_in_5_bits_uop_is_sfb,
  input  [19:0] io_in_5_bits_uop_br_mask,
  input  [4:0]  io_in_5_bits_uop_br_tag,
  input  [5:0]  io_in_5_bits_uop_ftq_idx,
  input         io_in_5_bits_uop_edge_inst,
  input  [5:0]  io_in_5_bits_uop_pc_lob,
  input         io_in_5_bits_uop_taken,
  input  [19:0] io_in_5_bits_uop_imm_packed,
  input  [11:0] io_in_5_bits_uop_csr_addr,
  input  [6:0]  io_in_5_bits_uop_rob_idx,
  input  [4:0]  io_in_5_bits_uop_ldq_idx,
                io_in_5_bits_uop_stq_idx,
  input  [1:0]  io_in_5_bits_uop_rxq_idx,
  input  [6:0]  io_in_5_bits_uop_pdst,
                io_in_5_bits_uop_prs1,
                io_in_5_bits_uop_prs2,
                io_in_5_bits_uop_prs3,
  input  [5:0]  io_in_5_bits_uop_ppred,
  input         io_in_5_bits_uop_prs1_busy,
                io_in_5_bits_uop_prs2_busy,
                io_in_5_bits_uop_prs3_busy,
                io_in_5_bits_uop_ppred_busy,
  input  [6:0]  io_in_5_bits_uop_stale_pdst,
  input         io_in_5_bits_uop_exception,
  input  [63:0] io_in_5_bits_uop_exc_cause,
  input         io_in_5_bits_uop_bypassable,
  input  [4:0]  io_in_5_bits_uop_mem_cmd,
  input  [1:0]  io_in_5_bits_uop_mem_size,
  input         io_in_5_bits_uop_mem_signed,
                io_in_5_bits_uop_is_fence,
                io_in_5_bits_uop_is_fencei,
                io_in_5_bits_uop_is_amo,
                io_in_5_bits_uop_uses_ldq,
                io_in_5_bits_uop_uses_stq,
                io_in_5_bits_uop_is_sys_pc2epc,
                io_in_5_bits_uop_is_unique,
                io_in_5_bits_uop_flush_on_commit,
                io_in_5_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_5_bits_uop_ldst,
                io_in_5_bits_uop_lrs1,
                io_in_5_bits_uop_lrs2,
                io_in_5_bits_uop_lrs3,
  input         io_in_5_bits_uop_ldst_val,
  input  [1:0]  io_in_5_bits_uop_dst_rtype,
                io_in_5_bits_uop_lrs1_rtype,
                io_in_5_bits_uop_lrs2_rtype,
  input         io_in_5_bits_uop_frs3_en,
                io_in_5_bits_uop_fp_val,
                io_in_5_bits_uop_fp_single,
                io_in_5_bits_uop_xcpt_pf_if,
                io_in_5_bits_uop_xcpt_ae_if,
                io_in_5_bits_uop_xcpt_ma_if,
                io_in_5_bits_uop_bp_debug_if,
                io_in_5_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_5_bits_uop_debug_fsrc,
                io_in_5_bits_uop_debug_tsrc,
  input  [39:0] io_in_5_bits_addr,
  input         io_in_5_bits_is_hella,
  input  [7:0]  io_in_5_bits_way_en,
  input  [4:0]  io_in_5_bits_sdq_id,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [6:0]  io_in_6_bits_uop_uopc,
  input  [31:0] io_in_6_bits_uop_inst,
                io_in_6_bits_uop_debug_inst,
  input         io_in_6_bits_uop_is_rvc,
  input  [39:0] io_in_6_bits_uop_debug_pc,
  input  [2:0]  io_in_6_bits_uop_iq_type,
  input  [9:0]  io_in_6_bits_uop_fu_code,
  input  [3:0]  io_in_6_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_6_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_6_bits_uop_ctrl_op2_sel,
                io_in_6_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_6_bits_uop_ctrl_op_fcn,
  input         io_in_6_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_6_bits_uop_ctrl_csr_cmd,
  input         io_in_6_bits_uop_ctrl_is_load,
                io_in_6_bits_uop_ctrl_is_sta,
                io_in_6_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_6_bits_uop_iw_state,
  input         io_in_6_bits_uop_iw_p1_poisoned,
                io_in_6_bits_uop_iw_p2_poisoned,
                io_in_6_bits_uop_is_br,
                io_in_6_bits_uop_is_jalr,
                io_in_6_bits_uop_is_jal,
                io_in_6_bits_uop_is_sfb,
  input  [19:0] io_in_6_bits_uop_br_mask,
  input  [4:0]  io_in_6_bits_uop_br_tag,
  input  [5:0]  io_in_6_bits_uop_ftq_idx,
  input         io_in_6_bits_uop_edge_inst,
  input  [5:0]  io_in_6_bits_uop_pc_lob,
  input         io_in_6_bits_uop_taken,
  input  [19:0] io_in_6_bits_uop_imm_packed,
  input  [11:0] io_in_6_bits_uop_csr_addr,
  input  [6:0]  io_in_6_bits_uop_rob_idx,
  input  [4:0]  io_in_6_bits_uop_ldq_idx,
                io_in_6_bits_uop_stq_idx,
  input  [1:0]  io_in_6_bits_uop_rxq_idx,
  input  [6:0]  io_in_6_bits_uop_pdst,
                io_in_6_bits_uop_prs1,
                io_in_6_bits_uop_prs2,
                io_in_6_bits_uop_prs3,
  input  [5:0]  io_in_6_bits_uop_ppred,
  input         io_in_6_bits_uop_prs1_busy,
                io_in_6_bits_uop_prs2_busy,
                io_in_6_bits_uop_prs3_busy,
                io_in_6_bits_uop_ppred_busy,
  input  [6:0]  io_in_6_bits_uop_stale_pdst,
  input         io_in_6_bits_uop_exception,
  input  [63:0] io_in_6_bits_uop_exc_cause,
  input         io_in_6_bits_uop_bypassable,
  input  [4:0]  io_in_6_bits_uop_mem_cmd,
  input  [1:0]  io_in_6_bits_uop_mem_size,
  input         io_in_6_bits_uop_mem_signed,
                io_in_6_bits_uop_is_fence,
                io_in_6_bits_uop_is_fencei,
                io_in_6_bits_uop_is_amo,
                io_in_6_bits_uop_uses_ldq,
                io_in_6_bits_uop_uses_stq,
                io_in_6_bits_uop_is_sys_pc2epc,
                io_in_6_bits_uop_is_unique,
                io_in_6_bits_uop_flush_on_commit,
                io_in_6_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_6_bits_uop_ldst,
                io_in_6_bits_uop_lrs1,
                io_in_6_bits_uop_lrs2,
                io_in_6_bits_uop_lrs3,
  input         io_in_6_bits_uop_ldst_val,
  input  [1:0]  io_in_6_bits_uop_dst_rtype,
                io_in_6_bits_uop_lrs1_rtype,
                io_in_6_bits_uop_lrs2_rtype,
  input         io_in_6_bits_uop_frs3_en,
                io_in_6_bits_uop_fp_val,
                io_in_6_bits_uop_fp_single,
                io_in_6_bits_uop_xcpt_pf_if,
                io_in_6_bits_uop_xcpt_ae_if,
                io_in_6_bits_uop_xcpt_ma_if,
                io_in_6_bits_uop_bp_debug_if,
                io_in_6_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_6_bits_uop_debug_fsrc,
                io_in_6_bits_uop_debug_tsrc,
  input  [39:0] io_in_6_bits_addr,
  input         io_in_6_bits_is_hella,
  input  [7:0]  io_in_6_bits_way_en,
  input  [4:0]  io_in_6_bits_sdq_id,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [6:0]  io_in_7_bits_uop_uopc,
  input  [31:0] io_in_7_bits_uop_inst,
                io_in_7_bits_uop_debug_inst,
  input         io_in_7_bits_uop_is_rvc,
  input  [39:0] io_in_7_bits_uop_debug_pc,
  input  [2:0]  io_in_7_bits_uop_iq_type,
  input  [9:0]  io_in_7_bits_uop_fu_code,
  input  [3:0]  io_in_7_bits_uop_ctrl_br_type,
  input  [1:0]  io_in_7_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_in_7_bits_uop_ctrl_op2_sel,
                io_in_7_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_in_7_bits_uop_ctrl_op_fcn,
  input         io_in_7_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_in_7_bits_uop_ctrl_csr_cmd,
  input         io_in_7_bits_uop_ctrl_is_load,
                io_in_7_bits_uop_ctrl_is_sta,
                io_in_7_bits_uop_ctrl_is_std,
  input  [1:0]  io_in_7_bits_uop_iw_state,
  input         io_in_7_bits_uop_iw_p1_poisoned,
                io_in_7_bits_uop_iw_p2_poisoned,
                io_in_7_bits_uop_is_br,
                io_in_7_bits_uop_is_jalr,
                io_in_7_bits_uop_is_jal,
                io_in_7_bits_uop_is_sfb,
  input  [19:0] io_in_7_bits_uop_br_mask,
  input  [4:0]  io_in_7_bits_uop_br_tag,
  input  [5:0]  io_in_7_bits_uop_ftq_idx,
  input         io_in_7_bits_uop_edge_inst,
  input  [5:0]  io_in_7_bits_uop_pc_lob,
  input         io_in_7_bits_uop_taken,
  input  [19:0] io_in_7_bits_uop_imm_packed,
  input  [11:0] io_in_7_bits_uop_csr_addr,
  input  [6:0]  io_in_7_bits_uop_rob_idx,
  input  [4:0]  io_in_7_bits_uop_ldq_idx,
                io_in_7_bits_uop_stq_idx,
  input  [1:0]  io_in_7_bits_uop_rxq_idx,
  input  [6:0]  io_in_7_bits_uop_pdst,
                io_in_7_bits_uop_prs1,
                io_in_7_bits_uop_prs2,
                io_in_7_bits_uop_prs3,
  input  [5:0]  io_in_7_bits_uop_ppred,
  input         io_in_7_bits_uop_prs1_busy,
                io_in_7_bits_uop_prs2_busy,
                io_in_7_bits_uop_prs3_busy,
                io_in_7_bits_uop_ppred_busy,
  input  [6:0]  io_in_7_bits_uop_stale_pdst,
  input         io_in_7_bits_uop_exception,
  input  [63:0] io_in_7_bits_uop_exc_cause,
  input         io_in_7_bits_uop_bypassable,
  input  [4:0]  io_in_7_bits_uop_mem_cmd,
  input  [1:0]  io_in_7_bits_uop_mem_size,
  input         io_in_7_bits_uop_mem_signed,
                io_in_7_bits_uop_is_fence,
                io_in_7_bits_uop_is_fencei,
                io_in_7_bits_uop_is_amo,
                io_in_7_bits_uop_uses_ldq,
                io_in_7_bits_uop_uses_stq,
                io_in_7_bits_uop_is_sys_pc2epc,
                io_in_7_bits_uop_is_unique,
                io_in_7_bits_uop_flush_on_commit,
                io_in_7_bits_uop_ldst_is_rs1,
  input  [5:0]  io_in_7_bits_uop_ldst,
                io_in_7_bits_uop_lrs1,
                io_in_7_bits_uop_lrs2,
                io_in_7_bits_uop_lrs3,
  input         io_in_7_bits_uop_ldst_val,
  input  [1:0]  io_in_7_bits_uop_dst_rtype,
                io_in_7_bits_uop_lrs1_rtype,
                io_in_7_bits_uop_lrs2_rtype,
  input         io_in_7_bits_uop_frs3_en,
                io_in_7_bits_uop_fp_val,
                io_in_7_bits_uop_fp_single,
                io_in_7_bits_uop_xcpt_pf_if,
                io_in_7_bits_uop_xcpt_ae_if,
                io_in_7_bits_uop_xcpt_ma_if,
                io_in_7_bits_uop_bp_debug_if,
                io_in_7_bits_uop_bp_xcpt_if,
  input  [1:0]  io_in_7_bits_uop_debug_fsrc,
                io_in_7_bits_uop_debug_tsrc,
  input  [39:0] io_in_7_bits_addr,
  input         io_in_7_bits_is_hella,
  input  [7:0]  io_in_7_bits_way_en,
  input  [4:0]  io_in_7_bits_sdq_id,
  input         io_out_ready,
  output        io_out_valid,
  output [6:0]  io_out_bits_uop_uopc,
  output [31:0] io_out_bits_uop_inst,
                io_out_bits_uop_debug_inst,
  output        io_out_bits_uop_is_rvc,
  output [39:0] io_out_bits_uop_debug_pc,
  output [2:0]  io_out_bits_uop_iq_type,
  output [9:0]  io_out_bits_uop_fu_code,
  output [3:0]  io_out_bits_uop_ctrl_br_type,
  output [1:0]  io_out_bits_uop_ctrl_op1_sel,
  output [2:0]  io_out_bits_uop_ctrl_op2_sel,
                io_out_bits_uop_ctrl_imm_sel,
  output [3:0]  io_out_bits_uop_ctrl_op_fcn,
  output        io_out_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_out_bits_uop_ctrl_csr_cmd,
  output        io_out_bits_uop_ctrl_is_load,
                io_out_bits_uop_ctrl_is_sta,
                io_out_bits_uop_ctrl_is_std,
  output [1:0]  io_out_bits_uop_iw_state,
  output        io_out_bits_uop_iw_p1_poisoned,
                io_out_bits_uop_iw_p2_poisoned,
                io_out_bits_uop_is_br,
                io_out_bits_uop_is_jalr,
                io_out_bits_uop_is_jal,
                io_out_bits_uop_is_sfb,
  output [19:0] io_out_bits_uop_br_mask,
  output [4:0]  io_out_bits_uop_br_tag,
  output [5:0]  io_out_bits_uop_ftq_idx,
  output        io_out_bits_uop_edge_inst,
  output [5:0]  io_out_bits_uop_pc_lob,
  output        io_out_bits_uop_taken,
  output [19:0] io_out_bits_uop_imm_packed,
  output [11:0] io_out_bits_uop_csr_addr,
  output [6:0]  io_out_bits_uop_rob_idx,
  output [4:0]  io_out_bits_uop_ldq_idx,
                io_out_bits_uop_stq_idx,
  output [1:0]  io_out_bits_uop_rxq_idx,
  output [6:0]  io_out_bits_uop_pdst,
                io_out_bits_uop_prs1,
                io_out_bits_uop_prs2,
                io_out_bits_uop_prs3,
  output [5:0]  io_out_bits_uop_ppred,
  output        io_out_bits_uop_prs1_busy,
                io_out_bits_uop_prs2_busy,
                io_out_bits_uop_prs3_busy,
                io_out_bits_uop_ppred_busy,
  output [6:0]  io_out_bits_uop_stale_pdst,
  output        io_out_bits_uop_exception,
  output [63:0] io_out_bits_uop_exc_cause,
  output        io_out_bits_uop_bypassable,
  output [4:0]  io_out_bits_uop_mem_cmd,
  output [1:0]  io_out_bits_uop_mem_size,
  output        io_out_bits_uop_mem_signed,
                io_out_bits_uop_is_fence,
                io_out_bits_uop_is_fencei,
                io_out_bits_uop_is_amo,
                io_out_bits_uop_uses_ldq,
                io_out_bits_uop_uses_stq,
                io_out_bits_uop_is_sys_pc2epc,
                io_out_bits_uop_is_unique,
                io_out_bits_uop_flush_on_commit,
                io_out_bits_uop_ldst_is_rs1,
  output [5:0]  io_out_bits_uop_ldst,
                io_out_bits_uop_lrs1,
                io_out_bits_uop_lrs2,
                io_out_bits_uop_lrs3,
  output        io_out_bits_uop_ldst_val,
  output [1:0]  io_out_bits_uop_dst_rtype,
                io_out_bits_uop_lrs1_rtype,
                io_out_bits_uop_lrs2_rtype,
  output        io_out_bits_uop_frs3_en,
                io_out_bits_uop_fp_val,
                io_out_bits_uop_fp_single,
                io_out_bits_uop_xcpt_pf_if,
                io_out_bits_uop_xcpt_ae_if,
                io_out_bits_uop_xcpt_ma_if,
                io_out_bits_uop_bp_debug_if,
                io_out_bits_uop_bp_xcpt_if,
  output [1:0]  io_out_bits_uop_debug_fsrc,
                io_out_bits_uop_debug_tsrc,
  output [39:0] io_out_bits_addr,
  output        io_out_bits_is_hella,
  output [7:0]  io_out_bits_way_en,
  output [4:0]  io_out_bits_sdq_id
);

  wire _grant_T = io_in_0_valid | io_in_1_valid;
  wire _grant_T_1 = _grant_T | io_in_2_valid;
  wire _grant_T_2 = _grant_T_1 | io_in_3_valid;
  wire _grant_T_3 = _grant_T_2 | io_in_4_valid;
  wire _grant_T_4 = _grant_T_3 | io_in_5_valid;
  wire _io_out_valid_T = _grant_T_4 | io_in_6_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = ~io_in_0_valid & io_out_ready;
  assign io_in_2_ready = ~_grant_T & io_out_ready;
  assign io_in_3_ready = ~_grant_T_1 & io_out_ready;
  assign io_in_4_ready = ~_grant_T_2 & io_out_ready;
  assign io_in_5_ready = ~_grant_T_3 & io_out_ready;
  assign io_in_6_ready = ~_grant_T_4 & io_out_ready;
  assign io_in_7_ready = ~_io_out_valid_T & io_out_ready;
  assign io_out_valid = _io_out_valid_T | io_in_7_valid;
  assign io_out_bits_uop_uopc = io_in_0_valid ? io_in_0_bits_uop_uopc : io_in_1_valid ? io_in_1_bits_uop_uopc : io_in_2_valid ? io_in_2_bits_uop_uopc : io_in_3_valid ? io_in_3_bits_uop_uopc : io_in_4_valid ? io_in_4_bits_uop_uopc : io_in_5_valid ? io_in_5_bits_uop_uopc : io_in_6_valid ? io_in_6_bits_uop_uopc : io_in_7_bits_uop_uopc;
  assign io_out_bits_uop_inst = io_in_0_valid ? io_in_0_bits_uop_inst : io_in_1_valid ? io_in_1_bits_uop_inst : io_in_2_valid ? io_in_2_bits_uop_inst : io_in_3_valid ? io_in_3_bits_uop_inst : io_in_4_valid ? io_in_4_bits_uop_inst : io_in_5_valid ? io_in_5_bits_uop_inst : io_in_6_valid ? io_in_6_bits_uop_inst : io_in_7_bits_uop_inst;
  assign io_out_bits_uop_debug_inst = io_in_0_valid ? io_in_0_bits_uop_debug_inst : io_in_1_valid ? io_in_1_bits_uop_debug_inst : io_in_2_valid ? io_in_2_bits_uop_debug_inst : io_in_3_valid ? io_in_3_bits_uop_debug_inst : io_in_4_valid ? io_in_4_bits_uop_debug_inst : io_in_5_valid ? io_in_5_bits_uop_debug_inst : io_in_6_valid ? io_in_6_bits_uop_debug_inst : io_in_7_bits_uop_debug_inst;
  assign io_out_bits_uop_is_rvc = io_in_0_valid ? io_in_0_bits_uop_is_rvc : io_in_1_valid ? io_in_1_bits_uop_is_rvc : io_in_2_valid ? io_in_2_bits_uop_is_rvc : io_in_3_valid ? io_in_3_bits_uop_is_rvc : io_in_4_valid ? io_in_4_bits_uop_is_rvc : io_in_5_valid ? io_in_5_bits_uop_is_rvc : io_in_6_valid ? io_in_6_bits_uop_is_rvc : io_in_7_bits_uop_is_rvc;
  assign io_out_bits_uop_debug_pc = io_in_0_valid ? io_in_0_bits_uop_debug_pc : io_in_1_valid ? io_in_1_bits_uop_debug_pc : io_in_2_valid ? io_in_2_bits_uop_debug_pc : io_in_3_valid ? io_in_3_bits_uop_debug_pc : io_in_4_valid ? io_in_4_bits_uop_debug_pc : io_in_5_valid ? io_in_5_bits_uop_debug_pc : io_in_6_valid ? io_in_6_bits_uop_debug_pc : io_in_7_bits_uop_debug_pc;
  assign io_out_bits_uop_iq_type = io_in_0_valid ? io_in_0_bits_uop_iq_type : io_in_1_valid ? io_in_1_bits_uop_iq_type : io_in_2_valid ? io_in_2_bits_uop_iq_type : io_in_3_valid ? io_in_3_bits_uop_iq_type : io_in_4_valid ? io_in_4_bits_uop_iq_type : io_in_5_valid ? io_in_5_bits_uop_iq_type : io_in_6_valid ? io_in_6_bits_uop_iq_type : io_in_7_bits_uop_iq_type;
  assign io_out_bits_uop_fu_code = io_in_0_valid ? io_in_0_bits_uop_fu_code : io_in_1_valid ? io_in_1_bits_uop_fu_code : io_in_2_valid ? io_in_2_bits_uop_fu_code : io_in_3_valid ? io_in_3_bits_uop_fu_code : io_in_4_valid ? io_in_4_bits_uop_fu_code : io_in_5_valid ? io_in_5_bits_uop_fu_code : io_in_6_valid ? io_in_6_bits_uop_fu_code : io_in_7_bits_uop_fu_code;
  assign io_out_bits_uop_ctrl_br_type = io_in_0_valid ? io_in_0_bits_uop_ctrl_br_type : io_in_1_valid ? io_in_1_bits_uop_ctrl_br_type : io_in_2_valid ? io_in_2_bits_uop_ctrl_br_type : io_in_3_valid ? io_in_3_bits_uop_ctrl_br_type : io_in_4_valid ? io_in_4_bits_uop_ctrl_br_type : io_in_5_valid ? io_in_5_bits_uop_ctrl_br_type : io_in_6_valid ? io_in_6_bits_uop_ctrl_br_type : io_in_7_bits_uop_ctrl_br_type;
  assign io_out_bits_uop_ctrl_op1_sel = io_in_0_valid ? io_in_0_bits_uop_ctrl_op1_sel : io_in_1_valid ? io_in_1_bits_uop_ctrl_op1_sel : io_in_2_valid ? io_in_2_bits_uop_ctrl_op1_sel : io_in_3_valid ? io_in_3_bits_uop_ctrl_op1_sel : io_in_4_valid ? io_in_4_bits_uop_ctrl_op1_sel : io_in_5_valid ? io_in_5_bits_uop_ctrl_op1_sel : io_in_6_valid ? io_in_6_bits_uop_ctrl_op1_sel : io_in_7_bits_uop_ctrl_op1_sel;
  assign io_out_bits_uop_ctrl_op2_sel = io_in_0_valid ? io_in_0_bits_uop_ctrl_op2_sel : io_in_1_valid ? io_in_1_bits_uop_ctrl_op2_sel : io_in_2_valid ? io_in_2_bits_uop_ctrl_op2_sel : io_in_3_valid ? io_in_3_bits_uop_ctrl_op2_sel : io_in_4_valid ? io_in_4_bits_uop_ctrl_op2_sel : io_in_5_valid ? io_in_5_bits_uop_ctrl_op2_sel : io_in_6_valid ? io_in_6_bits_uop_ctrl_op2_sel : io_in_7_bits_uop_ctrl_op2_sel;
  assign io_out_bits_uop_ctrl_imm_sel = io_in_0_valid ? io_in_0_bits_uop_ctrl_imm_sel : io_in_1_valid ? io_in_1_bits_uop_ctrl_imm_sel : io_in_2_valid ? io_in_2_bits_uop_ctrl_imm_sel : io_in_3_valid ? io_in_3_bits_uop_ctrl_imm_sel : io_in_4_valid ? io_in_4_bits_uop_ctrl_imm_sel : io_in_5_valid ? io_in_5_bits_uop_ctrl_imm_sel : io_in_6_valid ? io_in_6_bits_uop_ctrl_imm_sel : io_in_7_bits_uop_ctrl_imm_sel;
  assign io_out_bits_uop_ctrl_op_fcn = io_in_0_valid ? io_in_0_bits_uop_ctrl_op_fcn : io_in_1_valid ? io_in_1_bits_uop_ctrl_op_fcn : io_in_2_valid ? io_in_2_bits_uop_ctrl_op_fcn : io_in_3_valid ? io_in_3_bits_uop_ctrl_op_fcn : io_in_4_valid ? io_in_4_bits_uop_ctrl_op_fcn : io_in_5_valid ? io_in_5_bits_uop_ctrl_op_fcn : io_in_6_valid ? io_in_6_bits_uop_ctrl_op_fcn : io_in_7_bits_uop_ctrl_op_fcn;
  assign io_out_bits_uop_ctrl_fcn_dw = io_in_0_valid ? io_in_0_bits_uop_ctrl_fcn_dw : io_in_1_valid ? io_in_1_bits_uop_ctrl_fcn_dw : io_in_2_valid ? io_in_2_bits_uop_ctrl_fcn_dw : io_in_3_valid ? io_in_3_bits_uop_ctrl_fcn_dw : io_in_4_valid ? io_in_4_bits_uop_ctrl_fcn_dw : io_in_5_valid ? io_in_5_bits_uop_ctrl_fcn_dw : io_in_6_valid ? io_in_6_bits_uop_ctrl_fcn_dw : io_in_7_bits_uop_ctrl_fcn_dw;
  assign io_out_bits_uop_ctrl_csr_cmd = io_in_0_valid ? io_in_0_bits_uop_ctrl_csr_cmd : io_in_1_valid ? io_in_1_bits_uop_ctrl_csr_cmd : io_in_2_valid ? io_in_2_bits_uop_ctrl_csr_cmd : io_in_3_valid ? io_in_3_bits_uop_ctrl_csr_cmd : io_in_4_valid ? io_in_4_bits_uop_ctrl_csr_cmd : io_in_5_valid ? io_in_5_bits_uop_ctrl_csr_cmd : io_in_6_valid ? io_in_6_bits_uop_ctrl_csr_cmd : io_in_7_bits_uop_ctrl_csr_cmd;
  assign io_out_bits_uop_ctrl_is_load = io_in_0_valid ? io_in_0_bits_uop_ctrl_is_load : io_in_1_valid ? io_in_1_bits_uop_ctrl_is_load : io_in_2_valid ? io_in_2_bits_uop_ctrl_is_load : io_in_3_valid ? io_in_3_bits_uop_ctrl_is_load : io_in_4_valid ? io_in_4_bits_uop_ctrl_is_load : io_in_5_valid ? io_in_5_bits_uop_ctrl_is_load : io_in_6_valid ? io_in_6_bits_uop_ctrl_is_load : io_in_7_bits_uop_ctrl_is_load;
  assign io_out_bits_uop_ctrl_is_sta = io_in_0_valid ? io_in_0_bits_uop_ctrl_is_sta : io_in_1_valid ? io_in_1_bits_uop_ctrl_is_sta : io_in_2_valid ? io_in_2_bits_uop_ctrl_is_sta : io_in_3_valid ? io_in_3_bits_uop_ctrl_is_sta : io_in_4_valid ? io_in_4_bits_uop_ctrl_is_sta : io_in_5_valid ? io_in_5_bits_uop_ctrl_is_sta : io_in_6_valid ? io_in_6_bits_uop_ctrl_is_sta : io_in_7_bits_uop_ctrl_is_sta;
  assign io_out_bits_uop_ctrl_is_std = io_in_0_valid ? io_in_0_bits_uop_ctrl_is_std : io_in_1_valid ? io_in_1_bits_uop_ctrl_is_std : io_in_2_valid ? io_in_2_bits_uop_ctrl_is_std : io_in_3_valid ? io_in_3_bits_uop_ctrl_is_std : io_in_4_valid ? io_in_4_bits_uop_ctrl_is_std : io_in_5_valid ? io_in_5_bits_uop_ctrl_is_std : io_in_6_valid ? io_in_6_bits_uop_ctrl_is_std : io_in_7_bits_uop_ctrl_is_std;
  assign io_out_bits_uop_iw_state = io_in_0_valid ? io_in_0_bits_uop_iw_state : io_in_1_valid ? io_in_1_bits_uop_iw_state : io_in_2_valid ? io_in_2_bits_uop_iw_state : io_in_3_valid ? io_in_3_bits_uop_iw_state : io_in_4_valid ? io_in_4_bits_uop_iw_state : io_in_5_valid ? io_in_5_bits_uop_iw_state : io_in_6_valid ? io_in_6_bits_uop_iw_state : io_in_7_bits_uop_iw_state;
  assign io_out_bits_uop_iw_p1_poisoned = io_in_0_valid ? io_in_0_bits_uop_iw_p1_poisoned : io_in_1_valid ? io_in_1_bits_uop_iw_p1_poisoned : io_in_2_valid ? io_in_2_bits_uop_iw_p1_poisoned : io_in_3_valid ? io_in_3_bits_uop_iw_p1_poisoned : io_in_4_valid ? io_in_4_bits_uop_iw_p1_poisoned : io_in_5_valid ? io_in_5_bits_uop_iw_p1_poisoned : io_in_6_valid ? io_in_6_bits_uop_iw_p1_poisoned : io_in_7_bits_uop_iw_p1_poisoned;
  assign io_out_bits_uop_iw_p2_poisoned = io_in_0_valid ? io_in_0_bits_uop_iw_p2_poisoned : io_in_1_valid ? io_in_1_bits_uop_iw_p2_poisoned : io_in_2_valid ? io_in_2_bits_uop_iw_p2_poisoned : io_in_3_valid ? io_in_3_bits_uop_iw_p2_poisoned : io_in_4_valid ? io_in_4_bits_uop_iw_p2_poisoned : io_in_5_valid ? io_in_5_bits_uop_iw_p2_poisoned : io_in_6_valid ? io_in_6_bits_uop_iw_p2_poisoned : io_in_7_bits_uop_iw_p2_poisoned;
  assign io_out_bits_uop_is_br = io_in_0_valid ? io_in_0_bits_uop_is_br : io_in_1_valid ? io_in_1_bits_uop_is_br : io_in_2_valid ? io_in_2_bits_uop_is_br : io_in_3_valid ? io_in_3_bits_uop_is_br : io_in_4_valid ? io_in_4_bits_uop_is_br : io_in_5_valid ? io_in_5_bits_uop_is_br : io_in_6_valid ? io_in_6_bits_uop_is_br : io_in_7_bits_uop_is_br;
  assign io_out_bits_uop_is_jalr = io_in_0_valid ? io_in_0_bits_uop_is_jalr : io_in_1_valid ? io_in_1_bits_uop_is_jalr : io_in_2_valid ? io_in_2_bits_uop_is_jalr : io_in_3_valid ? io_in_3_bits_uop_is_jalr : io_in_4_valid ? io_in_4_bits_uop_is_jalr : io_in_5_valid ? io_in_5_bits_uop_is_jalr : io_in_6_valid ? io_in_6_bits_uop_is_jalr : io_in_7_bits_uop_is_jalr;
  assign io_out_bits_uop_is_jal = io_in_0_valid ? io_in_0_bits_uop_is_jal : io_in_1_valid ? io_in_1_bits_uop_is_jal : io_in_2_valid ? io_in_2_bits_uop_is_jal : io_in_3_valid ? io_in_3_bits_uop_is_jal : io_in_4_valid ? io_in_4_bits_uop_is_jal : io_in_5_valid ? io_in_5_bits_uop_is_jal : io_in_6_valid ? io_in_6_bits_uop_is_jal : io_in_7_bits_uop_is_jal;
  assign io_out_bits_uop_is_sfb = io_in_0_valid ? io_in_0_bits_uop_is_sfb : io_in_1_valid ? io_in_1_bits_uop_is_sfb : io_in_2_valid ? io_in_2_bits_uop_is_sfb : io_in_3_valid ? io_in_3_bits_uop_is_sfb : io_in_4_valid ? io_in_4_bits_uop_is_sfb : io_in_5_valid ? io_in_5_bits_uop_is_sfb : io_in_6_valid ? io_in_6_bits_uop_is_sfb : io_in_7_bits_uop_is_sfb;
  assign io_out_bits_uop_br_mask = io_in_0_valid ? io_in_0_bits_uop_br_mask : io_in_1_valid ? io_in_1_bits_uop_br_mask : io_in_2_valid ? io_in_2_bits_uop_br_mask : io_in_3_valid ? io_in_3_bits_uop_br_mask : io_in_4_valid ? io_in_4_bits_uop_br_mask : io_in_5_valid ? io_in_5_bits_uop_br_mask : io_in_6_valid ? io_in_6_bits_uop_br_mask : io_in_7_bits_uop_br_mask;
  assign io_out_bits_uop_br_tag = io_in_0_valid ? io_in_0_bits_uop_br_tag : io_in_1_valid ? io_in_1_bits_uop_br_tag : io_in_2_valid ? io_in_2_bits_uop_br_tag : io_in_3_valid ? io_in_3_bits_uop_br_tag : io_in_4_valid ? io_in_4_bits_uop_br_tag : io_in_5_valid ? io_in_5_bits_uop_br_tag : io_in_6_valid ? io_in_6_bits_uop_br_tag : io_in_7_bits_uop_br_tag;
  assign io_out_bits_uop_ftq_idx = io_in_0_valid ? io_in_0_bits_uop_ftq_idx : io_in_1_valid ? io_in_1_bits_uop_ftq_idx : io_in_2_valid ? io_in_2_bits_uop_ftq_idx : io_in_3_valid ? io_in_3_bits_uop_ftq_idx : io_in_4_valid ? io_in_4_bits_uop_ftq_idx : io_in_5_valid ? io_in_5_bits_uop_ftq_idx : io_in_6_valid ? io_in_6_bits_uop_ftq_idx : io_in_7_bits_uop_ftq_idx;
  assign io_out_bits_uop_edge_inst = io_in_0_valid ? io_in_0_bits_uop_edge_inst : io_in_1_valid ? io_in_1_bits_uop_edge_inst : io_in_2_valid ? io_in_2_bits_uop_edge_inst : io_in_3_valid ? io_in_3_bits_uop_edge_inst : io_in_4_valid ? io_in_4_bits_uop_edge_inst : io_in_5_valid ? io_in_5_bits_uop_edge_inst : io_in_6_valid ? io_in_6_bits_uop_edge_inst : io_in_7_bits_uop_edge_inst;
  assign io_out_bits_uop_pc_lob = io_in_0_valid ? io_in_0_bits_uop_pc_lob : io_in_1_valid ? io_in_1_bits_uop_pc_lob : io_in_2_valid ? io_in_2_bits_uop_pc_lob : io_in_3_valid ? io_in_3_bits_uop_pc_lob : io_in_4_valid ? io_in_4_bits_uop_pc_lob : io_in_5_valid ? io_in_5_bits_uop_pc_lob : io_in_6_valid ? io_in_6_bits_uop_pc_lob : io_in_7_bits_uop_pc_lob;
  assign io_out_bits_uop_taken = io_in_0_valid ? io_in_0_bits_uop_taken : io_in_1_valid ? io_in_1_bits_uop_taken : io_in_2_valid ? io_in_2_bits_uop_taken : io_in_3_valid ? io_in_3_bits_uop_taken : io_in_4_valid ? io_in_4_bits_uop_taken : io_in_5_valid ? io_in_5_bits_uop_taken : io_in_6_valid ? io_in_6_bits_uop_taken : io_in_7_bits_uop_taken;
  assign io_out_bits_uop_imm_packed = io_in_0_valid ? io_in_0_bits_uop_imm_packed : io_in_1_valid ? io_in_1_bits_uop_imm_packed : io_in_2_valid ? io_in_2_bits_uop_imm_packed : io_in_3_valid ? io_in_3_bits_uop_imm_packed : io_in_4_valid ? io_in_4_bits_uop_imm_packed : io_in_5_valid ? io_in_5_bits_uop_imm_packed : io_in_6_valid ? io_in_6_bits_uop_imm_packed : io_in_7_bits_uop_imm_packed;
  assign io_out_bits_uop_csr_addr = io_in_0_valid ? io_in_0_bits_uop_csr_addr : io_in_1_valid ? io_in_1_bits_uop_csr_addr : io_in_2_valid ? io_in_2_bits_uop_csr_addr : io_in_3_valid ? io_in_3_bits_uop_csr_addr : io_in_4_valid ? io_in_4_bits_uop_csr_addr : io_in_5_valid ? io_in_5_bits_uop_csr_addr : io_in_6_valid ? io_in_6_bits_uop_csr_addr : io_in_7_bits_uop_csr_addr;
  assign io_out_bits_uop_rob_idx = io_in_0_valid ? io_in_0_bits_uop_rob_idx : io_in_1_valid ? io_in_1_bits_uop_rob_idx : io_in_2_valid ? io_in_2_bits_uop_rob_idx : io_in_3_valid ? io_in_3_bits_uop_rob_idx : io_in_4_valid ? io_in_4_bits_uop_rob_idx : io_in_5_valid ? io_in_5_bits_uop_rob_idx : io_in_6_valid ? io_in_6_bits_uop_rob_idx : io_in_7_bits_uop_rob_idx;
  assign io_out_bits_uop_ldq_idx = io_in_0_valid ? io_in_0_bits_uop_ldq_idx : io_in_1_valid ? io_in_1_bits_uop_ldq_idx : io_in_2_valid ? io_in_2_bits_uop_ldq_idx : io_in_3_valid ? io_in_3_bits_uop_ldq_idx : io_in_4_valid ? io_in_4_bits_uop_ldq_idx : io_in_5_valid ? io_in_5_bits_uop_ldq_idx : io_in_6_valid ? io_in_6_bits_uop_ldq_idx : io_in_7_bits_uop_ldq_idx;
  assign io_out_bits_uop_stq_idx = io_in_0_valid ? io_in_0_bits_uop_stq_idx : io_in_1_valid ? io_in_1_bits_uop_stq_idx : io_in_2_valid ? io_in_2_bits_uop_stq_idx : io_in_3_valid ? io_in_3_bits_uop_stq_idx : io_in_4_valid ? io_in_4_bits_uop_stq_idx : io_in_5_valid ? io_in_5_bits_uop_stq_idx : io_in_6_valid ? io_in_6_bits_uop_stq_idx : io_in_7_bits_uop_stq_idx;
  assign io_out_bits_uop_rxq_idx = io_in_0_valid ? io_in_0_bits_uop_rxq_idx : io_in_1_valid ? io_in_1_bits_uop_rxq_idx : io_in_2_valid ? io_in_2_bits_uop_rxq_idx : io_in_3_valid ? io_in_3_bits_uop_rxq_idx : io_in_4_valid ? io_in_4_bits_uop_rxq_idx : io_in_5_valid ? io_in_5_bits_uop_rxq_idx : io_in_6_valid ? io_in_6_bits_uop_rxq_idx : io_in_7_bits_uop_rxq_idx;
  assign io_out_bits_uop_pdst = io_in_0_valid ? io_in_0_bits_uop_pdst : io_in_1_valid ? io_in_1_bits_uop_pdst : io_in_2_valid ? io_in_2_bits_uop_pdst : io_in_3_valid ? io_in_3_bits_uop_pdst : io_in_4_valid ? io_in_4_bits_uop_pdst : io_in_5_valid ? io_in_5_bits_uop_pdst : io_in_6_valid ? io_in_6_bits_uop_pdst : io_in_7_bits_uop_pdst;
  assign io_out_bits_uop_prs1 = io_in_0_valid ? io_in_0_bits_uop_prs1 : io_in_1_valid ? io_in_1_bits_uop_prs1 : io_in_2_valid ? io_in_2_bits_uop_prs1 : io_in_3_valid ? io_in_3_bits_uop_prs1 : io_in_4_valid ? io_in_4_bits_uop_prs1 : io_in_5_valid ? io_in_5_bits_uop_prs1 : io_in_6_valid ? io_in_6_bits_uop_prs1 : io_in_7_bits_uop_prs1;
  assign io_out_bits_uop_prs2 = io_in_0_valid ? io_in_0_bits_uop_prs2 : io_in_1_valid ? io_in_1_bits_uop_prs2 : io_in_2_valid ? io_in_2_bits_uop_prs2 : io_in_3_valid ? io_in_3_bits_uop_prs2 : io_in_4_valid ? io_in_4_bits_uop_prs2 : io_in_5_valid ? io_in_5_bits_uop_prs2 : io_in_6_valid ? io_in_6_bits_uop_prs2 : io_in_7_bits_uop_prs2;
  assign io_out_bits_uop_prs3 = io_in_0_valid ? io_in_0_bits_uop_prs3 : io_in_1_valid ? io_in_1_bits_uop_prs3 : io_in_2_valid ? io_in_2_bits_uop_prs3 : io_in_3_valid ? io_in_3_bits_uop_prs3 : io_in_4_valid ? io_in_4_bits_uop_prs3 : io_in_5_valid ? io_in_5_bits_uop_prs3 : io_in_6_valid ? io_in_6_bits_uop_prs3 : io_in_7_bits_uop_prs3;
  assign io_out_bits_uop_ppred = io_in_0_valid ? io_in_0_bits_uop_ppred : io_in_1_valid ? io_in_1_bits_uop_ppred : io_in_2_valid ? io_in_2_bits_uop_ppred : io_in_3_valid ? io_in_3_bits_uop_ppred : io_in_4_valid ? io_in_4_bits_uop_ppred : io_in_5_valid ? io_in_5_bits_uop_ppred : io_in_6_valid ? io_in_6_bits_uop_ppred : io_in_7_bits_uop_ppred;
  assign io_out_bits_uop_prs1_busy = io_in_0_valid ? io_in_0_bits_uop_prs1_busy : io_in_1_valid ? io_in_1_bits_uop_prs1_busy : io_in_2_valid ? io_in_2_bits_uop_prs1_busy : io_in_3_valid ? io_in_3_bits_uop_prs1_busy : io_in_4_valid ? io_in_4_bits_uop_prs1_busy : io_in_5_valid ? io_in_5_bits_uop_prs1_busy : io_in_6_valid ? io_in_6_bits_uop_prs1_busy : io_in_7_bits_uop_prs1_busy;
  assign io_out_bits_uop_prs2_busy = io_in_0_valid ? io_in_0_bits_uop_prs2_busy : io_in_1_valid ? io_in_1_bits_uop_prs2_busy : io_in_2_valid ? io_in_2_bits_uop_prs2_busy : io_in_3_valid ? io_in_3_bits_uop_prs2_busy : io_in_4_valid ? io_in_4_bits_uop_prs2_busy : io_in_5_valid ? io_in_5_bits_uop_prs2_busy : io_in_6_valid ? io_in_6_bits_uop_prs2_busy : io_in_7_bits_uop_prs2_busy;
  assign io_out_bits_uop_prs3_busy = io_in_0_valid ? io_in_0_bits_uop_prs3_busy : io_in_1_valid ? io_in_1_bits_uop_prs3_busy : io_in_2_valid ? io_in_2_bits_uop_prs3_busy : io_in_3_valid ? io_in_3_bits_uop_prs3_busy : io_in_4_valid ? io_in_4_bits_uop_prs3_busy : io_in_5_valid ? io_in_5_bits_uop_prs3_busy : io_in_6_valid ? io_in_6_bits_uop_prs3_busy : io_in_7_bits_uop_prs3_busy;
  assign io_out_bits_uop_ppred_busy = io_in_0_valid ? io_in_0_bits_uop_ppred_busy : io_in_1_valid ? io_in_1_bits_uop_ppred_busy : io_in_2_valid ? io_in_2_bits_uop_ppred_busy : io_in_3_valid ? io_in_3_bits_uop_ppred_busy : io_in_4_valid ? io_in_4_bits_uop_ppred_busy : io_in_5_valid ? io_in_5_bits_uop_ppred_busy : io_in_6_valid ? io_in_6_bits_uop_ppred_busy : io_in_7_bits_uop_ppred_busy;
  assign io_out_bits_uop_stale_pdst = io_in_0_valid ? io_in_0_bits_uop_stale_pdst : io_in_1_valid ? io_in_1_bits_uop_stale_pdst : io_in_2_valid ? io_in_2_bits_uop_stale_pdst : io_in_3_valid ? io_in_3_bits_uop_stale_pdst : io_in_4_valid ? io_in_4_bits_uop_stale_pdst : io_in_5_valid ? io_in_5_bits_uop_stale_pdst : io_in_6_valid ? io_in_6_bits_uop_stale_pdst : io_in_7_bits_uop_stale_pdst;
  assign io_out_bits_uop_exception = io_in_0_valid ? io_in_0_bits_uop_exception : io_in_1_valid ? io_in_1_bits_uop_exception : io_in_2_valid ? io_in_2_bits_uop_exception : io_in_3_valid ? io_in_3_bits_uop_exception : io_in_4_valid ? io_in_4_bits_uop_exception : io_in_5_valid ? io_in_5_bits_uop_exception : io_in_6_valid ? io_in_6_bits_uop_exception : io_in_7_bits_uop_exception;
  assign io_out_bits_uop_exc_cause = io_in_0_valid ? io_in_0_bits_uop_exc_cause : io_in_1_valid ? io_in_1_bits_uop_exc_cause : io_in_2_valid ? io_in_2_bits_uop_exc_cause : io_in_3_valid ? io_in_3_bits_uop_exc_cause : io_in_4_valid ? io_in_4_bits_uop_exc_cause : io_in_5_valid ? io_in_5_bits_uop_exc_cause : io_in_6_valid ? io_in_6_bits_uop_exc_cause : io_in_7_bits_uop_exc_cause;
  assign io_out_bits_uop_bypassable = io_in_0_valid ? io_in_0_bits_uop_bypassable : io_in_1_valid ? io_in_1_bits_uop_bypassable : io_in_2_valid ? io_in_2_bits_uop_bypassable : io_in_3_valid ? io_in_3_bits_uop_bypassable : io_in_4_valid ? io_in_4_bits_uop_bypassable : io_in_5_valid ? io_in_5_bits_uop_bypassable : io_in_6_valid ? io_in_6_bits_uop_bypassable : io_in_7_bits_uop_bypassable;
  assign io_out_bits_uop_mem_cmd = io_in_0_valid ? io_in_0_bits_uop_mem_cmd : io_in_1_valid ? io_in_1_bits_uop_mem_cmd : io_in_2_valid ? io_in_2_bits_uop_mem_cmd : io_in_3_valid ? io_in_3_bits_uop_mem_cmd : io_in_4_valid ? io_in_4_bits_uop_mem_cmd : io_in_5_valid ? io_in_5_bits_uop_mem_cmd : io_in_6_valid ? io_in_6_bits_uop_mem_cmd : io_in_7_bits_uop_mem_cmd;
  assign io_out_bits_uop_mem_size = io_in_0_valid ? io_in_0_bits_uop_mem_size : io_in_1_valid ? io_in_1_bits_uop_mem_size : io_in_2_valid ? io_in_2_bits_uop_mem_size : io_in_3_valid ? io_in_3_bits_uop_mem_size : io_in_4_valid ? io_in_4_bits_uop_mem_size : io_in_5_valid ? io_in_5_bits_uop_mem_size : io_in_6_valid ? io_in_6_bits_uop_mem_size : io_in_7_bits_uop_mem_size;
  assign io_out_bits_uop_mem_signed = io_in_0_valid ? io_in_0_bits_uop_mem_signed : io_in_1_valid ? io_in_1_bits_uop_mem_signed : io_in_2_valid ? io_in_2_bits_uop_mem_signed : io_in_3_valid ? io_in_3_bits_uop_mem_signed : io_in_4_valid ? io_in_4_bits_uop_mem_signed : io_in_5_valid ? io_in_5_bits_uop_mem_signed : io_in_6_valid ? io_in_6_bits_uop_mem_signed : io_in_7_bits_uop_mem_signed;
  assign io_out_bits_uop_is_fence = io_in_0_valid ? io_in_0_bits_uop_is_fence : io_in_1_valid ? io_in_1_bits_uop_is_fence : io_in_2_valid ? io_in_2_bits_uop_is_fence : io_in_3_valid ? io_in_3_bits_uop_is_fence : io_in_4_valid ? io_in_4_bits_uop_is_fence : io_in_5_valid ? io_in_5_bits_uop_is_fence : io_in_6_valid ? io_in_6_bits_uop_is_fence : io_in_7_bits_uop_is_fence;
  assign io_out_bits_uop_is_fencei = io_in_0_valid ? io_in_0_bits_uop_is_fencei : io_in_1_valid ? io_in_1_bits_uop_is_fencei : io_in_2_valid ? io_in_2_bits_uop_is_fencei : io_in_3_valid ? io_in_3_bits_uop_is_fencei : io_in_4_valid ? io_in_4_bits_uop_is_fencei : io_in_5_valid ? io_in_5_bits_uop_is_fencei : io_in_6_valid ? io_in_6_bits_uop_is_fencei : io_in_7_bits_uop_is_fencei;
  assign io_out_bits_uop_is_amo = io_in_0_valid ? io_in_0_bits_uop_is_amo : io_in_1_valid ? io_in_1_bits_uop_is_amo : io_in_2_valid ? io_in_2_bits_uop_is_amo : io_in_3_valid ? io_in_3_bits_uop_is_amo : io_in_4_valid ? io_in_4_bits_uop_is_amo : io_in_5_valid ? io_in_5_bits_uop_is_amo : io_in_6_valid ? io_in_6_bits_uop_is_amo : io_in_7_bits_uop_is_amo;
  assign io_out_bits_uop_uses_ldq = io_in_0_valid ? io_in_0_bits_uop_uses_ldq : io_in_1_valid ? io_in_1_bits_uop_uses_ldq : io_in_2_valid ? io_in_2_bits_uop_uses_ldq : io_in_3_valid ? io_in_3_bits_uop_uses_ldq : io_in_4_valid ? io_in_4_bits_uop_uses_ldq : io_in_5_valid ? io_in_5_bits_uop_uses_ldq : io_in_6_valid ? io_in_6_bits_uop_uses_ldq : io_in_7_bits_uop_uses_ldq;
  assign io_out_bits_uop_uses_stq = io_in_0_valid ? io_in_0_bits_uop_uses_stq : io_in_1_valid ? io_in_1_bits_uop_uses_stq : io_in_2_valid ? io_in_2_bits_uop_uses_stq : io_in_3_valid ? io_in_3_bits_uop_uses_stq : io_in_4_valid ? io_in_4_bits_uop_uses_stq : io_in_5_valid ? io_in_5_bits_uop_uses_stq : io_in_6_valid ? io_in_6_bits_uop_uses_stq : io_in_7_bits_uop_uses_stq;
  assign io_out_bits_uop_is_sys_pc2epc = io_in_0_valid ? io_in_0_bits_uop_is_sys_pc2epc : io_in_1_valid ? io_in_1_bits_uop_is_sys_pc2epc : io_in_2_valid ? io_in_2_bits_uop_is_sys_pc2epc : io_in_3_valid ? io_in_3_bits_uop_is_sys_pc2epc : io_in_4_valid ? io_in_4_bits_uop_is_sys_pc2epc : io_in_5_valid ? io_in_5_bits_uop_is_sys_pc2epc : io_in_6_valid ? io_in_6_bits_uop_is_sys_pc2epc : io_in_7_bits_uop_is_sys_pc2epc;
  assign io_out_bits_uop_is_unique = io_in_0_valid ? io_in_0_bits_uop_is_unique : io_in_1_valid ? io_in_1_bits_uop_is_unique : io_in_2_valid ? io_in_2_bits_uop_is_unique : io_in_3_valid ? io_in_3_bits_uop_is_unique : io_in_4_valid ? io_in_4_bits_uop_is_unique : io_in_5_valid ? io_in_5_bits_uop_is_unique : io_in_6_valid ? io_in_6_bits_uop_is_unique : io_in_7_bits_uop_is_unique;
  assign io_out_bits_uop_flush_on_commit = io_in_0_valid ? io_in_0_bits_uop_flush_on_commit : io_in_1_valid ? io_in_1_bits_uop_flush_on_commit : io_in_2_valid ? io_in_2_bits_uop_flush_on_commit : io_in_3_valid ? io_in_3_bits_uop_flush_on_commit : io_in_4_valid ? io_in_4_bits_uop_flush_on_commit : io_in_5_valid ? io_in_5_bits_uop_flush_on_commit : io_in_6_valid ? io_in_6_bits_uop_flush_on_commit : io_in_7_bits_uop_flush_on_commit;
  assign io_out_bits_uop_ldst_is_rs1 = io_in_0_valid ? io_in_0_bits_uop_ldst_is_rs1 : io_in_1_valid ? io_in_1_bits_uop_ldst_is_rs1 : io_in_2_valid ? io_in_2_bits_uop_ldst_is_rs1 : io_in_3_valid ? io_in_3_bits_uop_ldst_is_rs1 : io_in_4_valid ? io_in_4_bits_uop_ldst_is_rs1 : io_in_5_valid ? io_in_5_bits_uop_ldst_is_rs1 : io_in_6_valid ? io_in_6_bits_uop_ldst_is_rs1 : io_in_7_bits_uop_ldst_is_rs1;
  assign io_out_bits_uop_ldst = io_in_0_valid ? io_in_0_bits_uop_ldst : io_in_1_valid ? io_in_1_bits_uop_ldst : io_in_2_valid ? io_in_2_bits_uop_ldst : io_in_3_valid ? io_in_3_bits_uop_ldst : io_in_4_valid ? io_in_4_bits_uop_ldst : io_in_5_valid ? io_in_5_bits_uop_ldst : io_in_6_valid ? io_in_6_bits_uop_ldst : io_in_7_bits_uop_ldst;
  assign io_out_bits_uop_lrs1 = io_in_0_valid ? io_in_0_bits_uop_lrs1 : io_in_1_valid ? io_in_1_bits_uop_lrs1 : io_in_2_valid ? io_in_2_bits_uop_lrs1 : io_in_3_valid ? io_in_3_bits_uop_lrs1 : io_in_4_valid ? io_in_4_bits_uop_lrs1 : io_in_5_valid ? io_in_5_bits_uop_lrs1 : io_in_6_valid ? io_in_6_bits_uop_lrs1 : io_in_7_bits_uop_lrs1;
  assign io_out_bits_uop_lrs2 = io_in_0_valid ? io_in_0_bits_uop_lrs2 : io_in_1_valid ? io_in_1_bits_uop_lrs2 : io_in_2_valid ? io_in_2_bits_uop_lrs2 : io_in_3_valid ? io_in_3_bits_uop_lrs2 : io_in_4_valid ? io_in_4_bits_uop_lrs2 : io_in_5_valid ? io_in_5_bits_uop_lrs2 : io_in_6_valid ? io_in_6_bits_uop_lrs2 : io_in_7_bits_uop_lrs2;
  assign io_out_bits_uop_lrs3 = io_in_0_valid ? io_in_0_bits_uop_lrs3 : io_in_1_valid ? io_in_1_bits_uop_lrs3 : io_in_2_valid ? io_in_2_bits_uop_lrs3 : io_in_3_valid ? io_in_3_bits_uop_lrs3 : io_in_4_valid ? io_in_4_bits_uop_lrs3 : io_in_5_valid ? io_in_5_bits_uop_lrs3 : io_in_6_valid ? io_in_6_bits_uop_lrs3 : io_in_7_bits_uop_lrs3;
  assign io_out_bits_uop_ldst_val = io_in_0_valid ? io_in_0_bits_uop_ldst_val : io_in_1_valid ? io_in_1_bits_uop_ldst_val : io_in_2_valid ? io_in_2_bits_uop_ldst_val : io_in_3_valid ? io_in_3_bits_uop_ldst_val : io_in_4_valid ? io_in_4_bits_uop_ldst_val : io_in_5_valid ? io_in_5_bits_uop_ldst_val : io_in_6_valid ? io_in_6_bits_uop_ldst_val : io_in_7_bits_uop_ldst_val;
  assign io_out_bits_uop_dst_rtype = io_in_0_valid ? io_in_0_bits_uop_dst_rtype : io_in_1_valid ? io_in_1_bits_uop_dst_rtype : io_in_2_valid ? io_in_2_bits_uop_dst_rtype : io_in_3_valid ? io_in_3_bits_uop_dst_rtype : io_in_4_valid ? io_in_4_bits_uop_dst_rtype : io_in_5_valid ? io_in_5_bits_uop_dst_rtype : io_in_6_valid ? io_in_6_bits_uop_dst_rtype : io_in_7_bits_uop_dst_rtype;
  assign io_out_bits_uop_lrs1_rtype = io_in_0_valid ? io_in_0_bits_uop_lrs1_rtype : io_in_1_valid ? io_in_1_bits_uop_lrs1_rtype : io_in_2_valid ? io_in_2_bits_uop_lrs1_rtype : io_in_3_valid ? io_in_3_bits_uop_lrs1_rtype : io_in_4_valid ? io_in_4_bits_uop_lrs1_rtype : io_in_5_valid ? io_in_5_bits_uop_lrs1_rtype : io_in_6_valid ? io_in_6_bits_uop_lrs1_rtype : io_in_7_bits_uop_lrs1_rtype;
  assign io_out_bits_uop_lrs2_rtype = io_in_0_valid ? io_in_0_bits_uop_lrs2_rtype : io_in_1_valid ? io_in_1_bits_uop_lrs2_rtype : io_in_2_valid ? io_in_2_bits_uop_lrs2_rtype : io_in_3_valid ? io_in_3_bits_uop_lrs2_rtype : io_in_4_valid ? io_in_4_bits_uop_lrs2_rtype : io_in_5_valid ? io_in_5_bits_uop_lrs2_rtype : io_in_6_valid ? io_in_6_bits_uop_lrs2_rtype : io_in_7_bits_uop_lrs2_rtype;
  assign io_out_bits_uop_frs3_en = io_in_0_valid ? io_in_0_bits_uop_frs3_en : io_in_1_valid ? io_in_1_bits_uop_frs3_en : io_in_2_valid ? io_in_2_bits_uop_frs3_en : io_in_3_valid ? io_in_3_bits_uop_frs3_en : io_in_4_valid ? io_in_4_bits_uop_frs3_en : io_in_5_valid ? io_in_5_bits_uop_frs3_en : io_in_6_valid ? io_in_6_bits_uop_frs3_en : io_in_7_bits_uop_frs3_en;
  assign io_out_bits_uop_fp_val = io_in_0_valid ? io_in_0_bits_uop_fp_val : io_in_1_valid ? io_in_1_bits_uop_fp_val : io_in_2_valid ? io_in_2_bits_uop_fp_val : io_in_3_valid ? io_in_3_bits_uop_fp_val : io_in_4_valid ? io_in_4_bits_uop_fp_val : io_in_5_valid ? io_in_5_bits_uop_fp_val : io_in_6_valid ? io_in_6_bits_uop_fp_val : io_in_7_bits_uop_fp_val;
  assign io_out_bits_uop_fp_single = io_in_0_valid ? io_in_0_bits_uop_fp_single : io_in_1_valid ? io_in_1_bits_uop_fp_single : io_in_2_valid ? io_in_2_bits_uop_fp_single : io_in_3_valid ? io_in_3_bits_uop_fp_single : io_in_4_valid ? io_in_4_bits_uop_fp_single : io_in_5_valid ? io_in_5_bits_uop_fp_single : io_in_6_valid ? io_in_6_bits_uop_fp_single : io_in_7_bits_uop_fp_single;
  assign io_out_bits_uop_xcpt_pf_if = io_in_0_valid ? io_in_0_bits_uop_xcpt_pf_if : io_in_1_valid ? io_in_1_bits_uop_xcpt_pf_if : io_in_2_valid ? io_in_2_bits_uop_xcpt_pf_if : io_in_3_valid ? io_in_3_bits_uop_xcpt_pf_if : io_in_4_valid ? io_in_4_bits_uop_xcpt_pf_if : io_in_5_valid ? io_in_5_bits_uop_xcpt_pf_if : io_in_6_valid ? io_in_6_bits_uop_xcpt_pf_if : io_in_7_bits_uop_xcpt_pf_if;
  assign io_out_bits_uop_xcpt_ae_if = io_in_0_valid ? io_in_0_bits_uop_xcpt_ae_if : io_in_1_valid ? io_in_1_bits_uop_xcpt_ae_if : io_in_2_valid ? io_in_2_bits_uop_xcpt_ae_if : io_in_3_valid ? io_in_3_bits_uop_xcpt_ae_if : io_in_4_valid ? io_in_4_bits_uop_xcpt_ae_if : io_in_5_valid ? io_in_5_bits_uop_xcpt_ae_if : io_in_6_valid ? io_in_6_bits_uop_xcpt_ae_if : io_in_7_bits_uop_xcpt_ae_if;
  assign io_out_bits_uop_xcpt_ma_if = io_in_0_valid ? io_in_0_bits_uop_xcpt_ma_if : io_in_1_valid ? io_in_1_bits_uop_xcpt_ma_if : io_in_2_valid ? io_in_2_bits_uop_xcpt_ma_if : io_in_3_valid ? io_in_3_bits_uop_xcpt_ma_if : io_in_4_valid ? io_in_4_bits_uop_xcpt_ma_if : io_in_5_valid ? io_in_5_bits_uop_xcpt_ma_if : io_in_6_valid ? io_in_6_bits_uop_xcpt_ma_if : io_in_7_bits_uop_xcpt_ma_if;
  assign io_out_bits_uop_bp_debug_if = io_in_0_valid ? io_in_0_bits_uop_bp_debug_if : io_in_1_valid ? io_in_1_bits_uop_bp_debug_if : io_in_2_valid ? io_in_2_bits_uop_bp_debug_if : io_in_3_valid ? io_in_3_bits_uop_bp_debug_if : io_in_4_valid ? io_in_4_bits_uop_bp_debug_if : io_in_5_valid ? io_in_5_bits_uop_bp_debug_if : io_in_6_valid ? io_in_6_bits_uop_bp_debug_if : io_in_7_bits_uop_bp_debug_if;
  assign io_out_bits_uop_bp_xcpt_if = io_in_0_valid ? io_in_0_bits_uop_bp_xcpt_if : io_in_1_valid ? io_in_1_bits_uop_bp_xcpt_if : io_in_2_valid ? io_in_2_bits_uop_bp_xcpt_if : io_in_3_valid ? io_in_3_bits_uop_bp_xcpt_if : io_in_4_valid ? io_in_4_bits_uop_bp_xcpt_if : io_in_5_valid ? io_in_5_bits_uop_bp_xcpt_if : io_in_6_valid ? io_in_6_bits_uop_bp_xcpt_if : io_in_7_bits_uop_bp_xcpt_if;
  assign io_out_bits_uop_debug_fsrc = io_in_0_valid ? io_in_0_bits_uop_debug_fsrc : io_in_1_valid ? io_in_1_bits_uop_debug_fsrc : io_in_2_valid ? io_in_2_bits_uop_debug_fsrc : io_in_3_valid ? io_in_3_bits_uop_debug_fsrc : io_in_4_valid ? io_in_4_bits_uop_debug_fsrc : io_in_5_valid ? io_in_5_bits_uop_debug_fsrc : io_in_6_valid ? io_in_6_bits_uop_debug_fsrc : io_in_7_bits_uop_debug_fsrc;
  assign io_out_bits_uop_debug_tsrc = io_in_0_valid ? io_in_0_bits_uop_debug_tsrc : io_in_1_valid ? io_in_1_bits_uop_debug_tsrc : io_in_2_valid ? io_in_2_bits_uop_debug_tsrc : io_in_3_valid ? io_in_3_bits_uop_debug_tsrc : io_in_4_valid ? io_in_4_bits_uop_debug_tsrc : io_in_5_valid ? io_in_5_bits_uop_debug_tsrc : io_in_6_valid ? io_in_6_bits_uop_debug_tsrc : io_in_7_bits_uop_debug_tsrc;
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_valid ? io_in_1_bits_addr : io_in_2_valid ? io_in_2_bits_addr : io_in_3_valid ? io_in_3_bits_addr : io_in_4_valid ? io_in_4_bits_addr : io_in_5_valid ? io_in_5_bits_addr : io_in_6_valid ? io_in_6_bits_addr : io_in_7_bits_addr;
  assign io_out_bits_is_hella = io_in_0_valid ? io_in_0_bits_is_hella : io_in_1_valid ? io_in_1_bits_is_hella : io_in_2_valid ? io_in_2_bits_is_hella : io_in_3_valid ? io_in_3_bits_is_hella : io_in_4_valid ? io_in_4_bits_is_hella : io_in_5_valid ? io_in_5_bits_is_hella : io_in_6_valid ? io_in_6_bits_is_hella : io_in_7_bits_is_hella;
  assign io_out_bits_way_en = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_valid ? io_in_1_bits_way_en : io_in_2_valid ? io_in_2_bits_way_en : io_in_3_valid ? io_in_3_bits_way_en : io_in_4_valid ? io_in_4_bits_way_en : io_in_5_valid ? io_in_5_bits_way_en : io_in_6_valid ? io_in_6_bits_way_en : io_in_7_bits_way_en;
  assign io_out_bits_sdq_id = io_in_0_valid ? io_in_0_bits_sdq_id : io_in_1_valid ? io_in_1_bits_sdq_id : io_in_2_valid ? io_in_2_bits_sdq_id : io_in_3_valid ? io_in_3_bits_sdq_id : io_in_4_valid ? io_in_4_bits_sdq_id : io_in_5_valid ? io_in_5_bits_sdq_id : io_in_6_valid ? io_in_6_bits_sdq_id : io_in_7_bits_sdq_id;
endmodule

