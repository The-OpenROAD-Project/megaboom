// Standard header to adapt well known macros for prints and assertions.

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module IssueUnitCollapsing_1(
  input         clock,
                reset,
  output        io_dis_uops_0_ready,
  input         io_dis_uops_0_valid,
  input  [6:0]  io_dis_uops_0_bits_uopc,
  input  [31:0] io_dis_uops_0_bits_inst,
                io_dis_uops_0_bits_debug_inst,
  input         io_dis_uops_0_bits_is_rvc,
  input  [39:0] io_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_dis_uops_0_bits_iq_type,
  input  [9:0]  io_dis_uops_0_bits_fu_code,
  input         io_dis_uops_0_bits_is_br,
                io_dis_uops_0_bits_is_jalr,
                io_dis_uops_0_bits_is_jal,
                io_dis_uops_0_bits_is_sfb,
  input  [19:0] io_dis_uops_0_bits_br_mask,
  input  [4:0]  io_dis_uops_0_bits_br_tag,
  input  [5:0]  io_dis_uops_0_bits_ftq_idx,
  input         io_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_dis_uops_0_bits_pc_lob,
  input         io_dis_uops_0_bits_taken,
  input  [19:0] io_dis_uops_0_bits_imm_packed,
  input  [11:0] io_dis_uops_0_bits_csr_addr,
  input  [6:0]  io_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_dis_uops_0_bits_ldq_idx,
                io_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_dis_uops_0_bits_pdst,
                io_dis_uops_0_bits_prs1,
                io_dis_uops_0_bits_prs2,
                io_dis_uops_0_bits_prs3,
  input         io_dis_uops_0_bits_prs1_busy,
                io_dis_uops_0_bits_prs2_busy,
  input  [6:0]  io_dis_uops_0_bits_stale_pdst,
  input         io_dis_uops_0_bits_exception,
  input  [63:0] io_dis_uops_0_bits_exc_cause,
  input         io_dis_uops_0_bits_bypassable,
  input  [4:0]  io_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_dis_uops_0_bits_mem_size,
  input         io_dis_uops_0_bits_mem_signed,
                io_dis_uops_0_bits_is_fence,
                io_dis_uops_0_bits_is_fencei,
                io_dis_uops_0_bits_is_amo,
                io_dis_uops_0_bits_uses_ldq,
                io_dis_uops_0_bits_uses_stq,
                io_dis_uops_0_bits_is_sys_pc2epc,
                io_dis_uops_0_bits_is_unique,
                io_dis_uops_0_bits_flush_on_commit,
                io_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_0_bits_ldst,
                io_dis_uops_0_bits_lrs1,
                io_dis_uops_0_bits_lrs2,
                io_dis_uops_0_bits_lrs3,
  input         io_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_dis_uops_0_bits_dst_rtype,
                io_dis_uops_0_bits_lrs1_rtype,
                io_dis_uops_0_bits_lrs2_rtype,
  input         io_dis_uops_0_bits_frs3_en,
                io_dis_uops_0_bits_fp_val,
                io_dis_uops_0_bits_fp_single,
                io_dis_uops_0_bits_xcpt_pf_if,
                io_dis_uops_0_bits_xcpt_ae_if,
                io_dis_uops_0_bits_xcpt_ma_if,
                io_dis_uops_0_bits_bp_debug_if,
                io_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_0_bits_debug_fsrc,
                io_dis_uops_0_bits_debug_tsrc,
  output        io_dis_uops_1_ready,
  input         io_dis_uops_1_valid,
  input  [6:0]  io_dis_uops_1_bits_uopc,
  input  [31:0] io_dis_uops_1_bits_inst,
                io_dis_uops_1_bits_debug_inst,
  input         io_dis_uops_1_bits_is_rvc,
  input  [39:0] io_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_dis_uops_1_bits_iq_type,
  input  [9:0]  io_dis_uops_1_bits_fu_code,
  input         io_dis_uops_1_bits_is_br,
                io_dis_uops_1_bits_is_jalr,
                io_dis_uops_1_bits_is_jal,
                io_dis_uops_1_bits_is_sfb,
  input  [19:0] io_dis_uops_1_bits_br_mask,
  input  [4:0]  io_dis_uops_1_bits_br_tag,
  input  [5:0]  io_dis_uops_1_bits_ftq_idx,
  input         io_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_dis_uops_1_bits_pc_lob,
  input         io_dis_uops_1_bits_taken,
  input  [19:0] io_dis_uops_1_bits_imm_packed,
  input  [11:0] io_dis_uops_1_bits_csr_addr,
  input  [6:0]  io_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_dis_uops_1_bits_ldq_idx,
                io_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_dis_uops_1_bits_pdst,
                io_dis_uops_1_bits_prs1,
                io_dis_uops_1_bits_prs2,
                io_dis_uops_1_bits_prs3,
  input         io_dis_uops_1_bits_prs1_busy,
                io_dis_uops_1_bits_prs2_busy,
  input  [6:0]  io_dis_uops_1_bits_stale_pdst,
  input         io_dis_uops_1_bits_exception,
  input  [63:0] io_dis_uops_1_bits_exc_cause,
  input         io_dis_uops_1_bits_bypassable,
  input  [4:0]  io_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_dis_uops_1_bits_mem_size,
  input         io_dis_uops_1_bits_mem_signed,
                io_dis_uops_1_bits_is_fence,
                io_dis_uops_1_bits_is_fencei,
                io_dis_uops_1_bits_is_amo,
                io_dis_uops_1_bits_uses_ldq,
                io_dis_uops_1_bits_uses_stq,
                io_dis_uops_1_bits_is_sys_pc2epc,
                io_dis_uops_1_bits_is_unique,
                io_dis_uops_1_bits_flush_on_commit,
                io_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_1_bits_ldst,
                io_dis_uops_1_bits_lrs1,
                io_dis_uops_1_bits_lrs2,
                io_dis_uops_1_bits_lrs3,
  input         io_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_dis_uops_1_bits_dst_rtype,
                io_dis_uops_1_bits_lrs1_rtype,
                io_dis_uops_1_bits_lrs2_rtype,
  input         io_dis_uops_1_bits_frs3_en,
                io_dis_uops_1_bits_fp_val,
                io_dis_uops_1_bits_fp_single,
                io_dis_uops_1_bits_xcpt_pf_if,
                io_dis_uops_1_bits_xcpt_ae_if,
                io_dis_uops_1_bits_xcpt_ma_if,
                io_dis_uops_1_bits_bp_debug_if,
                io_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_1_bits_debug_fsrc,
                io_dis_uops_1_bits_debug_tsrc,
  output        io_dis_uops_2_ready,
  input         io_dis_uops_2_valid,
  input  [6:0]  io_dis_uops_2_bits_uopc,
  input  [31:0] io_dis_uops_2_bits_inst,
                io_dis_uops_2_bits_debug_inst,
  input         io_dis_uops_2_bits_is_rvc,
  input  [39:0] io_dis_uops_2_bits_debug_pc,
  input  [2:0]  io_dis_uops_2_bits_iq_type,
  input  [9:0]  io_dis_uops_2_bits_fu_code,
  input         io_dis_uops_2_bits_is_br,
                io_dis_uops_2_bits_is_jalr,
                io_dis_uops_2_bits_is_jal,
                io_dis_uops_2_bits_is_sfb,
  input  [19:0] io_dis_uops_2_bits_br_mask,
  input  [4:0]  io_dis_uops_2_bits_br_tag,
  input  [5:0]  io_dis_uops_2_bits_ftq_idx,
  input         io_dis_uops_2_bits_edge_inst,
  input  [5:0]  io_dis_uops_2_bits_pc_lob,
  input         io_dis_uops_2_bits_taken,
  input  [19:0] io_dis_uops_2_bits_imm_packed,
  input  [11:0] io_dis_uops_2_bits_csr_addr,
  input  [6:0]  io_dis_uops_2_bits_rob_idx,
  input  [4:0]  io_dis_uops_2_bits_ldq_idx,
                io_dis_uops_2_bits_stq_idx,
  input  [1:0]  io_dis_uops_2_bits_rxq_idx,
  input  [6:0]  io_dis_uops_2_bits_pdst,
                io_dis_uops_2_bits_prs1,
                io_dis_uops_2_bits_prs2,
                io_dis_uops_2_bits_prs3,
  input         io_dis_uops_2_bits_prs1_busy,
                io_dis_uops_2_bits_prs2_busy,
  input  [6:0]  io_dis_uops_2_bits_stale_pdst,
  input         io_dis_uops_2_bits_exception,
  input  [63:0] io_dis_uops_2_bits_exc_cause,
  input         io_dis_uops_2_bits_bypassable,
  input  [4:0]  io_dis_uops_2_bits_mem_cmd,
  input  [1:0]  io_dis_uops_2_bits_mem_size,
  input         io_dis_uops_2_bits_mem_signed,
                io_dis_uops_2_bits_is_fence,
                io_dis_uops_2_bits_is_fencei,
                io_dis_uops_2_bits_is_amo,
                io_dis_uops_2_bits_uses_ldq,
                io_dis_uops_2_bits_uses_stq,
                io_dis_uops_2_bits_is_sys_pc2epc,
                io_dis_uops_2_bits_is_unique,
                io_dis_uops_2_bits_flush_on_commit,
                io_dis_uops_2_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_2_bits_ldst,
                io_dis_uops_2_bits_lrs1,
                io_dis_uops_2_bits_lrs2,
                io_dis_uops_2_bits_lrs3,
  input         io_dis_uops_2_bits_ldst_val,
  input  [1:0]  io_dis_uops_2_bits_dst_rtype,
                io_dis_uops_2_bits_lrs1_rtype,
                io_dis_uops_2_bits_lrs2_rtype,
  input         io_dis_uops_2_bits_frs3_en,
                io_dis_uops_2_bits_fp_val,
                io_dis_uops_2_bits_fp_single,
                io_dis_uops_2_bits_xcpt_pf_if,
                io_dis_uops_2_bits_xcpt_ae_if,
                io_dis_uops_2_bits_xcpt_ma_if,
                io_dis_uops_2_bits_bp_debug_if,
                io_dis_uops_2_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_2_bits_debug_fsrc,
                io_dis_uops_2_bits_debug_tsrc,
  output        io_dis_uops_3_ready,
  input         io_dis_uops_3_valid,
  input  [6:0]  io_dis_uops_3_bits_uopc,
  input  [31:0] io_dis_uops_3_bits_inst,
                io_dis_uops_3_bits_debug_inst,
  input         io_dis_uops_3_bits_is_rvc,
  input  [39:0] io_dis_uops_3_bits_debug_pc,
  input  [2:0]  io_dis_uops_3_bits_iq_type,
  input  [9:0]  io_dis_uops_3_bits_fu_code,
  input         io_dis_uops_3_bits_is_br,
                io_dis_uops_3_bits_is_jalr,
                io_dis_uops_3_bits_is_jal,
                io_dis_uops_3_bits_is_sfb,
  input  [19:0] io_dis_uops_3_bits_br_mask,
  input  [4:0]  io_dis_uops_3_bits_br_tag,
  input  [5:0]  io_dis_uops_3_bits_ftq_idx,
  input         io_dis_uops_3_bits_edge_inst,
  input  [5:0]  io_dis_uops_3_bits_pc_lob,
  input         io_dis_uops_3_bits_taken,
  input  [19:0] io_dis_uops_3_bits_imm_packed,
  input  [11:0] io_dis_uops_3_bits_csr_addr,
  input  [6:0]  io_dis_uops_3_bits_rob_idx,
  input  [4:0]  io_dis_uops_3_bits_ldq_idx,
                io_dis_uops_3_bits_stq_idx,
  input  [1:0]  io_dis_uops_3_bits_rxq_idx,
  input  [6:0]  io_dis_uops_3_bits_pdst,
                io_dis_uops_3_bits_prs1,
                io_dis_uops_3_bits_prs2,
                io_dis_uops_3_bits_prs3,
  input         io_dis_uops_3_bits_prs1_busy,
                io_dis_uops_3_bits_prs2_busy,
  input  [6:0]  io_dis_uops_3_bits_stale_pdst,
  input         io_dis_uops_3_bits_exception,
  input  [63:0] io_dis_uops_3_bits_exc_cause,
  input         io_dis_uops_3_bits_bypassable,
  input  [4:0]  io_dis_uops_3_bits_mem_cmd,
  input  [1:0]  io_dis_uops_3_bits_mem_size,
  input         io_dis_uops_3_bits_mem_signed,
                io_dis_uops_3_bits_is_fence,
                io_dis_uops_3_bits_is_fencei,
                io_dis_uops_3_bits_is_amo,
                io_dis_uops_3_bits_uses_ldq,
                io_dis_uops_3_bits_uses_stq,
                io_dis_uops_3_bits_is_sys_pc2epc,
                io_dis_uops_3_bits_is_unique,
                io_dis_uops_3_bits_flush_on_commit,
                io_dis_uops_3_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_3_bits_ldst,
                io_dis_uops_3_bits_lrs1,
                io_dis_uops_3_bits_lrs2,
                io_dis_uops_3_bits_lrs3,
  input         io_dis_uops_3_bits_ldst_val,
  input  [1:0]  io_dis_uops_3_bits_dst_rtype,
                io_dis_uops_3_bits_lrs1_rtype,
                io_dis_uops_3_bits_lrs2_rtype,
  input         io_dis_uops_3_bits_frs3_en,
                io_dis_uops_3_bits_fp_val,
                io_dis_uops_3_bits_fp_single,
                io_dis_uops_3_bits_xcpt_pf_if,
                io_dis_uops_3_bits_xcpt_ae_if,
                io_dis_uops_3_bits_xcpt_ma_if,
                io_dis_uops_3_bits_bp_debug_if,
                io_dis_uops_3_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_3_bits_debug_fsrc,
                io_dis_uops_3_bits_debug_tsrc,
  output        io_iss_valids_0,
                io_iss_valids_1,
  output [6:0]  io_iss_uops_0_uopc,
  output [31:0] io_iss_uops_0_inst,
                io_iss_uops_0_debug_inst,
  output        io_iss_uops_0_is_rvc,
  output [39:0] io_iss_uops_0_debug_pc,
  output [2:0]  io_iss_uops_0_iq_type,
  output [9:0]  io_iss_uops_0_fu_code,
  output [1:0]  io_iss_uops_0_iw_state,
  output        io_iss_uops_0_iw_p1_poisoned,
                io_iss_uops_0_iw_p2_poisoned,
                io_iss_uops_0_is_br,
                io_iss_uops_0_is_jalr,
                io_iss_uops_0_is_jal,
                io_iss_uops_0_is_sfb,
  output [19:0] io_iss_uops_0_br_mask,
  output [4:0]  io_iss_uops_0_br_tag,
  output [5:0]  io_iss_uops_0_ftq_idx,
  output        io_iss_uops_0_edge_inst,
  output [5:0]  io_iss_uops_0_pc_lob,
  output        io_iss_uops_0_taken,
  output [19:0] io_iss_uops_0_imm_packed,
  output [11:0] io_iss_uops_0_csr_addr,
  output [6:0]  io_iss_uops_0_rob_idx,
  output [4:0]  io_iss_uops_0_ldq_idx,
                io_iss_uops_0_stq_idx,
  output [1:0]  io_iss_uops_0_rxq_idx,
  output [6:0]  io_iss_uops_0_pdst,
                io_iss_uops_0_prs1,
                io_iss_uops_0_prs2,
                io_iss_uops_0_prs3,
  output [5:0]  io_iss_uops_0_ppred,
  output        io_iss_uops_0_prs1_busy,
                io_iss_uops_0_prs2_busy,
                io_iss_uops_0_prs3_busy,
                io_iss_uops_0_ppred_busy,
  output [6:0]  io_iss_uops_0_stale_pdst,
  output        io_iss_uops_0_exception,
  output [63:0] io_iss_uops_0_exc_cause,
  output        io_iss_uops_0_bypassable,
  output [4:0]  io_iss_uops_0_mem_cmd,
  output [1:0]  io_iss_uops_0_mem_size,
  output        io_iss_uops_0_mem_signed,
                io_iss_uops_0_is_fence,
                io_iss_uops_0_is_fencei,
                io_iss_uops_0_is_amo,
                io_iss_uops_0_uses_ldq,
                io_iss_uops_0_uses_stq,
                io_iss_uops_0_is_sys_pc2epc,
                io_iss_uops_0_is_unique,
                io_iss_uops_0_flush_on_commit,
                io_iss_uops_0_ldst_is_rs1,
  output [5:0]  io_iss_uops_0_ldst,
                io_iss_uops_0_lrs1,
                io_iss_uops_0_lrs2,
                io_iss_uops_0_lrs3,
  output        io_iss_uops_0_ldst_val,
  output [1:0]  io_iss_uops_0_dst_rtype,
                io_iss_uops_0_lrs1_rtype,
                io_iss_uops_0_lrs2_rtype,
  output        io_iss_uops_0_frs3_en,
                io_iss_uops_0_fp_val,
                io_iss_uops_0_fp_single,
                io_iss_uops_0_xcpt_pf_if,
                io_iss_uops_0_xcpt_ae_if,
                io_iss_uops_0_xcpt_ma_if,
                io_iss_uops_0_bp_debug_if,
                io_iss_uops_0_bp_xcpt_if,
  output [1:0]  io_iss_uops_0_debug_fsrc,
                io_iss_uops_0_debug_tsrc,
  output [6:0]  io_iss_uops_1_uopc,
  output [31:0] io_iss_uops_1_inst,
                io_iss_uops_1_debug_inst,
  output        io_iss_uops_1_is_rvc,
  output [39:0] io_iss_uops_1_debug_pc,
  output [2:0]  io_iss_uops_1_iq_type,
  output [9:0]  io_iss_uops_1_fu_code,
  output [1:0]  io_iss_uops_1_iw_state,
  output        io_iss_uops_1_iw_p1_poisoned,
                io_iss_uops_1_iw_p2_poisoned,
                io_iss_uops_1_is_br,
                io_iss_uops_1_is_jalr,
                io_iss_uops_1_is_jal,
                io_iss_uops_1_is_sfb,
  output [19:0] io_iss_uops_1_br_mask,
  output [4:0]  io_iss_uops_1_br_tag,
  output [5:0]  io_iss_uops_1_ftq_idx,
  output        io_iss_uops_1_edge_inst,
  output [5:0]  io_iss_uops_1_pc_lob,
  output        io_iss_uops_1_taken,
  output [19:0] io_iss_uops_1_imm_packed,
  output [11:0] io_iss_uops_1_csr_addr,
  output [6:0]  io_iss_uops_1_rob_idx,
  output [4:0]  io_iss_uops_1_ldq_idx,
                io_iss_uops_1_stq_idx,
  output [1:0]  io_iss_uops_1_rxq_idx,
  output [6:0]  io_iss_uops_1_pdst,
                io_iss_uops_1_prs1,
                io_iss_uops_1_prs2,
                io_iss_uops_1_prs3,
  output [5:0]  io_iss_uops_1_ppred,
  output        io_iss_uops_1_prs1_busy,
                io_iss_uops_1_prs2_busy,
                io_iss_uops_1_prs3_busy,
                io_iss_uops_1_ppred_busy,
  output [6:0]  io_iss_uops_1_stale_pdst,
  output        io_iss_uops_1_exception,
  output [63:0] io_iss_uops_1_exc_cause,
  output        io_iss_uops_1_bypassable,
  output [4:0]  io_iss_uops_1_mem_cmd,
  output [1:0]  io_iss_uops_1_mem_size,
  output        io_iss_uops_1_mem_signed,
                io_iss_uops_1_is_fence,
                io_iss_uops_1_is_fencei,
                io_iss_uops_1_is_amo,
                io_iss_uops_1_uses_ldq,
                io_iss_uops_1_uses_stq,
                io_iss_uops_1_is_sys_pc2epc,
                io_iss_uops_1_is_unique,
                io_iss_uops_1_flush_on_commit,
                io_iss_uops_1_ldst_is_rs1,
  output [5:0]  io_iss_uops_1_ldst,
                io_iss_uops_1_lrs1,
                io_iss_uops_1_lrs2,
                io_iss_uops_1_lrs3,
  output        io_iss_uops_1_ldst_val,
  output [1:0]  io_iss_uops_1_dst_rtype,
                io_iss_uops_1_lrs1_rtype,
                io_iss_uops_1_lrs2_rtype,
  output        io_iss_uops_1_frs3_en,
                io_iss_uops_1_fp_val,
                io_iss_uops_1_fp_single,
                io_iss_uops_1_xcpt_pf_if,
                io_iss_uops_1_xcpt_ae_if,
                io_iss_uops_1_xcpt_ma_if,
                io_iss_uops_1_bp_debug_if,
                io_iss_uops_1_bp_xcpt_if,
  output [1:0]  io_iss_uops_1_debug_fsrc,
                io_iss_uops_1_debug_tsrc,
  input         io_wakeup_ports_0_valid,
  input  [6:0]  io_wakeup_ports_0_bits_pdst,
  input         io_wakeup_ports_1_valid,
  input  [6:0]  io_wakeup_ports_1_bits_pdst,
  input         io_wakeup_ports_2_valid,
  input  [6:0]  io_wakeup_ports_2_bits_pdst,
  input         io_wakeup_ports_3_valid,
  input  [6:0]  io_wakeup_ports_3_bits_pdst,
  input         io_wakeup_ports_4_valid,
  input  [6:0]  io_wakeup_ports_4_bits_pdst,
  input         io_wakeup_ports_5_valid,
  input  [6:0]  io_wakeup_ports_5_bits_pdst,
  input         io_wakeup_ports_6_valid,
  input  [6:0]  io_wakeup_ports_6_bits_pdst,
  input         io_wakeup_ports_7_valid,
  input  [6:0]  io_wakeup_ports_7_bits_pdst,
  input         io_wakeup_ports_8_valid,
  input  [6:0]  io_wakeup_ports_8_bits_pdst,
  input         io_wakeup_ports_9_valid,
  input  [6:0]  io_wakeup_ports_9_bits_pdst,
  input         io_spec_ld_wakeup_0_valid,
  input  [6:0]  io_spec_ld_wakeup_0_bits,
  input         io_spec_ld_wakeup_1_valid,
  input  [6:0]  io_spec_ld_wakeup_1_bits,
  input  [9:0]  io_fu_types_0,
                io_fu_types_1,
  input  [19:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input         io_flush_pipeline,
                io_ld_miss
);

  wire        issue_slots_23_grant;
  wire        issue_slots_22_grant;
  wire        issue_slots_21_grant;
  wire        issue_slots_20_grant;
  wire        issue_slots_19_grant;
  wire        issue_slots_18_grant;
  wire        issue_slots_17_grant;
  wire        issue_slots_16_grant;
  wire        issue_slots_15_grant;
  wire        issue_slots_14_grant;
  wire        issue_slots_13_grant;
  wire        issue_slots_12_grant;
  wire        issue_slots_11_grant;
  wire        issue_slots_10_grant;
  wire        issue_slots_9_grant;
  wire        issue_slots_8_grant;
  wire        issue_slots_7_grant;
  wire        issue_slots_6_grant;
  wire        issue_slots_5_grant;
  wire        issue_slots_4_grant;
  wire        issue_slots_3_grant;
  wire        issue_slots_2_grant;
  wire        issue_slots_1_grant;
  wire        issue_slots_0_grant;
  wire [3:0]  next_22;
  wire [3:0]  next_21;
  wire [3:0]  next_20;
  wire [3:0]  next_19;
  wire [3:0]  next_18;
  wire [3:0]  next_17;
  wire [3:0]  next_16;
  wire [3:0]  next_15;
  wire [3:0]  next_14;
  wire [3:0]  next_13;
  wire [3:0]  next_12;
  wire [3:0]  next_11;
  wire [3:0]  next_10;
  wire [3:0]  next_9;
  wire [3:0]  next_8;
  wire [3:0]  next_7;
  wire [3:0]  next_6;
  wire [3:0]  next_5;
  wire [3:0]  next_4;
  wire [3:0]  next_3;
  wire [3:0]  next_2;
  wire [1:0]  _next_1_1to0;
  wire        _slots_23_io_valid;
  wire        _slots_23_io_will_be_valid;
  wire        _slots_23_io_request;
  wire [6:0]  _slots_23_io_out_uop_uopc;
  wire [31:0] _slots_23_io_out_uop_inst;
  wire [31:0] _slots_23_io_out_uop_debug_inst;
  wire        _slots_23_io_out_uop_is_rvc;
  wire [39:0] _slots_23_io_out_uop_debug_pc;
  wire [2:0]  _slots_23_io_out_uop_iq_type;
  wire [9:0]  _slots_23_io_out_uop_fu_code;
  wire [1:0]  _slots_23_io_out_uop_iw_state;
  wire        _slots_23_io_out_uop_iw_p1_poisoned;
  wire        _slots_23_io_out_uop_iw_p2_poisoned;
  wire        _slots_23_io_out_uop_is_br;
  wire        _slots_23_io_out_uop_is_jalr;
  wire        _slots_23_io_out_uop_is_jal;
  wire        _slots_23_io_out_uop_is_sfb;
  wire [19:0] _slots_23_io_out_uop_br_mask;
  wire [4:0]  _slots_23_io_out_uop_br_tag;
  wire [5:0]  _slots_23_io_out_uop_ftq_idx;
  wire        _slots_23_io_out_uop_edge_inst;
  wire [5:0]  _slots_23_io_out_uop_pc_lob;
  wire        _slots_23_io_out_uop_taken;
  wire [19:0] _slots_23_io_out_uop_imm_packed;
  wire [11:0] _slots_23_io_out_uop_csr_addr;
  wire [6:0]  _slots_23_io_out_uop_rob_idx;
  wire [4:0]  _slots_23_io_out_uop_ldq_idx;
  wire [4:0]  _slots_23_io_out_uop_stq_idx;
  wire [1:0]  _slots_23_io_out_uop_rxq_idx;
  wire [6:0]  _slots_23_io_out_uop_pdst;
  wire [6:0]  _slots_23_io_out_uop_prs1;
  wire [6:0]  _slots_23_io_out_uop_prs2;
  wire [6:0]  _slots_23_io_out_uop_prs3;
  wire [5:0]  _slots_23_io_out_uop_ppred;
  wire        _slots_23_io_out_uop_prs1_busy;
  wire        _slots_23_io_out_uop_prs2_busy;
  wire        _slots_23_io_out_uop_prs3_busy;
  wire        _slots_23_io_out_uop_ppred_busy;
  wire [6:0]  _slots_23_io_out_uop_stale_pdst;
  wire        _slots_23_io_out_uop_exception;
  wire [63:0] _slots_23_io_out_uop_exc_cause;
  wire        _slots_23_io_out_uop_bypassable;
  wire [4:0]  _slots_23_io_out_uop_mem_cmd;
  wire [1:0]  _slots_23_io_out_uop_mem_size;
  wire        _slots_23_io_out_uop_mem_signed;
  wire        _slots_23_io_out_uop_is_fence;
  wire        _slots_23_io_out_uop_is_fencei;
  wire        _slots_23_io_out_uop_is_amo;
  wire        _slots_23_io_out_uop_uses_ldq;
  wire        _slots_23_io_out_uop_uses_stq;
  wire        _slots_23_io_out_uop_is_sys_pc2epc;
  wire        _slots_23_io_out_uop_is_unique;
  wire        _slots_23_io_out_uop_flush_on_commit;
  wire        _slots_23_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_23_io_out_uop_ldst;
  wire [5:0]  _slots_23_io_out_uop_lrs1;
  wire [5:0]  _slots_23_io_out_uop_lrs2;
  wire [5:0]  _slots_23_io_out_uop_lrs3;
  wire        _slots_23_io_out_uop_ldst_val;
  wire [1:0]  _slots_23_io_out_uop_dst_rtype;
  wire [1:0]  _slots_23_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_23_io_out_uop_lrs2_rtype;
  wire        _slots_23_io_out_uop_frs3_en;
  wire        _slots_23_io_out_uop_fp_val;
  wire        _slots_23_io_out_uop_fp_single;
  wire        _slots_23_io_out_uop_xcpt_pf_if;
  wire        _slots_23_io_out_uop_xcpt_ae_if;
  wire        _slots_23_io_out_uop_xcpt_ma_if;
  wire        _slots_23_io_out_uop_bp_debug_if;
  wire        _slots_23_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_23_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_23_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_23_io_uop_uopc;
  wire [31:0] _slots_23_io_uop_inst;
  wire [31:0] _slots_23_io_uop_debug_inst;
  wire        _slots_23_io_uop_is_rvc;
  wire [39:0] _slots_23_io_uop_debug_pc;
  wire [2:0]  _slots_23_io_uop_iq_type;
  wire [9:0]  _slots_23_io_uop_fu_code;
  wire [1:0]  _slots_23_io_uop_iw_state;
  wire        _slots_23_io_uop_iw_p1_poisoned;
  wire        _slots_23_io_uop_iw_p2_poisoned;
  wire        _slots_23_io_uop_is_br;
  wire        _slots_23_io_uop_is_jalr;
  wire        _slots_23_io_uop_is_jal;
  wire        _slots_23_io_uop_is_sfb;
  wire [19:0] _slots_23_io_uop_br_mask;
  wire [4:0]  _slots_23_io_uop_br_tag;
  wire [5:0]  _slots_23_io_uop_ftq_idx;
  wire        _slots_23_io_uop_edge_inst;
  wire [5:0]  _slots_23_io_uop_pc_lob;
  wire        _slots_23_io_uop_taken;
  wire [19:0] _slots_23_io_uop_imm_packed;
  wire [11:0] _slots_23_io_uop_csr_addr;
  wire [6:0]  _slots_23_io_uop_rob_idx;
  wire [4:0]  _slots_23_io_uop_ldq_idx;
  wire [4:0]  _slots_23_io_uop_stq_idx;
  wire [1:0]  _slots_23_io_uop_rxq_idx;
  wire [6:0]  _slots_23_io_uop_pdst;
  wire [6:0]  _slots_23_io_uop_prs1;
  wire [6:0]  _slots_23_io_uop_prs2;
  wire [6:0]  _slots_23_io_uop_prs3;
  wire [5:0]  _slots_23_io_uop_ppred;
  wire        _slots_23_io_uop_prs1_busy;
  wire        _slots_23_io_uop_prs2_busy;
  wire        _slots_23_io_uop_prs3_busy;
  wire        _slots_23_io_uop_ppred_busy;
  wire [6:0]  _slots_23_io_uop_stale_pdst;
  wire        _slots_23_io_uop_exception;
  wire [63:0] _slots_23_io_uop_exc_cause;
  wire        _slots_23_io_uop_bypassable;
  wire [4:0]  _slots_23_io_uop_mem_cmd;
  wire [1:0]  _slots_23_io_uop_mem_size;
  wire        _slots_23_io_uop_mem_signed;
  wire        _slots_23_io_uop_is_fence;
  wire        _slots_23_io_uop_is_fencei;
  wire        _slots_23_io_uop_is_amo;
  wire        _slots_23_io_uop_uses_ldq;
  wire        _slots_23_io_uop_uses_stq;
  wire        _slots_23_io_uop_is_sys_pc2epc;
  wire        _slots_23_io_uop_is_unique;
  wire        _slots_23_io_uop_flush_on_commit;
  wire        _slots_23_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_23_io_uop_ldst;
  wire [5:0]  _slots_23_io_uop_lrs1;
  wire [5:0]  _slots_23_io_uop_lrs2;
  wire [5:0]  _slots_23_io_uop_lrs3;
  wire        _slots_23_io_uop_ldst_val;
  wire [1:0]  _slots_23_io_uop_dst_rtype;
  wire [1:0]  _slots_23_io_uop_lrs1_rtype;
  wire [1:0]  _slots_23_io_uop_lrs2_rtype;
  wire        _slots_23_io_uop_frs3_en;
  wire        _slots_23_io_uop_fp_val;
  wire        _slots_23_io_uop_fp_single;
  wire        _slots_23_io_uop_xcpt_pf_if;
  wire        _slots_23_io_uop_xcpt_ae_if;
  wire        _slots_23_io_uop_xcpt_ma_if;
  wire        _slots_23_io_uop_bp_debug_if;
  wire        _slots_23_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_23_io_uop_debug_fsrc;
  wire [1:0]  _slots_23_io_uop_debug_tsrc;
  wire        _slots_22_io_valid;
  wire        _slots_22_io_will_be_valid;
  wire        _slots_22_io_request;
  wire [6:0]  _slots_22_io_out_uop_uopc;
  wire [31:0] _slots_22_io_out_uop_inst;
  wire [31:0] _slots_22_io_out_uop_debug_inst;
  wire        _slots_22_io_out_uop_is_rvc;
  wire [39:0] _slots_22_io_out_uop_debug_pc;
  wire [2:0]  _slots_22_io_out_uop_iq_type;
  wire [9:0]  _slots_22_io_out_uop_fu_code;
  wire [1:0]  _slots_22_io_out_uop_iw_state;
  wire        _slots_22_io_out_uop_iw_p1_poisoned;
  wire        _slots_22_io_out_uop_iw_p2_poisoned;
  wire        _slots_22_io_out_uop_is_br;
  wire        _slots_22_io_out_uop_is_jalr;
  wire        _slots_22_io_out_uop_is_jal;
  wire        _slots_22_io_out_uop_is_sfb;
  wire [19:0] _slots_22_io_out_uop_br_mask;
  wire [4:0]  _slots_22_io_out_uop_br_tag;
  wire [5:0]  _slots_22_io_out_uop_ftq_idx;
  wire        _slots_22_io_out_uop_edge_inst;
  wire [5:0]  _slots_22_io_out_uop_pc_lob;
  wire        _slots_22_io_out_uop_taken;
  wire [19:0] _slots_22_io_out_uop_imm_packed;
  wire [11:0] _slots_22_io_out_uop_csr_addr;
  wire [6:0]  _slots_22_io_out_uop_rob_idx;
  wire [4:0]  _slots_22_io_out_uop_ldq_idx;
  wire [4:0]  _slots_22_io_out_uop_stq_idx;
  wire [1:0]  _slots_22_io_out_uop_rxq_idx;
  wire [6:0]  _slots_22_io_out_uop_pdst;
  wire [6:0]  _slots_22_io_out_uop_prs1;
  wire [6:0]  _slots_22_io_out_uop_prs2;
  wire [6:0]  _slots_22_io_out_uop_prs3;
  wire [5:0]  _slots_22_io_out_uop_ppred;
  wire        _slots_22_io_out_uop_prs1_busy;
  wire        _slots_22_io_out_uop_prs2_busy;
  wire        _slots_22_io_out_uop_prs3_busy;
  wire        _slots_22_io_out_uop_ppred_busy;
  wire [6:0]  _slots_22_io_out_uop_stale_pdst;
  wire        _slots_22_io_out_uop_exception;
  wire [63:0] _slots_22_io_out_uop_exc_cause;
  wire        _slots_22_io_out_uop_bypassable;
  wire [4:0]  _slots_22_io_out_uop_mem_cmd;
  wire [1:0]  _slots_22_io_out_uop_mem_size;
  wire        _slots_22_io_out_uop_mem_signed;
  wire        _slots_22_io_out_uop_is_fence;
  wire        _slots_22_io_out_uop_is_fencei;
  wire        _slots_22_io_out_uop_is_amo;
  wire        _slots_22_io_out_uop_uses_ldq;
  wire        _slots_22_io_out_uop_uses_stq;
  wire        _slots_22_io_out_uop_is_sys_pc2epc;
  wire        _slots_22_io_out_uop_is_unique;
  wire        _slots_22_io_out_uop_flush_on_commit;
  wire        _slots_22_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_22_io_out_uop_ldst;
  wire [5:0]  _slots_22_io_out_uop_lrs1;
  wire [5:0]  _slots_22_io_out_uop_lrs2;
  wire [5:0]  _slots_22_io_out_uop_lrs3;
  wire        _slots_22_io_out_uop_ldst_val;
  wire [1:0]  _slots_22_io_out_uop_dst_rtype;
  wire [1:0]  _slots_22_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_22_io_out_uop_lrs2_rtype;
  wire        _slots_22_io_out_uop_frs3_en;
  wire        _slots_22_io_out_uop_fp_val;
  wire        _slots_22_io_out_uop_fp_single;
  wire        _slots_22_io_out_uop_xcpt_pf_if;
  wire        _slots_22_io_out_uop_xcpt_ae_if;
  wire        _slots_22_io_out_uop_xcpt_ma_if;
  wire        _slots_22_io_out_uop_bp_debug_if;
  wire        _slots_22_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_22_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_22_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_22_io_uop_uopc;
  wire [31:0] _slots_22_io_uop_inst;
  wire [31:0] _slots_22_io_uop_debug_inst;
  wire        _slots_22_io_uop_is_rvc;
  wire [39:0] _slots_22_io_uop_debug_pc;
  wire [2:0]  _slots_22_io_uop_iq_type;
  wire [9:0]  _slots_22_io_uop_fu_code;
  wire [1:0]  _slots_22_io_uop_iw_state;
  wire        _slots_22_io_uop_iw_p1_poisoned;
  wire        _slots_22_io_uop_iw_p2_poisoned;
  wire        _slots_22_io_uop_is_br;
  wire        _slots_22_io_uop_is_jalr;
  wire        _slots_22_io_uop_is_jal;
  wire        _slots_22_io_uop_is_sfb;
  wire [19:0] _slots_22_io_uop_br_mask;
  wire [4:0]  _slots_22_io_uop_br_tag;
  wire [5:0]  _slots_22_io_uop_ftq_idx;
  wire        _slots_22_io_uop_edge_inst;
  wire [5:0]  _slots_22_io_uop_pc_lob;
  wire        _slots_22_io_uop_taken;
  wire [19:0] _slots_22_io_uop_imm_packed;
  wire [11:0] _slots_22_io_uop_csr_addr;
  wire [6:0]  _slots_22_io_uop_rob_idx;
  wire [4:0]  _slots_22_io_uop_ldq_idx;
  wire [4:0]  _slots_22_io_uop_stq_idx;
  wire [1:0]  _slots_22_io_uop_rxq_idx;
  wire [6:0]  _slots_22_io_uop_pdst;
  wire [6:0]  _slots_22_io_uop_prs1;
  wire [6:0]  _slots_22_io_uop_prs2;
  wire [6:0]  _slots_22_io_uop_prs3;
  wire [5:0]  _slots_22_io_uop_ppred;
  wire        _slots_22_io_uop_prs1_busy;
  wire        _slots_22_io_uop_prs2_busy;
  wire        _slots_22_io_uop_prs3_busy;
  wire        _slots_22_io_uop_ppred_busy;
  wire [6:0]  _slots_22_io_uop_stale_pdst;
  wire        _slots_22_io_uop_exception;
  wire [63:0] _slots_22_io_uop_exc_cause;
  wire        _slots_22_io_uop_bypassable;
  wire [4:0]  _slots_22_io_uop_mem_cmd;
  wire [1:0]  _slots_22_io_uop_mem_size;
  wire        _slots_22_io_uop_mem_signed;
  wire        _slots_22_io_uop_is_fence;
  wire        _slots_22_io_uop_is_fencei;
  wire        _slots_22_io_uop_is_amo;
  wire        _slots_22_io_uop_uses_ldq;
  wire        _slots_22_io_uop_uses_stq;
  wire        _slots_22_io_uop_is_sys_pc2epc;
  wire        _slots_22_io_uop_is_unique;
  wire        _slots_22_io_uop_flush_on_commit;
  wire        _slots_22_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_22_io_uop_ldst;
  wire [5:0]  _slots_22_io_uop_lrs1;
  wire [5:0]  _slots_22_io_uop_lrs2;
  wire [5:0]  _slots_22_io_uop_lrs3;
  wire        _slots_22_io_uop_ldst_val;
  wire [1:0]  _slots_22_io_uop_dst_rtype;
  wire [1:0]  _slots_22_io_uop_lrs1_rtype;
  wire [1:0]  _slots_22_io_uop_lrs2_rtype;
  wire        _slots_22_io_uop_frs3_en;
  wire        _slots_22_io_uop_fp_val;
  wire        _slots_22_io_uop_fp_single;
  wire        _slots_22_io_uop_xcpt_pf_if;
  wire        _slots_22_io_uop_xcpt_ae_if;
  wire        _slots_22_io_uop_xcpt_ma_if;
  wire        _slots_22_io_uop_bp_debug_if;
  wire        _slots_22_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_22_io_uop_debug_fsrc;
  wire [1:0]  _slots_22_io_uop_debug_tsrc;
  wire        _slots_21_io_valid;
  wire        _slots_21_io_will_be_valid;
  wire        _slots_21_io_request;
  wire [6:0]  _slots_21_io_out_uop_uopc;
  wire [31:0] _slots_21_io_out_uop_inst;
  wire [31:0] _slots_21_io_out_uop_debug_inst;
  wire        _slots_21_io_out_uop_is_rvc;
  wire [39:0] _slots_21_io_out_uop_debug_pc;
  wire [2:0]  _slots_21_io_out_uop_iq_type;
  wire [9:0]  _slots_21_io_out_uop_fu_code;
  wire [1:0]  _slots_21_io_out_uop_iw_state;
  wire        _slots_21_io_out_uop_iw_p1_poisoned;
  wire        _slots_21_io_out_uop_iw_p2_poisoned;
  wire        _slots_21_io_out_uop_is_br;
  wire        _slots_21_io_out_uop_is_jalr;
  wire        _slots_21_io_out_uop_is_jal;
  wire        _slots_21_io_out_uop_is_sfb;
  wire [19:0] _slots_21_io_out_uop_br_mask;
  wire [4:0]  _slots_21_io_out_uop_br_tag;
  wire [5:0]  _slots_21_io_out_uop_ftq_idx;
  wire        _slots_21_io_out_uop_edge_inst;
  wire [5:0]  _slots_21_io_out_uop_pc_lob;
  wire        _slots_21_io_out_uop_taken;
  wire [19:0] _slots_21_io_out_uop_imm_packed;
  wire [11:0] _slots_21_io_out_uop_csr_addr;
  wire [6:0]  _slots_21_io_out_uop_rob_idx;
  wire [4:0]  _slots_21_io_out_uop_ldq_idx;
  wire [4:0]  _slots_21_io_out_uop_stq_idx;
  wire [1:0]  _slots_21_io_out_uop_rxq_idx;
  wire [6:0]  _slots_21_io_out_uop_pdst;
  wire [6:0]  _slots_21_io_out_uop_prs1;
  wire [6:0]  _slots_21_io_out_uop_prs2;
  wire [6:0]  _slots_21_io_out_uop_prs3;
  wire [5:0]  _slots_21_io_out_uop_ppred;
  wire        _slots_21_io_out_uop_prs1_busy;
  wire        _slots_21_io_out_uop_prs2_busy;
  wire        _slots_21_io_out_uop_prs3_busy;
  wire        _slots_21_io_out_uop_ppred_busy;
  wire [6:0]  _slots_21_io_out_uop_stale_pdst;
  wire        _slots_21_io_out_uop_exception;
  wire [63:0] _slots_21_io_out_uop_exc_cause;
  wire        _slots_21_io_out_uop_bypassable;
  wire [4:0]  _slots_21_io_out_uop_mem_cmd;
  wire [1:0]  _slots_21_io_out_uop_mem_size;
  wire        _slots_21_io_out_uop_mem_signed;
  wire        _slots_21_io_out_uop_is_fence;
  wire        _slots_21_io_out_uop_is_fencei;
  wire        _slots_21_io_out_uop_is_amo;
  wire        _slots_21_io_out_uop_uses_ldq;
  wire        _slots_21_io_out_uop_uses_stq;
  wire        _slots_21_io_out_uop_is_sys_pc2epc;
  wire        _slots_21_io_out_uop_is_unique;
  wire        _slots_21_io_out_uop_flush_on_commit;
  wire        _slots_21_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_21_io_out_uop_ldst;
  wire [5:0]  _slots_21_io_out_uop_lrs1;
  wire [5:0]  _slots_21_io_out_uop_lrs2;
  wire [5:0]  _slots_21_io_out_uop_lrs3;
  wire        _slots_21_io_out_uop_ldst_val;
  wire [1:0]  _slots_21_io_out_uop_dst_rtype;
  wire [1:0]  _slots_21_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_21_io_out_uop_lrs2_rtype;
  wire        _slots_21_io_out_uop_frs3_en;
  wire        _slots_21_io_out_uop_fp_val;
  wire        _slots_21_io_out_uop_fp_single;
  wire        _slots_21_io_out_uop_xcpt_pf_if;
  wire        _slots_21_io_out_uop_xcpt_ae_if;
  wire        _slots_21_io_out_uop_xcpt_ma_if;
  wire        _slots_21_io_out_uop_bp_debug_if;
  wire        _slots_21_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_21_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_21_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_21_io_uop_uopc;
  wire [31:0] _slots_21_io_uop_inst;
  wire [31:0] _slots_21_io_uop_debug_inst;
  wire        _slots_21_io_uop_is_rvc;
  wire [39:0] _slots_21_io_uop_debug_pc;
  wire [2:0]  _slots_21_io_uop_iq_type;
  wire [9:0]  _slots_21_io_uop_fu_code;
  wire [1:0]  _slots_21_io_uop_iw_state;
  wire        _slots_21_io_uop_iw_p1_poisoned;
  wire        _slots_21_io_uop_iw_p2_poisoned;
  wire        _slots_21_io_uop_is_br;
  wire        _slots_21_io_uop_is_jalr;
  wire        _slots_21_io_uop_is_jal;
  wire        _slots_21_io_uop_is_sfb;
  wire [19:0] _slots_21_io_uop_br_mask;
  wire [4:0]  _slots_21_io_uop_br_tag;
  wire [5:0]  _slots_21_io_uop_ftq_idx;
  wire        _slots_21_io_uop_edge_inst;
  wire [5:0]  _slots_21_io_uop_pc_lob;
  wire        _slots_21_io_uop_taken;
  wire [19:0] _slots_21_io_uop_imm_packed;
  wire [11:0] _slots_21_io_uop_csr_addr;
  wire [6:0]  _slots_21_io_uop_rob_idx;
  wire [4:0]  _slots_21_io_uop_ldq_idx;
  wire [4:0]  _slots_21_io_uop_stq_idx;
  wire [1:0]  _slots_21_io_uop_rxq_idx;
  wire [6:0]  _slots_21_io_uop_pdst;
  wire [6:0]  _slots_21_io_uop_prs1;
  wire [6:0]  _slots_21_io_uop_prs2;
  wire [6:0]  _slots_21_io_uop_prs3;
  wire [5:0]  _slots_21_io_uop_ppred;
  wire        _slots_21_io_uop_prs1_busy;
  wire        _slots_21_io_uop_prs2_busy;
  wire        _slots_21_io_uop_prs3_busy;
  wire        _slots_21_io_uop_ppred_busy;
  wire [6:0]  _slots_21_io_uop_stale_pdst;
  wire        _slots_21_io_uop_exception;
  wire [63:0] _slots_21_io_uop_exc_cause;
  wire        _slots_21_io_uop_bypassable;
  wire [4:0]  _slots_21_io_uop_mem_cmd;
  wire [1:0]  _slots_21_io_uop_mem_size;
  wire        _slots_21_io_uop_mem_signed;
  wire        _slots_21_io_uop_is_fence;
  wire        _slots_21_io_uop_is_fencei;
  wire        _slots_21_io_uop_is_amo;
  wire        _slots_21_io_uop_uses_ldq;
  wire        _slots_21_io_uop_uses_stq;
  wire        _slots_21_io_uop_is_sys_pc2epc;
  wire        _slots_21_io_uop_is_unique;
  wire        _slots_21_io_uop_flush_on_commit;
  wire        _slots_21_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_21_io_uop_ldst;
  wire [5:0]  _slots_21_io_uop_lrs1;
  wire [5:0]  _slots_21_io_uop_lrs2;
  wire [5:0]  _slots_21_io_uop_lrs3;
  wire        _slots_21_io_uop_ldst_val;
  wire [1:0]  _slots_21_io_uop_dst_rtype;
  wire [1:0]  _slots_21_io_uop_lrs1_rtype;
  wire [1:0]  _slots_21_io_uop_lrs2_rtype;
  wire        _slots_21_io_uop_frs3_en;
  wire        _slots_21_io_uop_fp_val;
  wire        _slots_21_io_uop_fp_single;
  wire        _slots_21_io_uop_xcpt_pf_if;
  wire        _slots_21_io_uop_xcpt_ae_if;
  wire        _slots_21_io_uop_xcpt_ma_if;
  wire        _slots_21_io_uop_bp_debug_if;
  wire        _slots_21_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_21_io_uop_debug_fsrc;
  wire [1:0]  _slots_21_io_uop_debug_tsrc;
  wire        _slots_20_io_valid;
  wire        _slots_20_io_will_be_valid;
  wire        _slots_20_io_request;
  wire [6:0]  _slots_20_io_out_uop_uopc;
  wire [31:0] _slots_20_io_out_uop_inst;
  wire [31:0] _slots_20_io_out_uop_debug_inst;
  wire        _slots_20_io_out_uop_is_rvc;
  wire [39:0] _slots_20_io_out_uop_debug_pc;
  wire [2:0]  _slots_20_io_out_uop_iq_type;
  wire [9:0]  _slots_20_io_out_uop_fu_code;
  wire [1:0]  _slots_20_io_out_uop_iw_state;
  wire        _slots_20_io_out_uop_iw_p1_poisoned;
  wire        _slots_20_io_out_uop_iw_p2_poisoned;
  wire        _slots_20_io_out_uop_is_br;
  wire        _slots_20_io_out_uop_is_jalr;
  wire        _slots_20_io_out_uop_is_jal;
  wire        _slots_20_io_out_uop_is_sfb;
  wire [19:0] _slots_20_io_out_uop_br_mask;
  wire [4:0]  _slots_20_io_out_uop_br_tag;
  wire [5:0]  _slots_20_io_out_uop_ftq_idx;
  wire        _slots_20_io_out_uop_edge_inst;
  wire [5:0]  _slots_20_io_out_uop_pc_lob;
  wire        _slots_20_io_out_uop_taken;
  wire [19:0] _slots_20_io_out_uop_imm_packed;
  wire [11:0] _slots_20_io_out_uop_csr_addr;
  wire [6:0]  _slots_20_io_out_uop_rob_idx;
  wire [4:0]  _slots_20_io_out_uop_ldq_idx;
  wire [4:0]  _slots_20_io_out_uop_stq_idx;
  wire [1:0]  _slots_20_io_out_uop_rxq_idx;
  wire [6:0]  _slots_20_io_out_uop_pdst;
  wire [6:0]  _slots_20_io_out_uop_prs1;
  wire [6:0]  _slots_20_io_out_uop_prs2;
  wire [6:0]  _slots_20_io_out_uop_prs3;
  wire [5:0]  _slots_20_io_out_uop_ppred;
  wire        _slots_20_io_out_uop_prs1_busy;
  wire        _slots_20_io_out_uop_prs2_busy;
  wire        _slots_20_io_out_uop_prs3_busy;
  wire        _slots_20_io_out_uop_ppred_busy;
  wire [6:0]  _slots_20_io_out_uop_stale_pdst;
  wire        _slots_20_io_out_uop_exception;
  wire [63:0] _slots_20_io_out_uop_exc_cause;
  wire        _slots_20_io_out_uop_bypassable;
  wire [4:0]  _slots_20_io_out_uop_mem_cmd;
  wire [1:0]  _slots_20_io_out_uop_mem_size;
  wire        _slots_20_io_out_uop_mem_signed;
  wire        _slots_20_io_out_uop_is_fence;
  wire        _slots_20_io_out_uop_is_fencei;
  wire        _slots_20_io_out_uop_is_amo;
  wire        _slots_20_io_out_uop_uses_ldq;
  wire        _slots_20_io_out_uop_uses_stq;
  wire        _slots_20_io_out_uop_is_sys_pc2epc;
  wire        _slots_20_io_out_uop_is_unique;
  wire        _slots_20_io_out_uop_flush_on_commit;
  wire        _slots_20_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_20_io_out_uop_ldst;
  wire [5:0]  _slots_20_io_out_uop_lrs1;
  wire [5:0]  _slots_20_io_out_uop_lrs2;
  wire [5:0]  _slots_20_io_out_uop_lrs3;
  wire        _slots_20_io_out_uop_ldst_val;
  wire [1:0]  _slots_20_io_out_uop_dst_rtype;
  wire [1:0]  _slots_20_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_20_io_out_uop_lrs2_rtype;
  wire        _slots_20_io_out_uop_frs3_en;
  wire        _slots_20_io_out_uop_fp_val;
  wire        _slots_20_io_out_uop_fp_single;
  wire        _slots_20_io_out_uop_xcpt_pf_if;
  wire        _slots_20_io_out_uop_xcpt_ae_if;
  wire        _slots_20_io_out_uop_xcpt_ma_if;
  wire        _slots_20_io_out_uop_bp_debug_if;
  wire        _slots_20_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_20_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_20_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_20_io_uop_uopc;
  wire [31:0] _slots_20_io_uop_inst;
  wire [31:0] _slots_20_io_uop_debug_inst;
  wire        _slots_20_io_uop_is_rvc;
  wire [39:0] _slots_20_io_uop_debug_pc;
  wire [2:0]  _slots_20_io_uop_iq_type;
  wire [9:0]  _slots_20_io_uop_fu_code;
  wire [1:0]  _slots_20_io_uop_iw_state;
  wire        _slots_20_io_uop_iw_p1_poisoned;
  wire        _slots_20_io_uop_iw_p2_poisoned;
  wire        _slots_20_io_uop_is_br;
  wire        _slots_20_io_uop_is_jalr;
  wire        _slots_20_io_uop_is_jal;
  wire        _slots_20_io_uop_is_sfb;
  wire [19:0] _slots_20_io_uop_br_mask;
  wire [4:0]  _slots_20_io_uop_br_tag;
  wire [5:0]  _slots_20_io_uop_ftq_idx;
  wire        _slots_20_io_uop_edge_inst;
  wire [5:0]  _slots_20_io_uop_pc_lob;
  wire        _slots_20_io_uop_taken;
  wire [19:0] _slots_20_io_uop_imm_packed;
  wire [11:0] _slots_20_io_uop_csr_addr;
  wire [6:0]  _slots_20_io_uop_rob_idx;
  wire [4:0]  _slots_20_io_uop_ldq_idx;
  wire [4:0]  _slots_20_io_uop_stq_idx;
  wire [1:0]  _slots_20_io_uop_rxq_idx;
  wire [6:0]  _slots_20_io_uop_pdst;
  wire [6:0]  _slots_20_io_uop_prs1;
  wire [6:0]  _slots_20_io_uop_prs2;
  wire [6:0]  _slots_20_io_uop_prs3;
  wire [5:0]  _slots_20_io_uop_ppred;
  wire        _slots_20_io_uop_prs1_busy;
  wire        _slots_20_io_uop_prs2_busy;
  wire        _slots_20_io_uop_prs3_busy;
  wire        _slots_20_io_uop_ppred_busy;
  wire [6:0]  _slots_20_io_uop_stale_pdst;
  wire        _slots_20_io_uop_exception;
  wire [63:0] _slots_20_io_uop_exc_cause;
  wire        _slots_20_io_uop_bypassable;
  wire [4:0]  _slots_20_io_uop_mem_cmd;
  wire [1:0]  _slots_20_io_uop_mem_size;
  wire        _slots_20_io_uop_mem_signed;
  wire        _slots_20_io_uop_is_fence;
  wire        _slots_20_io_uop_is_fencei;
  wire        _slots_20_io_uop_is_amo;
  wire        _slots_20_io_uop_uses_ldq;
  wire        _slots_20_io_uop_uses_stq;
  wire        _slots_20_io_uop_is_sys_pc2epc;
  wire        _slots_20_io_uop_is_unique;
  wire        _slots_20_io_uop_flush_on_commit;
  wire        _slots_20_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_20_io_uop_ldst;
  wire [5:0]  _slots_20_io_uop_lrs1;
  wire [5:0]  _slots_20_io_uop_lrs2;
  wire [5:0]  _slots_20_io_uop_lrs3;
  wire        _slots_20_io_uop_ldst_val;
  wire [1:0]  _slots_20_io_uop_dst_rtype;
  wire [1:0]  _slots_20_io_uop_lrs1_rtype;
  wire [1:0]  _slots_20_io_uop_lrs2_rtype;
  wire        _slots_20_io_uop_frs3_en;
  wire        _slots_20_io_uop_fp_val;
  wire        _slots_20_io_uop_fp_single;
  wire        _slots_20_io_uop_xcpt_pf_if;
  wire        _slots_20_io_uop_xcpt_ae_if;
  wire        _slots_20_io_uop_xcpt_ma_if;
  wire        _slots_20_io_uop_bp_debug_if;
  wire        _slots_20_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_20_io_uop_debug_fsrc;
  wire [1:0]  _slots_20_io_uop_debug_tsrc;
  wire        _slots_19_io_valid;
  wire        _slots_19_io_will_be_valid;
  wire        _slots_19_io_request;
  wire [6:0]  _slots_19_io_out_uop_uopc;
  wire [31:0] _slots_19_io_out_uop_inst;
  wire [31:0] _slots_19_io_out_uop_debug_inst;
  wire        _slots_19_io_out_uop_is_rvc;
  wire [39:0] _slots_19_io_out_uop_debug_pc;
  wire [2:0]  _slots_19_io_out_uop_iq_type;
  wire [9:0]  _slots_19_io_out_uop_fu_code;
  wire [1:0]  _slots_19_io_out_uop_iw_state;
  wire        _slots_19_io_out_uop_iw_p1_poisoned;
  wire        _slots_19_io_out_uop_iw_p2_poisoned;
  wire        _slots_19_io_out_uop_is_br;
  wire        _slots_19_io_out_uop_is_jalr;
  wire        _slots_19_io_out_uop_is_jal;
  wire        _slots_19_io_out_uop_is_sfb;
  wire [19:0] _slots_19_io_out_uop_br_mask;
  wire [4:0]  _slots_19_io_out_uop_br_tag;
  wire [5:0]  _slots_19_io_out_uop_ftq_idx;
  wire        _slots_19_io_out_uop_edge_inst;
  wire [5:0]  _slots_19_io_out_uop_pc_lob;
  wire        _slots_19_io_out_uop_taken;
  wire [19:0] _slots_19_io_out_uop_imm_packed;
  wire [11:0] _slots_19_io_out_uop_csr_addr;
  wire [6:0]  _slots_19_io_out_uop_rob_idx;
  wire [4:0]  _slots_19_io_out_uop_ldq_idx;
  wire [4:0]  _slots_19_io_out_uop_stq_idx;
  wire [1:0]  _slots_19_io_out_uop_rxq_idx;
  wire [6:0]  _slots_19_io_out_uop_pdst;
  wire [6:0]  _slots_19_io_out_uop_prs1;
  wire [6:0]  _slots_19_io_out_uop_prs2;
  wire [6:0]  _slots_19_io_out_uop_prs3;
  wire [5:0]  _slots_19_io_out_uop_ppred;
  wire        _slots_19_io_out_uop_prs1_busy;
  wire        _slots_19_io_out_uop_prs2_busy;
  wire        _slots_19_io_out_uop_prs3_busy;
  wire        _slots_19_io_out_uop_ppred_busy;
  wire [6:0]  _slots_19_io_out_uop_stale_pdst;
  wire        _slots_19_io_out_uop_exception;
  wire [63:0] _slots_19_io_out_uop_exc_cause;
  wire        _slots_19_io_out_uop_bypassable;
  wire [4:0]  _slots_19_io_out_uop_mem_cmd;
  wire [1:0]  _slots_19_io_out_uop_mem_size;
  wire        _slots_19_io_out_uop_mem_signed;
  wire        _slots_19_io_out_uop_is_fence;
  wire        _slots_19_io_out_uop_is_fencei;
  wire        _slots_19_io_out_uop_is_amo;
  wire        _slots_19_io_out_uop_uses_ldq;
  wire        _slots_19_io_out_uop_uses_stq;
  wire        _slots_19_io_out_uop_is_sys_pc2epc;
  wire        _slots_19_io_out_uop_is_unique;
  wire        _slots_19_io_out_uop_flush_on_commit;
  wire        _slots_19_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_19_io_out_uop_ldst;
  wire [5:0]  _slots_19_io_out_uop_lrs1;
  wire [5:0]  _slots_19_io_out_uop_lrs2;
  wire [5:0]  _slots_19_io_out_uop_lrs3;
  wire        _slots_19_io_out_uop_ldst_val;
  wire [1:0]  _slots_19_io_out_uop_dst_rtype;
  wire [1:0]  _slots_19_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_19_io_out_uop_lrs2_rtype;
  wire        _slots_19_io_out_uop_frs3_en;
  wire        _slots_19_io_out_uop_fp_val;
  wire        _slots_19_io_out_uop_fp_single;
  wire        _slots_19_io_out_uop_xcpt_pf_if;
  wire        _slots_19_io_out_uop_xcpt_ae_if;
  wire        _slots_19_io_out_uop_xcpt_ma_if;
  wire        _slots_19_io_out_uop_bp_debug_if;
  wire        _slots_19_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_19_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_19_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_19_io_uop_uopc;
  wire [31:0] _slots_19_io_uop_inst;
  wire [31:0] _slots_19_io_uop_debug_inst;
  wire        _slots_19_io_uop_is_rvc;
  wire [39:0] _slots_19_io_uop_debug_pc;
  wire [2:0]  _slots_19_io_uop_iq_type;
  wire [9:0]  _slots_19_io_uop_fu_code;
  wire [1:0]  _slots_19_io_uop_iw_state;
  wire        _slots_19_io_uop_iw_p1_poisoned;
  wire        _slots_19_io_uop_iw_p2_poisoned;
  wire        _slots_19_io_uop_is_br;
  wire        _slots_19_io_uop_is_jalr;
  wire        _slots_19_io_uop_is_jal;
  wire        _slots_19_io_uop_is_sfb;
  wire [19:0] _slots_19_io_uop_br_mask;
  wire [4:0]  _slots_19_io_uop_br_tag;
  wire [5:0]  _slots_19_io_uop_ftq_idx;
  wire        _slots_19_io_uop_edge_inst;
  wire [5:0]  _slots_19_io_uop_pc_lob;
  wire        _slots_19_io_uop_taken;
  wire [19:0] _slots_19_io_uop_imm_packed;
  wire [11:0] _slots_19_io_uop_csr_addr;
  wire [6:0]  _slots_19_io_uop_rob_idx;
  wire [4:0]  _slots_19_io_uop_ldq_idx;
  wire [4:0]  _slots_19_io_uop_stq_idx;
  wire [1:0]  _slots_19_io_uop_rxq_idx;
  wire [6:0]  _slots_19_io_uop_pdst;
  wire [6:0]  _slots_19_io_uop_prs1;
  wire [6:0]  _slots_19_io_uop_prs2;
  wire [6:0]  _slots_19_io_uop_prs3;
  wire [5:0]  _slots_19_io_uop_ppred;
  wire        _slots_19_io_uop_prs1_busy;
  wire        _slots_19_io_uop_prs2_busy;
  wire        _slots_19_io_uop_prs3_busy;
  wire        _slots_19_io_uop_ppred_busy;
  wire [6:0]  _slots_19_io_uop_stale_pdst;
  wire        _slots_19_io_uop_exception;
  wire [63:0] _slots_19_io_uop_exc_cause;
  wire        _slots_19_io_uop_bypassable;
  wire [4:0]  _slots_19_io_uop_mem_cmd;
  wire [1:0]  _slots_19_io_uop_mem_size;
  wire        _slots_19_io_uop_mem_signed;
  wire        _slots_19_io_uop_is_fence;
  wire        _slots_19_io_uop_is_fencei;
  wire        _slots_19_io_uop_is_amo;
  wire        _slots_19_io_uop_uses_ldq;
  wire        _slots_19_io_uop_uses_stq;
  wire        _slots_19_io_uop_is_sys_pc2epc;
  wire        _slots_19_io_uop_is_unique;
  wire        _slots_19_io_uop_flush_on_commit;
  wire        _slots_19_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_19_io_uop_ldst;
  wire [5:0]  _slots_19_io_uop_lrs1;
  wire [5:0]  _slots_19_io_uop_lrs2;
  wire [5:0]  _slots_19_io_uop_lrs3;
  wire        _slots_19_io_uop_ldst_val;
  wire [1:0]  _slots_19_io_uop_dst_rtype;
  wire [1:0]  _slots_19_io_uop_lrs1_rtype;
  wire [1:0]  _slots_19_io_uop_lrs2_rtype;
  wire        _slots_19_io_uop_frs3_en;
  wire        _slots_19_io_uop_fp_val;
  wire        _slots_19_io_uop_fp_single;
  wire        _slots_19_io_uop_xcpt_pf_if;
  wire        _slots_19_io_uop_xcpt_ae_if;
  wire        _slots_19_io_uop_xcpt_ma_if;
  wire        _slots_19_io_uop_bp_debug_if;
  wire        _slots_19_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_19_io_uop_debug_fsrc;
  wire [1:0]  _slots_19_io_uop_debug_tsrc;
  wire        _slots_18_io_valid;
  wire        _slots_18_io_will_be_valid;
  wire        _slots_18_io_request;
  wire [6:0]  _slots_18_io_out_uop_uopc;
  wire [31:0] _slots_18_io_out_uop_inst;
  wire [31:0] _slots_18_io_out_uop_debug_inst;
  wire        _slots_18_io_out_uop_is_rvc;
  wire [39:0] _slots_18_io_out_uop_debug_pc;
  wire [2:0]  _slots_18_io_out_uop_iq_type;
  wire [9:0]  _slots_18_io_out_uop_fu_code;
  wire [1:0]  _slots_18_io_out_uop_iw_state;
  wire        _slots_18_io_out_uop_iw_p1_poisoned;
  wire        _slots_18_io_out_uop_iw_p2_poisoned;
  wire        _slots_18_io_out_uop_is_br;
  wire        _slots_18_io_out_uop_is_jalr;
  wire        _slots_18_io_out_uop_is_jal;
  wire        _slots_18_io_out_uop_is_sfb;
  wire [19:0] _slots_18_io_out_uop_br_mask;
  wire [4:0]  _slots_18_io_out_uop_br_tag;
  wire [5:0]  _slots_18_io_out_uop_ftq_idx;
  wire        _slots_18_io_out_uop_edge_inst;
  wire [5:0]  _slots_18_io_out_uop_pc_lob;
  wire        _slots_18_io_out_uop_taken;
  wire [19:0] _slots_18_io_out_uop_imm_packed;
  wire [11:0] _slots_18_io_out_uop_csr_addr;
  wire [6:0]  _slots_18_io_out_uop_rob_idx;
  wire [4:0]  _slots_18_io_out_uop_ldq_idx;
  wire [4:0]  _slots_18_io_out_uop_stq_idx;
  wire [1:0]  _slots_18_io_out_uop_rxq_idx;
  wire [6:0]  _slots_18_io_out_uop_pdst;
  wire [6:0]  _slots_18_io_out_uop_prs1;
  wire [6:0]  _slots_18_io_out_uop_prs2;
  wire [6:0]  _slots_18_io_out_uop_prs3;
  wire [5:0]  _slots_18_io_out_uop_ppred;
  wire        _slots_18_io_out_uop_prs1_busy;
  wire        _slots_18_io_out_uop_prs2_busy;
  wire        _slots_18_io_out_uop_prs3_busy;
  wire        _slots_18_io_out_uop_ppred_busy;
  wire [6:0]  _slots_18_io_out_uop_stale_pdst;
  wire        _slots_18_io_out_uop_exception;
  wire [63:0] _slots_18_io_out_uop_exc_cause;
  wire        _slots_18_io_out_uop_bypassable;
  wire [4:0]  _slots_18_io_out_uop_mem_cmd;
  wire [1:0]  _slots_18_io_out_uop_mem_size;
  wire        _slots_18_io_out_uop_mem_signed;
  wire        _slots_18_io_out_uop_is_fence;
  wire        _slots_18_io_out_uop_is_fencei;
  wire        _slots_18_io_out_uop_is_amo;
  wire        _slots_18_io_out_uop_uses_ldq;
  wire        _slots_18_io_out_uop_uses_stq;
  wire        _slots_18_io_out_uop_is_sys_pc2epc;
  wire        _slots_18_io_out_uop_is_unique;
  wire        _slots_18_io_out_uop_flush_on_commit;
  wire        _slots_18_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_18_io_out_uop_ldst;
  wire [5:0]  _slots_18_io_out_uop_lrs1;
  wire [5:0]  _slots_18_io_out_uop_lrs2;
  wire [5:0]  _slots_18_io_out_uop_lrs3;
  wire        _slots_18_io_out_uop_ldst_val;
  wire [1:0]  _slots_18_io_out_uop_dst_rtype;
  wire [1:0]  _slots_18_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_18_io_out_uop_lrs2_rtype;
  wire        _slots_18_io_out_uop_frs3_en;
  wire        _slots_18_io_out_uop_fp_val;
  wire        _slots_18_io_out_uop_fp_single;
  wire        _slots_18_io_out_uop_xcpt_pf_if;
  wire        _slots_18_io_out_uop_xcpt_ae_if;
  wire        _slots_18_io_out_uop_xcpt_ma_if;
  wire        _slots_18_io_out_uop_bp_debug_if;
  wire        _slots_18_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_18_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_18_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_18_io_uop_uopc;
  wire [31:0] _slots_18_io_uop_inst;
  wire [31:0] _slots_18_io_uop_debug_inst;
  wire        _slots_18_io_uop_is_rvc;
  wire [39:0] _slots_18_io_uop_debug_pc;
  wire [2:0]  _slots_18_io_uop_iq_type;
  wire [9:0]  _slots_18_io_uop_fu_code;
  wire [1:0]  _slots_18_io_uop_iw_state;
  wire        _slots_18_io_uop_iw_p1_poisoned;
  wire        _slots_18_io_uop_iw_p2_poisoned;
  wire        _slots_18_io_uop_is_br;
  wire        _slots_18_io_uop_is_jalr;
  wire        _slots_18_io_uop_is_jal;
  wire        _slots_18_io_uop_is_sfb;
  wire [19:0] _slots_18_io_uop_br_mask;
  wire [4:0]  _slots_18_io_uop_br_tag;
  wire [5:0]  _slots_18_io_uop_ftq_idx;
  wire        _slots_18_io_uop_edge_inst;
  wire [5:0]  _slots_18_io_uop_pc_lob;
  wire        _slots_18_io_uop_taken;
  wire [19:0] _slots_18_io_uop_imm_packed;
  wire [11:0] _slots_18_io_uop_csr_addr;
  wire [6:0]  _slots_18_io_uop_rob_idx;
  wire [4:0]  _slots_18_io_uop_ldq_idx;
  wire [4:0]  _slots_18_io_uop_stq_idx;
  wire [1:0]  _slots_18_io_uop_rxq_idx;
  wire [6:0]  _slots_18_io_uop_pdst;
  wire [6:0]  _slots_18_io_uop_prs1;
  wire [6:0]  _slots_18_io_uop_prs2;
  wire [6:0]  _slots_18_io_uop_prs3;
  wire [5:0]  _slots_18_io_uop_ppred;
  wire        _slots_18_io_uop_prs1_busy;
  wire        _slots_18_io_uop_prs2_busy;
  wire        _slots_18_io_uop_prs3_busy;
  wire        _slots_18_io_uop_ppred_busy;
  wire [6:0]  _slots_18_io_uop_stale_pdst;
  wire        _slots_18_io_uop_exception;
  wire [63:0] _slots_18_io_uop_exc_cause;
  wire        _slots_18_io_uop_bypassable;
  wire [4:0]  _slots_18_io_uop_mem_cmd;
  wire [1:0]  _slots_18_io_uop_mem_size;
  wire        _slots_18_io_uop_mem_signed;
  wire        _slots_18_io_uop_is_fence;
  wire        _slots_18_io_uop_is_fencei;
  wire        _slots_18_io_uop_is_amo;
  wire        _slots_18_io_uop_uses_ldq;
  wire        _slots_18_io_uop_uses_stq;
  wire        _slots_18_io_uop_is_sys_pc2epc;
  wire        _slots_18_io_uop_is_unique;
  wire        _slots_18_io_uop_flush_on_commit;
  wire        _slots_18_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_18_io_uop_ldst;
  wire [5:0]  _slots_18_io_uop_lrs1;
  wire [5:0]  _slots_18_io_uop_lrs2;
  wire [5:0]  _slots_18_io_uop_lrs3;
  wire        _slots_18_io_uop_ldst_val;
  wire [1:0]  _slots_18_io_uop_dst_rtype;
  wire [1:0]  _slots_18_io_uop_lrs1_rtype;
  wire [1:0]  _slots_18_io_uop_lrs2_rtype;
  wire        _slots_18_io_uop_frs3_en;
  wire        _slots_18_io_uop_fp_val;
  wire        _slots_18_io_uop_fp_single;
  wire        _slots_18_io_uop_xcpt_pf_if;
  wire        _slots_18_io_uop_xcpt_ae_if;
  wire        _slots_18_io_uop_xcpt_ma_if;
  wire        _slots_18_io_uop_bp_debug_if;
  wire        _slots_18_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_18_io_uop_debug_fsrc;
  wire [1:0]  _slots_18_io_uop_debug_tsrc;
  wire        _slots_17_io_valid;
  wire        _slots_17_io_will_be_valid;
  wire        _slots_17_io_request;
  wire [6:0]  _slots_17_io_out_uop_uopc;
  wire [31:0] _slots_17_io_out_uop_inst;
  wire [31:0] _slots_17_io_out_uop_debug_inst;
  wire        _slots_17_io_out_uop_is_rvc;
  wire [39:0] _slots_17_io_out_uop_debug_pc;
  wire [2:0]  _slots_17_io_out_uop_iq_type;
  wire [9:0]  _slots_17_io_out_uop_fu_code;
  wire [1:0]  _slots_17_io_out_uop_iw_state;
  wire        _slots_17_io_out_uop_iw_p1_poisoned;
  wire        _slots_17_io_out_uop_iw_p2_poisoned;
  wire        _slots_17_io_out_uop_is_br;
  wire        _slots_17_io_out_uop_is_jalr;
  wire        _slots_17_io_out_uop_is_jal;
  wire        _slots_17_io_out_uop_is_sfb;
  wire [19:0] _slots_17_io_out_uop_br_mask;
  wire [4:0]  _slots_17_io_out_uop_br_tag;
  wire [5:0]  _slots_17_io_out_uop_ftq_idx;
  wire        _slots_17_io_out_uop_edge_inst;
  wire [5:0]  _slots_17_io_out_uop_pc_lob;
  wire        _slots_17_io_out_uop_taken;
  wire [19:0] _slots_17_io_out_uop_imm_packed;
  wire [11:0] _slots_17_io_out_uop_csr_addr;
  wire [6:0]  _slots_17_io_out_uop_rob_idx;
  wire [4:0]  _slots_17_io_out_uop_ldq_idx;
  wire [4:0]  _slots_17_io_out_uop_stq_idx;
  wire [1:0]  _slots_17_io_out_uop_rxq_idx;
  wire [6:0]  _slots_17_io_out_uop_pdst;
  wire [6:0]  _slots_17_io_out_uop_prs1;
  wire [6:0]  _slots_17_io_out_uop_prs2;
  wire [6:0]  _slots_17_io_out_uop_prs3;
  wire [5:0]  _slots_17_io_out_uop_ppred;
  wire        _slots_17_io_out_uop_prs1_busy;
  wire        _slots_17_io_out_uop_prs2_busy;
  wire        _slots_17_io_out_uop_prs3_busy;
  wire        _slots_17_io_out_uop_ppred_busy;
  wire [6:0]  _slots_17_io_out_uop_stale_pdst;
  wire        _slots_17_io_out_uop_exception;
  wire [63:0] _slots_17_io_out_uop_exc_cause;
  wire        _slots_17_io_out_uop_bypassable;
  wire [4:0]  _slots_17_io_out_uop_mem_cmd;
  wire [1:0]  _slots_17_io_out_uop_mem_size;
  wire        _slots_17_io_out_uop_mem_signed;
  wire        _slots_17_io_out_uop_is_fence;
  wire        _slots_17_io_out_uop_is_fencei;
  wire        _slots_17_io_out_uop_is_amo;
  wire        _slots_17_io_out_uop_uses_ldq;
  wire        _slots_17_io_out_uop_uses_stq;
  wire        _slots_17_io_out_uop_is_sys_pc2epc;
  wire        _slots_17_io_out_uop_is_unique;
  wire        _slots_17_io_out_uop_flush_on_commit;
  wire        _slots_17_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_17_io_out_uop_ldst;
  wire [5:0]  _slots_17_io_out_uop_lrs1;
  wire [5:0]  _slots_17_io_out_uop_lrs2;
  wire [5:0]  _slots_17_io_out_uop_lrs3;
  wire        _slots_17_io_out_uop_ldst_val;
  wire [1:0]  _slots_17_io_out_uop_dst_rtype;
  wire [1:0]  _slots_17_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_17_io_out_uop_lrs2_rtype;
  wire        _slots_17_io_out_uop_frs3_en;
  wire        _slots_17_io_out_uop_fp_val;
  wire        _slots_17_io_out_uop_fp_single;
  wire        _slots_17_io_out_uop_xcpt_pf_if;
  wire        _slots_17_io_out_uop_xcpt_ae_if;
  wire        _slots_17_io_out_uop_xcpt_ma_if;
  wire        _slots_17_io_out_uop_bp_debug_if;
  wire        _slots_17_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_17_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_17_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_17_io_uop_uopc;
  wire [31:0] _slots_17_io_uop_inst;
  wire [31:0] _slots_17_io_uop_debug_inst;
  wire        _slots_17_io_uop_is_rvc;
  wire [39:0] _slots_17_io_uop_debug_pc;
  wire [2:0]  _slots_17_io_uop_iq_type;
  wire [9:0]  _slots_17_io_uop_fu_code;
  wire [1:0]  _slots_17_io_uop_iw_state;
  wire        _slots_17_io_uop_iw_p1_poisoned;
  wire        _slots_17_io_uop_iw_p2_poisoned;
  wire        _slots_17_io_uop_is_br;
  wire        _slots_17_io_uop_is_jalr;
  wire        _slots_17_io_uop_is_jal;
  wire        _slots_17_io_uop_is_sfb;
  wire [19:0] _slots_17_io_uop_br_mask;
  wire [4:0]  _slots_17_io_uop_br_tag;
  wire [5:0]  _slots_17_io_uop_ftq_idx;
  wire        _slots_17_io_uop_edge_inst;
  wire [5:0]  _slots_17_io_uop_pc_lob;
  wire        _slots_17_io_uop_taken;
  wire [19:0] _slots_17_io_uop_imm_packed;
  wire [11:0] _slots_17_io_uop_csr_addr;
  wire [6:0]  _slots_17_io_uop_rob_idx;
  wire [4:0]  _slots_17_io_uop_ldq_idx;
  wire [4:0]  _slots_17_io_uop_stq_idx;
  wire [1:0]  _slots_17_io_uop_rxq_idx;
  wire [6:0]  _slots_17_io_uop_pdst;
  wire [6:0]  _slots_17_io_uop_prs1;
  wire [6:0]  _slots_17_io_uop_prs2;
  wire [6:0]  _slots_17_io_uop_prs3;
  wire [5:0]  _slots_17_io_uop_ppred;
  wire        _slots_17_io_uop_prs1_busy;
  wire        _slots_17_io_uop_prs2_busy;
  wire        _slots_17_io_uop_prs3_busy;
  wire        _slots_17_io_uop_ppred_busy;
  wire [6:0]  _slots_17_io_uop_stale_pdst;
  wire        _slots_17_io_uop_exception;
  wire [63:0] _slots_17_io_uop_exc_cause;
  wire        _slots_17_io_uop_bypassable;
  wire [4:0]  _slots_17_io_uop_mem_cmd;
  wire [1:0]  _slots_17_io_uop_mem_size;
  wire        _slots_17_io_uop_mem_signed;
  wire        _slots_17_io_uop_is_fence;
  wire        _slots_17_io_uop_is_fencei;
  wire        _slots_17_io_uop_is_amo;
  wire        _slots_17_io_uop_uses_ldq;
  wire        _slots_17_io_uop_uses_stq;
  wire        _slots_17_io_uop_is_sys_pc2epc;
  wire        _slots_17_io_uop_is_unique;
  wire        _slots_17_io_uop_flush_on_commit;
  wire        _slots_17_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_17_io_uop_ldst;
  wire [5:0]  _slots_17_io_uop_lrs1;
  wire [5:0]  _slots_17_io_uop_lrs2;
  wire [5:0]  _slots_17_io_uop_lrs3;
  wire        _slots_17_io_uop_ldst_val;
  wire [1:0]  _slots_17_io_uop_dst_rtype;
  wire [1:0]  _slots_17_io_uop_lrs1_rtype;
  wire [1:0]  _slots_17_io_uop_lrs2_rtype;
  wire        _slots_17_io_uop_frs3_en;
  wire        _slots_17_io_uop_fp_val;
  wire        _slots_17_io_uop_fp_single;
  wire        _slots_17_io_uop_xcpt_pf_if;
  wire        _slots_17_io_uop_xcpt_ae_if;
  wire        _slots_17_io_uop_xcpt_ma_if;
  wire        _slots_17_io_uop_bp_debug_if;
  wire        _slots_17_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_17_io_uop_debug_fsrc;
  wire [1:0]  _slots_17_io_uop_debug_tsrc;
  wire        _slots_16_io_valid;
  wire        _slots_16_io_will_be_valid;
  wire        _slots_16_io_request;
  wire [6:0]  _slots_16_io_out_uop_uopc;
  wire [31:0] _slots_16_io_out_uop_inst;
  wire [31:0] _slots_16_io_out_uop_debug_inst;
  wire        _slots_16_io_out_uop_is_rvc;
  wire [39:0] _slots_16_io_out_uop_debug_pc;
  wire [2:0]  _slots_16_io_out_uop_iq_type;
  wire [9:0]  _slots_16_io_out_uop_fu_code;
  wire [1:0]  _slots_16_io_out_uop_iw_state;
  wire        _slots_16_io_out_uop_iw_p1_poisoned;
  wire        _slots_16_io_out_uop_iw_p2_poisoned;
  wire        _slots_16_io_out_uop_is_br;
  wire        _slots_16_io_out_uop_is_jalr;
  wire        _slots_16_io_out_uop_is_jal;
  wire        _slots_16_io_out_uop_is_sfb;
  wire [19:0] _slots_16_io_out_uop_br_mask;
  wire [4:0]  _slots_16_io_out_uop_br_tag;
  wire [5:0]  _slots_16_io_out_uop_ftq_idx;
  wire        _slots_16_io_out_uop_edge_inst;
  wire [5:0]  _slots_16_io_out_uop_pc_lob;
  wire        _slots_16_io_out_uop_taken;
  wire [19:0] _slots_16_io_out_uop_imm_packed;
  wire [11:0] _slots_16_io_out_uop_csr_addr;
  wire [6:0]  _slots_16_io_out_uop_rob_idx;
  wire [4:0]  _slots_16_io_out_uop_ldq_idx;
  wire [4:0]  _slots_16_io_out_uop_stq_idx;
  wire [1:0]  _slots_16_io_out_uop_rxq_idx;
  wire [6:0]  _slots_16_io_out_uop_pdst;
  wire [6:0]  _slots_16_io_out_uop_prs1;
  wire [6:0]  _slots_16_io_out_uop_prs2;
  wire [6:0]  _slots_16_io_out_uop_prs3;
  wire [5:0]  _slots_16_io_out_uop_ppred;
  wire        _slots_16_io_out_uop_prs1_busy;
  wire        _slots_16_io_out_uop_prs2_busy;
  wire        _slots_16_io_out_uop_prs3_busy;
  wire        _slots_16_io_out_uop_ppred_busy;
  wire [6:0]  _slots_16_io_out_uop_stale_pdst;
  wire        _slots_16_io_out_uop_exception;
  wire [63:0] _slots_16_io_out_uop_exc_cause;
  wire        _slots_16_io_out_uop_bypassable;
  wire [4:0]  _slots_16_io_out_uop_mem_cmd;
  wire [1:0]  _slots_16_io_out_uop_mem_size;
  wire        _slots_16_io_out_uop_mem_signed;
  wire        _slots_16_io_out_uop_is_fence;
  wire        _slots_16_io_out_uop_is_fencei;
  wire        _slots_16_io_out_uop_is_amo;
  wire        _slots_16_io_out_uop_uses_ldq;
  wire        _slots_16_io_out_uop_uses_stq;
  wire        _slots_16_io_out_uop_is_sys_pc2epc;
  wire        _slots_16_io_out_uop_is_unique;
  wire        _slots_16_io_out_uop_flush_on_commit;
  wire        _slots_16_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_16_io_out_uop_ldst;
  wire [5:0]  _slots_16_io_out_uop_lrs1;
  wire [5:0]  _slots_16_io_out_uop_lrs2;
  wire [5:0]  _slots_16_io_out_uop_lrs3;
  wire        _slots_16_io_out_uop_ldst_val;
  wire [1:0]  _slots_16_io_out_uop_dst_rtype;
  wire [1:0]  _slots_16_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_16_io_out_uop_lrs2_rtype;
  wire        _slots_16_io_out_uop_frs3_en;
  wire        _slots_16_io_out_uop_fp_val;
  wire        _slots_16_io_out_uop_fp_single;
  wire        _slots_16_io_out_uop_xcpt_pf_if;
  wire        _slots_16_io_out_uop_xcpt_ae_if;
  wire        _slots_16_io_out_uop_xcpt_ma_if;
  wire        _slots_16_io_out_uop_bp_debug_if;
  wire        _slots_16_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_16_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_16_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_16_io_uop_uopc;
  wire [31:0] _slots_16_io_uop_inst;
  wire [31:0] _slots_16_io_uop_debug_inst;
  wire        _slots_16_io_uop_is_rvc;
  wire [39:0] _slots_16_io_uop_debug_pc;
  wire [2:0]  _slots_16_io_uop_iq_type;
  wire [9:0]  _slots_16_io_uop_fu_code;
  wire [1:0]  _slots_16_io_uop_iw_state;
  wire        _slots_16_io_uop_iw_p1_poisoned;
  wire        _slots_16_io_uop_iw_p2_poisoned;
  wire        _slots_16_io_uop_is_br;
  wire        _slots_16_io_uop_is_jalr;
  wire        _slots_16_io_uop_is_jal;
  wire        _slots_16_io_uop_is_sfb;
  wire [19:0] _slots_16_io_uop_br_mask;
  wire [4:0]  _slots_16_io_uop_br_tag;
  wire [5:0]  _slots_16_io_uop_ftq_idx;
  wire        _slots_16_io_uop_edge_inst;
  wire [5:0]  _slots_16_io_uop_pc_lob;
  wire        _slots_16_io_uop_taken;
  wire [19:0] _slots_16_io_uop_imm_packed;
  wire [11:0] _slots_16_io_uop_csr_addr;
  wire [6:0]  _slots_16_io_uop_rob_idx;
  wire [4:0]  _slots_16_io_uop_ldq_idx;
  wire [4:0]  _slots_16_io_uop_stq_idx;
  wire [1:0]  _slots_16_io_uop_rxq_idx;
  wire [6:0]  _slots_16_io_uop_pdst;
  wire [6:0]  _slots_16_io_uop_prs1;
  wire [6:0]  _slots_16_io_uop_prs2;
  wire [6:0]  _slots_16_io_uop_prs3;
  wire [5:0]  _slots_16_io_uop_ppred;
  wire        _slots_16_io_uop_prs1_busy;
  wire        _slots_16_io_uop_prs2_busy;
  wire        _slots_16_io_uop_prs3_busy;
  wire        _slots_16_io_uop_ppred_busy;
  wire [6:0]  _slots_16_io_uop_stale_pdst;
  wire        _slots_16_io_uop_exception;
  wire [63:0] _slots_16_io_uop_exc_cause;
  wire        _slots_16_io_uop_bypassable;
  wire [4:0]  _slots_16_io_uop_mem_cmd;
  wire [1:0]  _slots_16_io_uop_mem_size;
  wire        _slots_16_io_uop_mem_signed;
  wire        _slots_16_io_uop_is_fence;
  wire        _slots_16_io_uop_is_fencei;
  wire        _slots_16_io_uop_is_amo;
  wire        _slots_16_io_uop_uses_ldq;
  wire        _slots_16_io_uop_uses_stq;
  wire        _slots_16_io_uop_is_sys_pc2epc;
  wire        _slots_16_io_uop_is_unique;
  wire        _slots_16_io_uop_flush_on_commit;
  wire        _slots_16_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_16_io_uop_ldst;
  wire [5:0]  _slots_16_io_uop_lrs1;
  wire [5:0]  _slots_16_io_uop_lrs2;
  wire [5:0]  _slots_16_io_uop_lrs3;
  wire        _slots_16_io_uop_ldst_val;
  wire [1:0]  _slots_16_io_uop_dst_rtype;
  wire [1:0]  _slots_16_io_uop_lrs1_rtype;
  wire [1:0]  _slots_16_io_uop_lrs2_rtype;
  wire        _slots_16_io_uop_frs3_en;
  wire        _slots_16_io_uop_fp_val;
  wire        _slots_16_io_uop_fp_single;
  wire        _slots_16_io_uop_xcpt_pf_if;
  wire        _slots_16_io_uop_xcpt_ae_if;
  wire        _slots_16_io_uop_xcpt_ma_if;
  wire        _slots_16_io_uop_bp_debug_if;
  wire        _slots_16_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_16_io_uop_debug_fsrc;
  wire [1:0]  _slots_16_io_uop_debug_tsrc;
  wire        _slots_15_io_valid;
  wire        _slots_15_io_will_be_valid;
  wire        _slots_15_io_request;
  wire [6:0]  _slots_15_io_out_uop_uopc;
  wire [31:0] _slots_15_io_out_uop_inst;
  wire [31:0] _slots_15_io_out_uop_debug_inst;
  wire        _slots_15_io_out_uop_is_rvc;
  wire [39:0] _slots_15_io_out_uop_debug_pc;
  wire [2:0]  _slots_15_io_out_uop_iq_type;
  wire [9:0]  _slots_15_io_out_uop_fu_code;
  wire [1:0]  _slots_15_io_out_uop_iw_state;
  wire        _slots_15_io_out_uop_iw_p1_poisoned;
  wire        _slots_15_io_out_uop_iw_p2_poisoned;
  wire        _slots_15_io_out_uop_is_br;
  wire        _slots_15_io_out_uop_is_jalr;
  wire        _slots_15_io_out_uop_is_jal;
  wire        _slots_15_io_out_uop_is_sfb;
  wire [19:0] _slots_15_io_out_uop_br_mask;
  wire [4:0]  _slots_15_io_out_uop_br_tag;
  wire [5:0]  _slots_15_io_out_uop_ftq_idx;
  wire        _slots_15_io_out_uop_edge_inst;
  wire [5:0]  _slots_15_io_out_uop_pc_lob;
  wire        _slots_15_io_out_uop_taken;
  wire [19:0] _slots_15_io_out_uop_imm_packed;
  wire [11:0] _slots_15_io_out_uop_csr_addr;
  wire [6:0]  _slots_15_io_out_uop_rob_idx;
  wire [4:0]  _slots_15_io_out_uop_ldq_idx;
  wire [4:0]  _slots_15_io_out_uop_stq_idx;
  wire [1:0]  _slots_15_io_out_uop_rxq_idx;
  wire [6:0]  _slots_15_io_out_uop_pdst;
  wire [6:0]  _slots_15_io_out_uop_prs1;
  wire [6:0]  _slots_15_io_out_uop_prs2;
  wire [6:0]  _slots_15_io_out_uop_prs3;
  wire [5:0]  _slots_15_io_out_uop_ppred;
  wire        _slots_15_io_out_uop_prs1_busy;
  wire        _slots_15_io_out_uop_prs2_busy;
  wire        _slots_15_io_out_uop_prs3_busy;
  wire        _slots_15_io_out_uop_ppred_busy;
  wire [6:0]  _slots_15_io_out_uop_stale_pdst;
  wire        _slots_15_io_out_uop_exception;
  wire [63:0] _slots_15_io_out_uop_exc_cause;
  wire        _slots_15_io_out_uop_bypassable;
  wire [4:0]  _slots_15_io_out_uop_mem_cmd;
  wire [1:0]  _slots_15_io_out_uop_mem_size;
  wire        _slots_15_io_out_uop_mem_signed;
  wire        _slots_15_io_out_uop_is_fence;
  wire        _slots_15_io_out_uop_is_fencei;
  wire        _slots_15_io_out_uop_is_amo;
  wire        _slots_15_io_out_uop_uses_ldq;
  wire        _slots_15_io_out_uop_uses_stq;
  wire        _slots_15_io_out_uop_is_sys_pc2epc;
  wire        _slots_15_io_out_uop_is_unique;
  wire        _slots_15_io_out_uop_flush_on_commit;
  wire        _slots_15_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_15_io_out_uop_ldst;
  wire [5:0]  _slots_15_io_out_uop_lrs1;
  wire [5:0]  _slots_15_io_out_uop_lrs2;
  wire [5:0]  _slots_15_io_out_uop_lrs3;
  wire        _slots_15_io_out_uop_ldst_val;
  wire [1:0]  _slots_15_io_out_uop_dst_rtype;
  wire [1:0]  _slots_15_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_15_io_out_uop_lrs2_rtype;
  wire        _slots_15_io_out_uop_frs3_en;
  wire        _slots_15_io_out_uop_fp_val;
  wire        _slots_15_io_out_uop_fp_single;
  wire        _slots_15_io_out_uop_xcpt_pf_if;
  wire        _slots_15_io_out_uop_xcpt_ae_if;
  wire        _slots_15_io_out_uop_xcpt_ma_if;
  wire        _slots_15_io_out_uop_bp_debug_if;
  wire        _slots_15_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_15_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_15_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_15_io_uop_uopc;
  wire [31:0] _slots_15_io_uop_inst;
  wire [31:0] _slots_15_io_uop_debug_inst;
  wire        _slots_15_io_uop_is_rvc;
  wire [39:0] _slots_15_io_uop_debug_pc;
  wire [2:0]  _slots_15_io_uop_iq_type;
  wire [9:0]  _slots_15_io_uop_fu_code;
  wire [1:0]  _slots_15_io_uop_iw_state;
  wire        _slots_15_io_uop_iw_p1_poisoned;
  wire        _slots_15_io_uop_iw_p2_poisoned;
  wire        _slots_15_io_uop_is_br;
  wire        _slots_15_io_uop_is_jalr;
  wire        _slots_15_io_uop_is_jal;
  wire        _slots_15_io_uop_is_sfb;
  wire [19:0] _slots_15_io_uop_br_mask;
  wire [4:0]  _slots_15_io_uop_br_tag;
  wire [5:0]  _slots_15_io_uop_ftq_idx;
  wire        _slots_15_io_uop_edge_inst;
  wire [5:0]  _slots_15_io_uop_pc_lob;
  wire        _slots_15_io_uop_taken;
  wire [19:0] _slots_15_io_uop_imm_packed;
  wire [11:0] _slots_15_io_uop_csr_addr;
  wire [6:0]  _slots_15_io_uop_rob_idx;
  wire [4:0]  _slots_15_io_uop_ldq_idx;
  wire [4:0]  _slots_15_io_uop_stq_idx;
  wire [1:0]  _slots_15_io_uop_rxq_idx;
  wire [6:0]  _slots_15_io_uop_pdst;
  wire [6:0]  _slots_15_io_uop_prs1;
  wire [6:0]  _slots_15_io_uop_prs2;
  wire [6:0]  _slots_15_io_uop_prs3;
  wire [5:0]  _slots_15_io_uop_ppred;
  wire        _slots_15_io_uop_prs1_busy;
  wire        _slots_15_io_uop_prs2_busy;
  wire        _slots_15_io_uop_prs3_busy;
  wire        _slots_15_io_uop_ppred_busy;
  wire [6:0]  _slots_15_io_uop_stale_pdst;
  wire        _slots_15_io_uop_exception;
  wire [63:0] _slots_15_io_uop_exc_cause;
  wire        _slots_15_io_uop_bypassable;
  wire [4:0]  _slots_15_io_uop_mem_cmd;
  wire [1:0]  _slots_15_io_uop_mem_size;
  wire        _slots_15_io_uop_mem_signed;
  wire        _slots_15_io_uop_is_fence;
  wire        _slots_15_io_uop_is_fencei;
  wire        _slots_15_io_uop_is_amo;
  wire        _slots_15_io_uop_uses_ldq;
  wire        _slots_15_io_uop_uses_stq;
  wire        _slots_15_io_uop_is_sys_pc2epc;
  wire        _slots_15_io_uop_is_unique;
  wire        _slots_15_io_uop_flush_on_commit;
  wire        _slots_15_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_15_io_uop_ldst;
  wire [5:0]  _slots_15_io_uop_lrs1;
  wire [5:0]  _slots_15_io_uop_lrs2;
  wire [5:0]  _slots_15_io_uop_lrs3;
  wire        _slots_15_io_uop_ldst_val;
  wire [1:0]  _slots_15_io_uop_dst_rtype;
  wire [1:0]  _slots_15_io_uop_lrs1_rtype;
  wire [1:0]  _slots_15_io_uop_lrs2_rtype;
  wire        _slots_15_io_uop_frs3_en;
  wire        _slots_15_io_uop_fp_val;
  wire        _slots_15_io_uop_fp_single;
  wire        _slots_15_io_uop_xcpt_pf_if;
  wire        _slots_15_io_uop_xcpt_ae_if;
  wire        _slots_15_io_uop_xcpt_ma_if;
  wire        _slots_15_io_uop_bp_debug_if;
  wire        _slots_15_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_15_io_uop_debug_fsrc;
  wire [1:0]  _slots_15_io_uop_debug_tsrc;
  wire        _slots_14_io_valid;
  wire        _slots_14_io_will_be_valid;
  wire        _slots_14_io_request;
  wire [6:0]  _slots_14_io_out_uop_uopc;
  wire [31:0] _slots_14_io_out_uop_inst;
  wire [31:0] _slots_14_io_out_uop_debug_inst;
  wire        _slots_14_io_out_uop_is_rvc;
  wire [39:0] _slots_14_io_out_uop_debug_pc;
  wire [2:0]  _slots_14_io_out_uop_iq_type;
  wire [9:0]  _slots_14_io_out_uop_fu_code;
  wire [1:0]  _slots_14_io_out_uop_iw_state;
  wire        _slots_14_io_out_uop_iw_p1_poisoned;
  wire        _slots_14_io_out_uop_iw_p2_poisoned;
  wire        _slots_14_io_out_uop_is_br;
  wire        _slots_14_io_out_uop_is_jalr;
  wire        _slots_14_io_out_uop_is_jal;
  wire        _slots_14_io_out_uop_is_sfb;
  wire [19:0] _slots_14_io_out_uop_br_mask;
  wire [4:0]  _slots_14_io_out_uop_br_tag;
  wire [5:0]  _slots_14_io_out_uop_ftq_idx;
  wire        _slots_14_io_out_uop_edge_inst;
  wire [5:0]  _slots_14_io_out_uop_pc_lob;
  wire        _slots_14_io_out_uop_taken;
  wire [19:0] _slots_14_io_out_uop_imm_packed;
  wire [11:0] _slots_14_io_out_uop_csr_addr;
  wire [6:0]  _slots_14_io_out_uop_rob_idx;
  wire [4:0]  _slots_14_io_out_uop_ldq_idx;
  wire [4:0]  _slots_14_io_out_uop_stq_idx;
  wire [1:0]  _slots_14_io_out_uop_rxq_idx;
  wire [6:0]  _slots_14_io_out_uop_pdst;
  wire [6:0]  _slots_14_io_out_uop_prs1;
  wire [6:0]  _slots_14_io_out_uop_prs2;
  wire [6:0]  _slots_14_io_out_uop_prs3;
  wire [5:0]  _slots_14_io_out_uop_ppred;
  wire        _slots_14_io_out_uop_prs1_busy;
  wire        _slots_14_io_out_uop_prs2_busy;
  wire        _slots_14_io_out_uop_prs3_busy;
  wire        _slots_14_io_out_uop_ppred_busy;
  wire [6:0]  _slots_14_io_out_uop_stale_pdst;
  wire        _slots_14_io_out_uop_exception;
  wire [63:0] _slots_14_io_out_uop_exc_cause;
  wire        _slots_14_io_out_uop_bypassable;
  wire [4:0]  _slots_14_io_out_uop_mem_cmd;
  wire [1:0]  _slots_14_io_out_uop_mem_size;
  wire        _slots_14_io_out_uop_mem_signed;
  wire        _slots_14_io_out_uop_is_fence;
  wire        _slots_14_io_out_uop_is_fencei;
  wire        _slots_14_io_out_uop_is_amo;
  wire        _slots_14_io_out_uop_uses_ldq;
  wire        _slots_14_io_out_uop_uses_stq;
  wire        _slots_14_io_out_uop_is_sys_pc2epc;
  wire        _slots_14_io_out_uop_is_unique;
  wire        _slots_14_io_out_uop_flush_on_commit;
  wire        _slots_14_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_14_io_out_uop_ldst;
  wire [5:0]  _slots_14_io_out_uop_lrs1;
  wire [5:0]  _slots_14_io_out_uop_lrs2;
  wire [5:0]  _slots_14_io_out_uop_lrs3;
  wire        _slots_14_io_out_uop_ldst_val;
  wire [1:0]  _slots_14_io_out_uop_dst_rtype;
  wire [1:0]  _slots_14_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_14_io_out_uop_lrs2_rtype;
  wire        _slots_14_io_out_uop_frs3_en;
  wire        _slots_14_io_out_uop_fp_val;
  wire        _slots_14_io_out_uop_fp_single;
  wire        _slots_14_io_out_uop_xcpt_pf_if;
  wire        _slots_14_io_out_uop_xcpt_ae_if;
  wire        _slots_14_io_out_uop_xcpt_ma_if;
  wire        _slots_14_io_out_uop_bp_debug_if;
  wire        _slots_14_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_14_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_14_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_14_io_uop_uopc;
  wire [31:0] _slots_14_io_uop_inst;
  wire [31:0] _slots_14_io_uop_debug_inst;
  wire        _slots_14_io_uop_is_rvc;
  wire [39:0] _slots_14_io_uop_debug_pc;
  wire [2:0]  _slots_14_io_uop_iq_type;
  wire [9:0]  _slots_14_io_uop_fu_code;
  wire [1:0]  _slots_14_io_uop_iw_state;
  wire        _slots_14_io_uop_iw_p1_poisoned;
  wire        _slots_14_io_uop_iw_p2_poisoned;
  wire        _slots_14_io_uop_is_br;
  wire        _slots_14_io_uop_is_jalr;
  wire        _slots_14_io_uop_is_jal;
  wire        _slots_14_io_uop_is_sfb;
  wire [19:0] _slots_14_io_uop_br_mask;
  wire [4:0]  _slots_14_io_uop_br_tag;
  wire [5:0]  _slots_14_io_uop_ftq_idx;
  wire        _slots_14_io_uop_edge_inst;
  wire [5:0]  _slots_14_io_uop_pc_lob;
  wire        _slots_14_io_uop_taken;
  wire [19:0] _slots_14_io_uop_imm_packed;
  wire [11:0] _slots_14_io_uop_csr_addr;
  wire [6:0]  _slots_14_io_uop_rob_idx;
  wire [4:0]  _slots_14_io_uop_ldq_idx;
  wire [4:0]  _slots_14_io_uop_stq_idx;
  wire [1:0]  _slots_14_io_uop_rxq_idx;
  wire [6:0]  _slots_14_io_uop_pdst;
  wire [6:0]  _slots_14_io_uop_prs1;
  wire [6:0]  _slots_14_io_uop_prs2;
  wire [6:0]  _slots_14_io_uop_prs3;
  wire [5:0]  _slots_14_io_uop_ppred;
  wire        _slots_14_io_uop_prs1_busy;
  wire        _slots_14_io_uop_prs2_busy;
  wire        _slots_14_io_uop_prs3_busy;
  wire        _slots_14_io_uop_ppred_busy;
  wire [6:0]  _slots_14_io_uop_stale_pdst;
  wire        _slots_14_io_uop_exception;
  wire [63:0] _slots_14_io_uop_exc_cause;
  wire        _slots_14_io_uop_bypassable;
  wire [4:0]  _slots_14_io_uop_mem_cmd;
  wire [1:0]  _slots_14_io_uop_mem_size;
  wire        _slots_14_io_uop_mem_signed;
  wire        _slots_14_io_uop_is_fence;
  wire        _slots_14_io_uop_is_fencei;
  wire        _slots_14_io_uop_is_amo;
  wire        _slots_14_io_uop_uses_ldq;
  wire        _slots_14_io_uop_uses_stq;
  wire        _slots_14_io_uop_is_sys_pc2epc;
  wire        _slots_14_io_uop_is_unique;
  wire        _slots_14_io_uop_flush_on_commit;
  wire        _slots_14_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_14_io_uop_ldst;
  wire [5:0]  _slots_14_io_uop_lrs1;
  wire [5:0]  _slots_14_io_uop_lrs2;
  wire [5:0]  _slots_14_io_uop_lrs3;
  wire        _slots_14_io_uop_ldst_val;
  wire [1:0]  _slots_14_io_uop_dst_rtype;
  wire [1:0]  _slots_14_io_uop_lrs1_rtype;
  wire [1:0]  _slots_14_io_uop_lrs2_rtype;
  wire        _slots_14_io_uop_frs3_en;
  wire        _slots_14_io_uop_fp_val;
  wire        _slots_14_io_uop_fp_single;
  wire        _slots_14_io_uop_xcpt_pf_if;
  wire        _slots_14_io_uop_xcpt_ae_if;
  wire        _slots_14_io_uop_xcpt_ma_if;
  wire        _slots_14_io_uop_bp_debug_if;
  wire        _slots_14_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_14_io_uop_debug_fsrc;
  wire [1:0]  _slots_14_io_uop_debug_tsrc;
  wire        _slots_13_io_valid;
  wire        _slots_13_io_will_be_valid;
  wire        _slots_13_io_request;
  wire [6:0]  _slots_13_io_out_uop_uopc;
  wire [31:0] _slots_13_io_out_uop_inst;
  wire [31:0] _slots_13_io_out_uop_debug_inst;
  wire        _slots_13_io_out_uop_is_rvc;
  wire [39:0] _slots_13_io_out_uop_debug_pc;
  wire [2:0]  _slots_13_io_out_uop_iq_type;
  wire [9:0]  _slots_13_io_out_uop_fu_code;
  wire [1:0]  _slots_13_io_out_uop_iw_state;
  wire        _slots_13_io_out_uop_iw_p1_poisoned;
  wire        _slots_13_io_out_uop_iw_p2_poisoned;
  wire        _slots_13_io_out_uop_is_br;
  wire        _slots_13_io_out_uop_is_jalr;
  wire        _slots_13_io_out_uop_is_jal;
  wire        _slots_13_io_out_uop_is_sfb;
  wire [19:0] _slots_13_io_out_uop_br_mask;
  wire [4:0]  _slots_13_io_out_uop_br_tag;
  wire [5:0]  _slots_13_io_out_uop_ftq_idx;
  wire        _slots_13_io_out_uop_edge_inst;
  wire [5:0]  _slots_13_io_out_uop_pc_lob;
  wire        _slots_13_io_out_uop_taken;
  wire [19:0] _slots_13_io_out_uop_imm_packed;
  wire [11:0] _slots_13_io_out_uop_csr_addr;
  wire [6:0]  _slots_13_io_out_uop_rob_idx;
  wire [4:0]  _slots_13_io_out_uop_ldq_idx;
  wire [4:0]  _slots_13_io_out_uop_stq_idx;
  wire [1:0]  _slots_13_io_out_uop_rxq_idx;
  wire [6:0]  _slots_13_io_out_uop_pdst;
  wire [6:0]  _slots_13_io_out_uop_prs1;
  wire [6:0]  _slots_13_io_out_uop_prs2;
  wire [6:0]  _slots_13_io_out_uop_prs3;
  wire [5:0]  _slots_13_io_out_uop_ppred;
  wire        _slots_13_io_out_uop_prs1_busy;
  wire        _slots_13_io_out_uop_prs2_busy;
  wire        _slots_13_io_out_uop_prs3_busy;
  wire        _slots_13_io_out_uop_ppred_busy;
  wire [6:0]  _slots_13_io_out_uop_stale_pdst;
  wire        _slots_13_io_out_uop_exception;
  wire [63:0] _slots_13_io_out_uop_exc_cause;
  wire        _slots_13_io_out_uop_bypassable;
  wire [4:0]  _slots_13_io_out_uop_mem_cmd;
  wire [1:0]  _slots_13_io_out_uop_mem_size;
  wire        _slots_13_io_out_uop_mem_signed;
  wire        _slots_13_io_out_uop_is_fence;
  wire        _slots_13_io_out_uop_is_fencei;
  wire        _slots_13_io_out_uop_is_amo;
  wire        _slots_13_io_out_uop_uses_ldq;
  wire        _slots_13_io_out_uop_uses_stq;
  wire        _slots_13_io_out_uop_is_sys_pc2epc;
  wire        _slots_13_io_out_uop_is_unique;
  wire        _slots_13_io_out_uop_flush_on_commit;
  wire        _slots_13_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_13_io_out_uop_ldst;
  wire [5:0]  _slots_13_io_out_uop_lrs1;
  wire [5:0]  _slots_13_io_out_uop_lrs2;
  wire [5:0]  _slots_13_io_out_uop_lrs3;
  wire        _slots_13_io_out_uop_ldst_val;
  wire [1:0]  _slots_13_io_out_uop_dst_rtype;
  wire [1:0]  _slots_13_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_13_io_out_uop_lrs2_rtype;
  wire        _slots_13_io_out_uop_frs3_en;
  wire        _slots_13_io_out_uop_fp_val;
  wire        _slots_13_io_out_uop_fp_single;
  wire        _slots_13_io_out_uop_xcpt_pf_if;
  wire        _slots_13_io_out_uop_xcpt_ae_if;
  wire        _slots_13_io_out_uop_xcpt_ma_if;
  wire        _slots_13_io_out_uop_bp_debug_if;
  wire        _slots_13_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_13_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_13_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_13_io_uop_uopc;
  wire [31:0] _slots_13_io_uop_inst;
  wire [31:0] _slots_13_io_uop_debug_inst;
  wire        _slots_13_io_uop_is_rvc;
  wire [39:0] _slots_13_io_uop_debug_pc;
  wire [2:0]  _slots_13_io_uop_iq_type;
  wire [9:0]  _slots_13_io_uop_fu_code;
  wire [1:0]  _slots_13_io_uop_iw_state;
  wire        _slots_13_io_uop_iw_p1_poisoned;
  wire        _slots_13_io_uop_iw_p2_poisoned;
  wire        _slots_13_io_uop_is_br;
  wire        _slots_13_io_uop_is_jalr;
  wire        _slots_13_io_uop_is_jal;
  wire        _slots_13_io_uop_is_sfb;
  wire [19:0] _slots_13_io_uop_br_mask;
  wire [4:0]  _slots_13_io_uop_br_tag;
  wire [5:0]  _slots_13_io_uop_ftq_idx;
  wire        _slots_13_io_uop_edge_inst;
  wire [5:0]  _slots_13_io_uop_pc_lob;
  wire        _slots_13_io_uop_taken;
  wire [19:0] _slots_13_io_uop_imm_packed;
  wire [11:0] _slots_13_io_uop_csr_addr;
  wire [6:0]  _slots_13_io_uop_rob_idx;
  wire [4:0]  _slots_13_io_uop_ldq_idx;
  wire [4:0]  _slots_13_io_uop_stq_idx;
  wire [1:0]  _slots_13_io_uop_rxq_idx;
  wire [6:0]  _slots_13_io_uop_pdst;
  wire [6:0]  _slots_13_io_uop_prs1;
  wire [6:0]  _slots_13_io_uop_prs2;
  wire [6:0]  _slots_13_io_uop_prs3;
  wire [5:0]  _slots_13_io_uop_ppred;
  wire        _slots_13_io_uop_prs1_busy;
  wire        _slots_13_io_uop_prs2_busy;
  wire        _slots_13_io_uop_prs3_busy;
  wire        _slots_13_io_uop_ppred_busy;
  wire [6:0]  _slots_13_io_uop_stale_pdst;
  wire        _slots_13_io_uop_exception;
  wire [63:0] _slots_13_io_uop_exc_cause;
  wire        _slots_13_io_uop_bypassable;
  wire [4:0]  _slots_13_io_uop_mem_cmd;
  wire [1:0]  _slots_13_io_uop_mem_size;
  wire        _slots_13_io_uop_mem_signed;
  wire        _slots_13_io_uop_is_fence;
  wire        _slots_13_io_uop_is_fencei;
  wire        _slots_13_io_uop_is_amo;
  wire        _slots_13_io_uop_uses_ldq;
  wire        _slots_13_io_uop_uses_stq;
  wire        _slots_13_io_uop_is_sys_pc2epc;
  wire        _slots_13_io_uop_is_unique;
  wire        _slots_13_io_uop_flush_on_commit;
  wire        _slots_13_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_13_io_uop_ldst;
  wire [5:0]  _slots_13_io_uop_lrs1;
  wire [5:0]  _slots_13_io_uop_lrs2;
  wire [5:0]  _slots_13_io_uop_lrs3;
  wire        _slots_13_io_uop_ldst_val;
  wire [1:0]  _slots_13_io_uop_dst_rtype;
  wire [1:0]  _slots_13_io_uop_lrs1_rtype;
  wire [1:0]  _slots_13_io_uop_lrs2_rtype;
  wire        _slots_13_io_uop_frs3_en;
  wire        _slots_13_io_uop_fp_val;
  wire        _slots_13_io_uop_fp_single;
  wire        _slots_13_io_uop_xcpt_pf_if;
  wire        _slots_13_io_uop_xcpt_ae_if;
  wire        _slots_13_io_uop_xcpt_ma_if;
  wire        _slots_13_io_uop_bp_debug_if;
  wire        _slots_13_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_13_io_uop_debug_fsrc;
  wire [1:0]  _slots_13_io_uop_debug_tsrc;
  wire        _slots_12_io_valid;
  wire        _slots_12_io_will_be_valid;
  wire        _slots_12_io_request;
  wire [6:0]  _slots_12_io_out_uop_uopc;
  wire [31:0] _slots_12_io_out_uop_inst;
  wire [31:0] _slots_12_io_out_uop_debug_inst;
  wire        _slots_12_io_out_uop_is_rvc;
  wire [39:0] _slots_12_io_out_uop_debug_pc;
  wire [2:0]  _slots_12_io_out_uop_iq_type;
  wire [9:0]  _slots_12_io_out_uop_fu_code;
  wire [1:0]  _slots_12_io_out_uop_iw_state;
  wire        _slots_12_io_out_uop_iw_p1_poisoned;
  wire        _slots_12_io_out_uop_iw_p2_poisoned;
  wire        _slots_12_io_out_uop_is_br;
  wire        _slots_12_io_out_uop_is_jalr;
  wire        _slots_12_io_out_uop_is_jal;
  wire        _slots_12_io_out_uop_is_sfb;
  wire [19:0] _slots_12_io_out_uop_br_mask;
  wire [4:0]  _slots_12_io_out_uop_br_tag;
  wire [5:0]  _slots_12_io_out_uop_ftq_idx;
  wire        _slots_12_io_out_uop_edge_inst;
  wire [5:0]  _slots_12_io_out_uop_pc_lob;
  wire        _slots_12_io_out_uop_taken;
  wire [19:0] _slots_12_io_out_uop_imm_packed;
  wire [11:0] _slots_12_io_out_uop_csr_addr;
  wire [6:0]  _slots_12_io_out_uop_rob_idx;
  wire [4:0]  _slots_12_io_out_uop_ldq_idx;
  wire [4:0]  _slots_12_io_out_uop_stq_idx;
  wire [1:0]  _slots_12_io_out_uop_rxq_idx;
  wire [6:0]  _slots_12_io_out_uop_pdst;
  wire [6:0]  _slots_12_io_out_uop_prs1;
  wire [6:0]  _slots_12_io_out_uop_prs2;
  wire [6:0]  _slots_12_io_out_uop_prs3;
  wire [5:0]  _slots_12_io_out_uop_ppred;
  wire        _slots_12_io_out_uop_prs1_busy;
  wire        _slots_12_io_out_uop_prs2_busy;
  wire        _slots_12_io_out_uop_prs3_busy;
  wire        _slots_12_io_out_uop_ppred_busy;
  wire [6:0]  _slots_12_io_out_uop_stale_pdst;
  wire        _slots_12_io_out_uop_exception;
  wire [63:0] _slots_12_io_out_uop_exc_cause;
  wire        _slots_12_io_out_uop_bypassable;
  wire [4:0]  _slots_12_io_out_uop_mem_cmd;
  wire [1:0]  _slots_12_io_out_uop_mem_size;
  wire        _slots_12_io_out_uop_mem_signed;
  wire        _slots_12_io_out_uop_is_fence;
  wire        _slots_12_io_out_uop_is_fencei;
  wire        _slots_12_io_out_uop_is_amo;
  wire        _slots_12_io_out_uop_uses_ldq;
  wire        _slots_12_io_out_uop_uses_stq;
  wire        _slots_12_io_out_uop_is_sys_pc2epc;
  wire        _slots_12_io_out_uop_is_unique;
  wire        _slots_12_io_out_uop_flush_on_commit;
  wire        _slots_12_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_12_io_out_uop_ldst;
  wire [5:0]  _slots_12_io_out_uop_lrs1;
  wire [5:0]  _slots_12_io_out_uop_lrs2;
  wire [5:0]  _slots_12_io_out_uop_lrs3;
  wire        _slots_12_io_out_uop_ldst_val;
  wire [1:0]  _slots_12_io_out_uop_dst_rtype;
  wire [1:0]  _slots_12_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_12_io_out_uop_lrs2_rtype;
  wire        _slots_12_io_out_uop_frs3_en;
  wire        _slots_12_io_out_uop_fp_val;
  wire        _slots_12_io_out_uop_fp_single;
  wire        _slots_12_io_out_uop_xcpt_pf_if;
  wire        _slots_12_io_out_uop_xcpt_ae_if;
  wire        _slots_12_io_out_uop_xcpt_ma_if;
  wire        _slots_12_io_out_uop_bp_debug_if;
  wire        _slots_12_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_12_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_12_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_12_io_uop_uopc;
  wire [31:0] _slots_12_io_uop_inst;
  wire [31:0] _slots_12_io_uop_debug_inst;
  wire        _slots_12_io_uop_is_rvc;
  wire [39:0] _slots_12_io_uop_debug_pc;
  wire [2:0]  _slots_12_io_uop_iq_type;
  wire [9:0]  _slots_12_io_uop_fu_code;
  wire [1:0]  _slots_12_io_uop_iw_state;
  wire        _slots_12_io_uop_iw_p1_poisoned;
  wire        _slots_12_io_uop_iw_p2_poisoned;
  wire        _slots_12_io_uop_is_br;
  wire        _slots_12_io_uop_is_jalr;
  wire        _slots_12_io_uop_is_jal;
  wire        _slots_12_io_uop_is_sfb;
  wire [19:0] _slots_12_io_uop_br_mask;
  wire [4:0]  _slots_12_io_uop_br_tag;
  wire [5:0]  _slots_12_io_uop_ftq_idx;
  wire        _slots_12_io_uop_edge_inst;
  wire [5:0]  _slots_12_io_uop_pc_lob;
  wire        _slots_12_io_uop_taken;
  wire [19:0] _slots_12_io_uop_imm_packed;
  wire [11:0] _slots_12_io_uop_csr_addr;
  wire [6:0]  _slots_12_io_uop_rob_idx;
  wire [4:0]  _slots_12_io_uop_ldq_idx;
  wire [4:0]  _slots_12_io_uop_stq_idx;
  wire [1:0]  _slots_12_io_uop_rxq_idx;
  wire [6:0]  _slots_12_io_uop_pdst;
  wire [6:0]  _slots_12_io_uop_prs1;
  wire [6:0]  _slots_12_io_uop_prs2;
  wire [6:0]  _slots_12_io_uop_prs3;
  wire [5:0]  _slots_12_io_uop_ppred;
  wire        _slots_12_io_uop_prs1_busy;
  wire        _slots_12_io_uop_prs2_busy;
  wire        _slots_12_io_uop_prs3_busy;
  wire        _slots_12_io_uop_ppred_busy;
  wire [6:0]  _slots_12_io_uop_stale_pdst;
  wire        _slots_12_io_uop_exception;
  wire [63:0] _slots_12_io_uop_exc_cause;
  wire        _slots_12_io_uop_bypassable;
  wire [4:0]  _slots_12_io_uop_mem_cmd;
  wire [1:0]  _slots_12_io_uop_mem_size;
  wire        _slots_12_io_uop_mem_signed;
  wire        _slots_12_io_uop_is_fence;
  wire        _slots_12_io_uop_is_fencei;
  wire        _slots_12_io_uop_is_amo;
  wire        _slots_12_io_uop_uses_ldq;
  wire        _slots_12_io_uop_uses_stq;
  wire        _slots_12_io_uop_is_sys_pc2epc;
  wire        _slots_12_io_uop_is_unique;
  wire        _slots_12_io_uop_flush_on_commit;
  wire        _slots_12_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_12_io_uop_ldst;
  wire [5:0]  _slots_12_io_uop_lrs1;
  wire [5:0]  _slots_12_io_uop_lrs2;
  wire [5:0]  _slots_12_io_uop_lrs3;
  wire        _slots_12_io_uop_ldst_val;
  wire [1:0]  _slots_12_io_uop_dst_rtype;
  wire [1:0]  _slots_12_io_uop_lrs1_rtype;
  wire [1:0]  _slots_12_io_uop_lrs2_rtype;
  wire        _slots_12_io_uop_frs3_en;
  wire        _slots_12_io_uop_fp_val;
  wire        _slots_12_io_uop_fp_single;
  wire        _slots_12_io_uop_xcpt_pf_if;
  wire        _slots_12_io_uop_xcpt_ae_if;
  wire        _slots_12_io_uop_xcpt_ma_if;
  wire        _slots_12_io_uop_bp_debug_if;
  wire        _slots_12_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_12_io_uop_debug_fsrc;
  wire [1:0]  _slots_12_io_uop_debug_tsrc;
  wire        _slots_11_io_valid;
  wire        _slots_11_io_will_be_valid;
  wire        _slots_11_io_request;
  wire [6:0]  _slots_11_io_out_uop_uopc;
  wire [31:0] _slots_11_io_out_uop_inst;
  wire [31:0] _slots_11_io_out_uop_debug_inst;
  wire        _slots_11_io_out_uop_is_rvc;
  wire [39:0] _slots_11_io_out_uop_debug_pc;
  wire [2:0]  _slots_11_io_out_uop_iq_type;
  wire [9:0]  _slots_11_io_out_uop_fu_code;
  wire [1:0]  _slots_11_io_out_uop_iw_state;
  wire        _slots_11_io_out_uop_iw_p1_poisoned;
  wire        _slots_11_io_out_uop_iw_p2_poisoned;
  wire        _slots_11_io_out_uop_is_br;
  wire        _slots_11_io_out_uop_is_jalr;
  wire        _slots_11_io_out_uop_is_jal;
  wire        _slots_11_io_out_uop_is_sfb;
  wire [19:0] _slots_11_io_out_uop_br_mask;
  wire [4:0]  _slots_11_io_out_uop_br_tag;
  wire [5:0]  _slots_11_io_out_uop_ftq_idx;
  wire        _slots_11_io_out_uop_edge_inst;
  wire [5:0]  _slots_11_io_out_uop_pc_lob;
  wire        _slots_11_io_out_uop_taken;
  wire [19:0] _slots_11_io_out_uop_imm_packed;
  wire [11:0] _slots_11_io_out_uop_csr_addr;
  wire [6:0]  _slots_11_io_out_uop_rob_idx;
  wire [4:0]  _slots_11_io_out_uop_ldq_idx;
  wire [4:0]  _slots_11_io_out_uop_stq_idx;
  wire [1:0]  _slots_11_io_out_uop_rxq_idx;
  wire [6:0]  _slots_11_io_out_uop_pdst;
  wire [6:0]  _slots_11_io_out_uop_prs1;
  wire [6:0]  _slots_11_io_out_uop_prs2;
  wire [6:0]  _slots_11_io_out_uop_prs3;
  wire [5:0]  _slots_11_io_out_uop_ppred;
  wire        _slots_11_io_out_uop_prs1_busy;
  wire        _slots_11_io_out_uop_prs2_busy;
  wire        _slots_11_io_out_uop_prs3_busy;
  wire        _slots_11_io_out_uop_ppred_busy;
  wire [6:0]  _slots_11_io_out_uop_stale_pdst;
  wire        _slots_11_io_out_uop_exception;
  wire [63:0] _slots_11_io_out_uop_exc_cause;
  wire        _slots_11_io_out_uop_bypassable;
  wire [4:0]  _slots_11_io_out_uop_mem_cmd;
  wire [1:0]  _slots_11_io_out_uop_mem_size;
  wire        _slots_11_io_out_uop_mem_signed;
  wire        _slots_11_io_out_uop_is_fence;
  wire        _slots_11_io_out_uop_is_fencei;
  wire        _slots_11_io_out_uop_is_amo;
  wire        _slots_11_io_out_uop_uses_ldq;
  wire        _slots_11_io_out_uop_uses_stq;
  wire        _slots_11_io_out_uop_is_sys_pc2epc;
  wire        _slots_11_io_out_uop_is_unique;
  wire        _slots_11_io_out_uop_flush_on_commit;
  wire        _slots_11_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_11_io_out_uop_ldst;
  wire [5:0]  _slots_11_io_out_uop_lrs1;
  wire [5:0]  _slots_11_io_out_uop_lrs2;
  wire [5:0]  _slots_11_io_out_uop_lrs3;
  wire        _slots_11_io_out_uop_ldst_val;
  wire [1:0]  _slots_11_io_out_uop_dst_rtype;
  wire [1:0]  _slots_11_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_11_io_out_uop_lrs2_rtype;
  wire        _slots_11_io_out_uop_frs3_en;
  wire        _slots_11_io_out_uop_fp_val;
  wire        _slots_11_io_out_uop_fp_single;
  wire        _slots_11_io_out_uop_xcpt_pf_if;
  wire        _slots_11_io_out_uop_xcpt_ae_if;
  wire        _slots_11_io_out_uop_xcpt_ma_if;
  wire        _slots_11_io_out_uop_bp_debug_if;
  wire        _slots_11_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_11_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_11_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_11_io_uop_uopc;
  wire [31:0] _slots_11_io_uop_inst;
  wire [31:0] _slots_11_io_uop_debug_inst;
  wire        _slots_11_io_uop_is_rvc;
  wire [39:0] _slots_11_io_uop_debug_pc;
  wire [2:0]  _slots_11_io_uop_iq_type;
  wire [9:0]  _slots_11_io_uop_fu_code;
  wire [1:0]  _slots_11_io_uop_iw_state;
  wire        _slots_11_io_uop_iw_p1_poisoned;
  wire        _slots_11_io_uop_iw_p2_poisoned;
  wire        _slots_11_io_uop_is_br;
  wire        _slots_11_io_uop_is_jalr;
  wire        _slots_11_io_uop_is_jal;
  wire        _slots_11_io_uop_is_sfb;
  wire [19:0] _slots_11_io_uop_br_mask;
  wire [4:0]  _slots_11_io_uop_br_tag;
  wire [5:0]  _slots_11_io_uop_ftq_idx;
  wire        _slots_11_io_uop_edge_inst;
  wire [5:0]  _slots_11_io_uop_pc_lob;
  wire        _slots_11_io_uop_taken;
  wire [19:0] _slots_11_io_uop_imm_packed;
  wire [11:0] _slots_11_io_uop_csr_addr;
  wire [6:0]  _slots_11_io_uop_rob_idx;
  wire [4:0]  _slots_11_io_uop_ldq_idx;
  wire [4:0]  _slots_11_io_uop_stq_idx;
  wire [1:0]  _slots_11_io_uop_rxq_idx;
  wire [6:0]  _slots_11_io_uop_pdst;
  wire [6:0]  _slots_11_io_uop_prs1;
  wire [6:0]  _slots_11_io_uop_prs2;
  wire [6:0]  _slots_11_io_uop_prs3;
  wire [5:0]  _slots_11_io_uop_ppred;
  wire        _slots_11_io_uop_prs1_busy;
  wire        _slots_11_io_uop_prs2_busy;
  wire        _slots_11_io_uop_prs3_busy;
  wire        _slots_11_io_uop_ppred_busy;
  wire [6:0]  _slots_11_io_uop_stale_pdst;
  wire        _slots_11_io_uop_exception;
  wire [63:0] _slots_11_io_uop_exc_cause;
  wire        _slots_11_io_uop_bypassable;
  wire [4:0]  _slots_11_io_uop_mem_cmd;
  wire [1:0]  _slots_11_io_uop_mem_size;
  wire        _slots_11_io_uop_mem_signed;
  wire        _slots_11_io_uop_is_fence;
  wire        _slots_11_io_uop_is_fencei;
  wire        _slots_11_io_uop_is_amo;
  wire        _slots_11_io_uop_uses_ldq;
  wire        _slots_11_io_uop_uses_stq;
  wire        _slots_11_io_uop_is_sys_pc2epc;
  wire        _slots_11_io_uop_is_unique;
  wire        _slots_11_io_uop_flush_on_commit;
  wire        _slots_11_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_11_io_uop_ldst;
  wire [5:0]  _slots_11_io_uop_lrs1;
  wire [5:0]  _slots_11_io_uop_lrs2;
  wire [5:0]  _slots_11_io_uop_lrs3;
  wire        _slots_11_io_uop_ldst_val;
  wire [1:0]  _slots_11_io_uop_dst_rtype;
  wire [1:0]  _slots_11_io_uop_lrs1_rtype;
  wire [1:0]  _slots_11_io_uop_lrs2_rtype;
  wire        _slots_11_io_uop_frs3_en;
  wire        _slots_11_io_uop_fp_val;
  wire        _slots_11_io_uop_fp_single;
  wire        _slots_11_io_uop_xcpt_pf_if;
  wire        _slots_11_io_uop_xcpt_ae_if;
  wire        _slots_11_io_uop_xcpt_ma_if;
  wire        _slots_11_io_uop_bp_debug_if;
  wire        _slots_11_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_11_io_uop_debug_fsrc;
  wire [1:0]  _slots_11_io_uop_debug_tsrc;
  wire        _slots_10_io_valid;
  wire        _slots_10_io_will_be_valid;
  wire        _slots_10_io_request;
  wire [6:0]  _slots_10_io_out_uop_uopc;
  wire [31:0] _slots_10_io_out_uop_inst;
  wire [31:0] _slots_10_io_out_uop_debug_inst;
  wire        _slots_10_io_out_uop_is_rvc;
  wire [39:0] _slots_10_io_out_uop_debug_pc;
  wire [2:0]  _slots_10_io_out_uop_iq_type;
  wire [9:0]  _slots_10_io_out_uop_fu_code;
  wire [1:0]  _slots_10_io_out_uop_iw_state;
  wire        _slots_10_io_out_uop_iw_p1_poisoned;
  wire        _slots_10_io_out_uop_iw_p2_poisoned;
  wire        _slots_10_io_out_uop_is_br;
  wire        _slots_10_io_out_uop_is_jalr;
  wire        _slots_10_io_out_uop_is_jal;
  wire        _slots_10_io_out_uop_is_sfb;
  wire [19:0] _slots_10_io_out_uop_br_mask;
  wire [4:0]  _slots_10_io_out_uop_br_tag;
  wire [5:0]  _slots_10_io_out_uop_ftq_idx;
  wire        _slots_10_io_out_uop_edge_inst;
  wire [5:0]  _slots_10_io_out_uop_pc_lob;
  wire        _slots_10_io_out_uop_taken;
  wire [19:0] _slots_10_io_out_uop_imm_packed;
  wire [11:0] _slots_10_io_out_uop_csr_addr;
  wire [6:0]  _slots_10_io_out_uop_rob_idx;
  wire [4:0]  _slots_10_io_out_uop_ldq_idx;
  wire [4:0]  _slots_10_io_out_uop_stq_idx;
  wire [1:0]  _slots_10_io_out_uop_rxq_idx;
  wire [6:0]  _slots_10_io_out_uop_pdst;
  wire [6:0]  _slots_10_io_out_uop_prs1;
  wire [6:0]  _slots_10_io_out_uop_prs2;
  wire [6:0]  _slots_10_io_out_uop_prs3;
  wire [5:0]  _slots_10_io_out_uop_ppred;
  wire        _slots_10_io_out_uop_prs1_busy;
  wire        _slots_10_io_out_uop_prs2_busy;
  wire        _slots_10_io_out_uop_prs3_busy;
  wire        _slots_10_io_out_uop_ppred_busy;
  wire [6:0]  _slots_10_io_out_uop_stale_pdst;
  wire        _slots_10_io_out_uop_exception;
  wire [63:0] _slots_10_io_out_uop_exc_cause;
  wire        _slots_10_io_out_uop_bypassable;
  wire [4:0]  _slots_10_io_out_uop_mem_cmd;
  wire [1:0]  _slots_10_io_out_uop_mem_size;
  wire        _slots_10_io_out_uop_mem_signed;
  wire        _slots_10_io_out_uop_is_fence;
  wire        _slots_10_io_out_uop_is_fencei;
  wire        _slots_10_io_out_uop_is_amo;
  wire        _slots_10_io_out_uop_uses_ldq;
  wire        _slots_10_io_out_uop_uses_stq;
  wire        _slots_10_io_out_uop_is_sys_pc2epc;
  wire        _slots_10_io_out_uop_is_unique;
  wire        _slots_10_io_out_uop_flush_on_commit;
  wire        _slots_10_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_10_io_out_uop_ldst;
  wire [5:0]  _slots_10_io_out_uop_lrs1;
  wire [5:0]  _slots_10_io_out_uop_lrs2;
  wire [5:0]  _slots_10_io_out_uop_lrs3;
  wire        _slots_10_io_out_uop_ldst_val;
  wire [1:0]  _slots_10_io_out_uop_dst_rtype;
  wire [1:0]  _slots_10_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_10_io_out_uop_lrs2_rtype;
  wire        _slots_10_io_out_uop_frs3_en;
  wire        _slots_10_io_out_uop_fp_val;
  wire        _slots_10_io_out_uop_fp_single;
  wire        _slots_10_io_out_uop_xcpt_pf_if;
  wire        _slots_10_io_out_uop_xcpt_ae_if;
  wire        _slots_10_io_out_uop_xcpt_ma_if;
  wire        _slots_10_io_out_uop_bp_debug_if;
  wire        _slots_10_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_10_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_10_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_10_io_uop_uopc;
  wire [31:0] _slots_10_io_uop_inst;
  wire [31:0] _slots_10_io_uop_debug_inst;
  wire        _slots_10_io_uop_is_rvc;
  wire [39:0] _slots_10_io_uop_debug_pc;
  wire [2:0]  _slots_10_io_uop_iq_type;
  wire [9:0]  _slots_10_io_uop_fu_code;
  wire [1:0]  _slots_10_io_uop_iw_state;
  wire        _slots_10_io_uop_iw_p1_poisoned;
  wire        _slots_10_io_uop_iw_p2_poisoned;
  wire        _slots_10_io_uop_is_br;
  wire        _slots_10_io_uop_is_jalr;
  wire        _slots_10_io_uop_is_jal;
  wire        _slots_10_io_uop_is_sfb;
  wire [19:0] _slots_10_io_uop_br_mask;
  wire [4:0]  _slots_10_io_uop_br_tag;
  wire [5:0]  _slots_10_io_uop_ftq_idx;
  wire        _slots_10_io_uop_edge_inst;
  wire [5:0]  _slots_10_io_uop_pc_lob;
  wire        _slots_10_io_uop_taken;
  wire [19:0] _slots_10_io_uop_imm_packed;
  wire [11:0] _slots_10_io_uop_csr_addr;
  wire [6:0]  _slots_10_io_uop_rob_idx;
  wire [4:0]  _slots_10_io_uop_ldq_idx;
  wire [4:0]  _slots_10_io_uop_stq_idx;
  wire [1:0]  _slots_10_io_uop_rxq_idx;
  wire [6:0]  _slots_10_io_uop_pdst;
  wire [6:0]  _slots_10_io_uop_prs1;
  wire [6:0]  _slots_10_io_uop_prs2;
  wire [6:0]  _slots_10_io_uop_prs3;
  wire [5:0]  _slots_10_io_uop_ppred;
  wire        _slots_10_io_uop_prs1_busy;
  wire        _slots_10_io_uop_prs2_busy;
  wire        _slots_10_io_uop_prs3_busy;
  wire        _slots_10_io_uop_ppred_busy;
  wire [6:0]  _slots_10_io_uop_stale_pdst;
  wire        _slots_10_io_uop_exception;
  wire [63:0] _slots_10_io_uop_exc_cause;
  wire        _slots_10_io_uop_bypassable;
  wire [4:0]  _slots_10_io_uop_mem_cmd;
  wire [1:0]  _slots_10_io_uop_mem_size;
  wire        _slots_10_io_uop_mem_signed;
  wire        _slots_10_io_uop_is_fence;
  wire        _slots_10_io_uop_is_fencei;
  wire        _slots_10_io_uop_is_amo;
  wire        _slots_10_io_uop_uses_ldq;
  wire        _slots_10_io_uop_uses_stq;
  wire        _slots_10_io_uop_is_sys_pc2epc;
  wire        _slots_10_io_uop_is_unique;
  wire        _slots_10_io_uop_flush_on_commit;
  wire        _slots_10_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_10_io_uop_ldst;
  wire [5:0]  _slots_10_io_uop_lrs1;
  wire [5:0]  _slots_10_io_uop_lrs2;
  wire [5:0]  _slots_10_io_uop_lrs3;
  wire        _slots_10_io_uop_ldst_val;
  wire [1:0]  _slots_10_io_uop_dst_rtype;
  wire [1:0]  _slots_10_io_uop_lrs1_rtype;
  wire [1:0]  _slots_10_io_uop_lrs2_rtype;
  wire        _slots_10_io_uop_frs3_en;
  wire        _slots_10_io_uop_fp_val;
  wire        _slots_10_io_uop_fp_single;
  wire        _slots_10_io_uop_xcpt_pf_if;
  wire        _slots_10_io_uop_xcpt_ae_if;
  wire        _slots_10_io_uop_xcpt_ma_if;
  wire        _slots_10_io_uop_bp_debug_if;
  wire        _slots_10_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_10_io_uop_debug_fsrc;
  wire [1:0]  _slots_10_io_uop_debug_tsrc;
  wire        _slots_9_io_valid;
  wire        _slots_9_io_will_be_valid;
  wire        _slots_9_io_request;
  wire [6:0]  _slots_9_io_out_uop_uopc;
  wire [31:0] _slots_9_io_out_uop_inst;
  wire [31:0] _slots_9_io_out_uop_debug_inst;
  wire        _slots_9_io_out_uop_is_rvc;
  wire [39:0] _slots_9_io_out_uop_debug_pc;
  wire [2:0]  _slots_9_io_out_uop_iq_type;
  wire [9:0]  _slots_9_io_out_uop_fu_code;
  wire [1:0]  _slots_9_io_out_uop_iw_state;
  wire        _slots_9_io_out_uop_iw_p1_poisoned;
  wire        _slots_9_io_out_uop_iw_p2_poisoned;
  wire        _slots_9_io_out_uop_is_br;
  wire        _slots_9_io_out_uop_is_jalr;
  wire        _slots_9_io_out_uop_is_jal;
  wire        _slots_9_io_out_uop_is_sfb;
  wire [19:0] _slots_9_io_out_uop_br_mask;
  wire [4:0]  _slots_9_io_out_uop_br_tag;
  wire [5:0]  _slots_9_io_out_uop_ftq_idx;
  wire        _slots_9_io_out_uop_edge_inst;
  wire [5:0]  _slots_9_io_out_uop_pc_lob;
  wire        _slots_9_io_out_uop_taken;
  wire [19:0] _slots_9_io_out_uop_imm_packed;
  wire [11:0] _slots_9_io_out_uop_csr_addr;
  wire [6:0]  _slots_9_io_out_uop_rob_idx;
  wire [4:0]  _slots_9_io_out_uop_ldq_idx;
  wire [4:0]  _slots_9_io_out_uop_stq_idx;
  wire [1:0]  _slots_9_io_out_uop_rxq_idx;
  wire [6:0]  _slots_9_io_out_uop_pdst;
  wire [6:0]  _slots_9_io_out_uop_prs1;
  wire [6:0]  _slots_9_io_out_uop_prs2;
  wire [6:0]  _slots_9_io_out_uop_prs3;
  wire [5:0]  _slots_9_io_out_uop_ppred;
  wire        _slots_9_io_out_uop_prs1_busy;
  wire        _slots_9_io_out_uop_prs2_busy;
  wire        _slots_9_io_out_uop_prs3_busy;
  wire        _slots_9_io_out_uop_ppred_busy;
  wire [6:0]  _slots_9_io_out_uop_stale_pdst;
  wire        _slots_9_io_out_uop_exception;
  wire [63:0] _slots_9_io_out_uop_exc_cause;
  wire        _slots_9_io_out_uop_bypassable;
  wire [4:0]  _slots_9_io_out_uop_mem_cmd;
  wire [1:0]  _slots_9_io_out_uop_mem_size;
  wire        _slots_9_io_out_uop_mem_signed;
  wire        _slots_9_io_out_uop_is_fence;
  wire        _slots_9_io_out_uop_is_fencei;
  wire        _slots_9_io_out_uop_is_amo;
  wire        _slots_9_io_out_uop_uses_ldq;
  wire        _slots_9_io_out_uop_uses_stq;
  wire        _slots_9_io_out_uop_is_sys_pc2epc;
  wire        _slots_9_io_out_uop_is_unique;
  wire        _slots_9_io_out_uop_flush_on_commit;
  wire        _slots_9_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_9_io_out_uop_ldst;
  wire [5:0]  _slots_9_io_out_uop_lrs1;
  wire [5:0]  _slots_9_io_out_uop_lrs2;
  wire [5:0]  _slots_9_io_out_uop_lrs3;
  wire        _slots_9_io_out_uop_ldst_val;
  wire [1:0]  _slots_9_io_out_uop_dst_rtype;
  wire [1:0]  _slots_9_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_9_io_out_uop_lrs2_rtype;
  wire        _slots_9_io_out_uop_frs3_en;
  wire        _slots_9_io_out_uop_fp_val;
  wire        _slots_9_io_out_uop_fp_single;
  wire        _slots_9_io_out_uop_xcpt_pf_if;
  wire        _slots_9_io_out_uop_xcpt_ae_if;
  wire        _slots_9_io_out_uop_xcpt_ma_if;
  wire        _slots_9_io_out_uop_bp_debug_if;
  wire        _slots_9_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_9_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_9_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_9_io_uop_uopc;
  wire [31:0] _slots_9_io_uop_inst;
  wire [31:0] _slots_9_io_uop_debug_inst;
  wire        _slots_9_io_uop_is_rvc;
  wire [39:0] _slots_9_io_uop_debug_pc;
  wire [2:0]  _slots_9_io_uop_iq_type;
  wire [9:0]  _slots_9_io_uop_fu_code;
  wire [1:0]  _slots_9_io_uop_iw_state;
  wire        _slots_9_io_uop_iw_p1_poisoned;
  wire        _slots_9_io_uop_iw_p2_poisoned;
  wire        _slots_9_io_uop_is_br;
  wire        _slots_9_io_uop_is_jalr;
  wire        _slots_9_io_uop_is_jal;
  wire        _slots_9_io_uop_is_sfb;
  wire [19:0] _slots_9_io_uop_br_mask;
  wire [4:0]  _slots_9_io_uop_br_tag;
  wire [5:0]  _slots_9_io_uop_ftq_idx;
  wire        _slots_9_io_uop_edge_inst;
  wire [5:0]  _slots_9_io_uop_pc_lob;
  wire        _slots_9_io_uop_taken;
  wire [19:0] _slots_9_io_uop_imm_packed;
  wire [11:0] _slots_9_io_uop_csr_addr;
  wire [6:0]  _slots_9_io_uop_rob_idx;
  wire [4:0]  _slots_9_io_uop_ldq_idx;
  wire [4:0]  _slots_9_io_uop_stq_idx;
  wire [1:0]  _slots_9_io_uop_rxq_idx;
  wire [6:0]  _slots_9_io_uop_pdst;
  wire [6:0]  _slots_9_io_uop_prs1;
  wire [6:0]  _slots_9_io_uop_prs2;
  wire [6:0]  _slots_9_io_uop_prs3;
  wire [5:0]  _slots_9_io_uop_ppred;
  wire        _slots_9_io_uop_prs1_busy;
  wire        _slots_9_io_uop_prs2_busy;
  wire        _slots_9_io_uop_prs3_busy;
  wire        _slots_9_io_uop_ppred_busy;
  wire [6:0]  _slots_9_io_uop_stale_pdst;
  wire        _slots_9_io_uop_exception;
  wire [63:0] _slots_9_io_uop_exc_cause;
  wire        _slots_9_io_uop_bypassable;
  wire [4:0]  _slots_9_io_uop_mem_cmd;
  wire [1:0]  _slots_9_io_uop_mem_size;
  wire        _slots_9_io_uop_mem_signed;
  wire        _slots_9_io_uop_is_fence;
  wire        _slots_9_io_uop_is_fencei;
  wire        _slots_9_io_uop_is_amo;
  wire        _slots_9_io_uop_uses_ldq;
  wire        _slots_9_io_uop_uses_stq;
  wire        _slots_9_io_uop_is_sys_pc2epc;
  wire        _slots_9_io_uop_is_unique;
  wire        _slots_9_io_uop_flush_on_commit;
  wire        _slots_9_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_9_io_uop_ldst;
  wire [5:0]  _slots_9_io_uop_lrs1;
  wire [5:0]  _slots_9_io_uop_lrs2;
  wire [5:0]  _slots_9_io_uop_lrs3;
  wire        _slots_9_io_uop_ldst_val;
  wire [1:0]  _slots_9_io_uop_dst_rtype;
  wire [1:0]  _slots_9_io_uop_lrs1_rtype;
  wire [1:0]  _slots_9_io_uop_lrs2_rtype;
  wire        _slots_9_io_uop_frs3_en;
  wire        _slots_9_io_uop_fp_val;
  wire        _slots_9_io_uop_fp_single;
  wire        _slots_9_io_uop_xcpt_pf_if;
  wire        _slots_9_io_uop_xcpt_ae_if;
  wire        _slots_9_io_uop_xcpt_ma_if;
  wire        _slots_9_io_uop_bp_debug_if;
  wire        _slots_9_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_9_io_uop_debug_fsrc;
  wire [1:0]  _slots_9_io_uop_debug_tsrc;
  wire        _slots_8_io_valid;
  wire        _slots_8_io_will_be_valid;
  wire        _slots_8_io_request;
  wire [6:0]  _slots_8_io_out_uop_uopc;
  wire [31:0] _slots_8_io_out_uop_inst;
  wire [31:0] _slots_8_io_out_uop_debug_inst;
  wire        _slots_8_io_out_uop_is_rvc;
  wire [39:0] _slots_8_io_out_uop_debug_pc;
  wire [2:0]  _slots_8_io_out_uop_iq_type;
  wire [9:0]  _slots_8_io_out_uop_fu_code;
  wire [1:0]  _slots_8_io_out_uop_iw_state;
  wire        _slots_8_io_out_uop_iw_p1_poisoned;
  wire        _slots_8_io_out_uop_iw_p2_poisoned;
  wire        _slots_8_io_out_uop_is_br;
  wire        _slots_8_io_out_uop_is_jalr;
  wire        _slots_8_io_out_uop_is_jal;
  wire        _slots_8_io_out_uop_is_sfb;
  wire [19:0] _slots_8_io_out_uop_br_mask;
  wire [4:0]  _slots_8_io_out_uop_br_tag;
  wire [5:0]  _slots_8_io_out_uop_ftq_idx;
  wire        _slots_8_io_out_uop_edge_inst;
  wire [5:0]  _slots_8_io_out_uop_pc_lob;
  wire        _slots_8_io_out_uop_taken;
  wire [19:0] _slots_8_io_out_uop_imm_packed;
  wire [11:0] _slots_8_io_out_uop_csr_addr;
  wire [6:0]  _slots_8_io_out_uop_rob_idx;
  wire [4:0]  _slots_8_io_out_uop_ldq_idx;
  wire [4:0]  _slots_8_io_out_uop_stq_idx;
  wire [1:0]  _slots_8_io_out_uop_rxq_idx;
  wire [6:0]  _slots_8_io_out_uop_pdst;
  wire [6:0]  _slots_8_io_out_uop_prs1;
  wire [6:0]  _slots_8_io_out_uop_prs2;
  wire [6:0]  _slots_8_io_out_uop_prs3;
  wire [5:0]  _slots_8_io_out_uop_ppred;
  wire        _slots_8_io_out_uop_prs1_busy;
  wire        _slots_8_io_out_uop_prs2_busy;
  wire        _slots_8_io_out_uop_prs3_busy;
  wire        _slots_8_io_out_uop_ppred_busy;
  wire [6:0]  _slots_8_io_out_uop_stale_pdst;
  wire        _slots_8_io_out_uop_exception;
  wire [63:0] _slots_8_io_out_uop_exc_cause;
  wire        _slots_8_io_out_uop_bypassable;
  wire [4:0]  _slots_8_io_out_uop_mem_cmd;
  wire [1:0]  _slots_8_io_out_uop_mem_size;
  wire        _slots_8_io_out_uop_mem_signed;
  wire        _slots_8_io_out_uop_is_fence;
  wire        _slots_8_io_out_uop_is_fencei;
  wire        _slots_8_io_out_uop_is_amo;
  wire        _slots_8_io_out_uop_uses_ldq;
  wire        _slots_8_io_out_uop_uses_stq;
  wire        _slots_8_io_out_uop_is_sys_pc2epc;
  wire        _slots_8_io_out_uop_is_unique;
  wire        _slots_8_io_out_uop_flush_on_commit;
  wire        _slots_8_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_8_io_out_uop_ldst;
  wire [5:0]  _slots_8_io_out_uop_lrs1;
  wire [5:0]  _slots_8_io_out_uop_lrs2;
  wire [5:0]  _slots_8_io_out_uop_lrs3;
  wire        _slots_8_io_out_uop_ldst_val;
  wire [1:0]  _slots_8_io_out_uop_dst_rtype;
  wire [1:0]  _slots_8_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_8_io_out_uop_lrs2_rtype;
  wire        _slots_8_io_out_uop_frs3_en;
  wire        _slots_8_io_out_uop_fp_val;
  wire        _slots_8_io_out_uop_fp_single;
  wire        _slots_8_io_out_uop_xcpt_pf_if;
  wire        _slots_8_io_out_uop_xcpt_ae_if;
  wire        _slots_8_io_out_uop_xcpt_ma_if;
  wire        _slots_8_io_out_uop_bp_debug_if;
  wire        _slots_8_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_8_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_8_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_8_io_uop_uopc;
  wire [31:0] _slots_8_io_uop_inst;
  wire [31:0] _slots_8_io_uop_debug_inst;
  wire        _slots_8_io_uop_is_rvc;
  wire [39:0] _slots_8_io_uop_debug_pc;
  wire [2:0]  _slots_8_io_uop_iq_type;
  wire [9:0]  _slots_8_io_uop_fu_code;
  wire [1:0]  _slots_8_io_uop_iw_state;
  wire        _slots_8_io_uop_iw_p1_poisoned;
  wire        _slots_8_io_uop_iw_p2_poisoned;
  wire        _slots_8_io_uop_is_br;
  wire        _slots_8_io_uop_is_jalr;
  wire        _slots_8_io_uop_is_jal;
  wire        _slots_8_io_uop_is_sfb;
  wire [19:0] _slots_8_io_uop_br_mask;
  wire [4:0]  _slots_8_io_uop_br_tag;
  wire [5:0]  _slots_8_io_uop_ftq_idx;
  wire        _slots_8_io_uop_edge_inst;
  wire [5:0]  _slots_8_io_uop_pc_lob;
  wire        _slots_8_io_uop_taken;
  wire [19:0] _slots_8_io_uop_imm_packed;
  wire [11:0] _slots_8_io_uop_csr_addr;
  wire [6:0]  _slots_8_io_uop_rob_idx;
  wire [4:0]  _slots_8_io_uop_ldq_idx;
  wire [4:0]  _slots_8_io_uop_stq_idx;
  wire [1:0]  _slots_8_io_uop_rxq_idx;
  wire [6:0]  _slots_8_io_uop_pdst;
  wire [6:0]  _slots_8_io_uop_prs1;
  wire [6:0]  _slots_8_io_uop_prs2;
  wire [6:0]  _slots_8_io_uop_prs3;
  wire [5:0]  _slots_8_io_uop_ppred;
  wire        _slots_8_io_uop_prs1_busy;
  wire        _slots_8_io_uop_prs2_busy;
  wire        _slots_8_io_uop_prs3_busy;
  wire        _slots_8_io_uop_ppred_busy;
  wire [6:0]  _slots_8_io_uop_stale_pdst;
  wire        _slots_8_io_uop_exception;
  wire [63:0] _slots_8_io_uop_exc_cause;
  wire        _slots_8_io_uop_bypassable;
  wire [4:0]  _slots_8_io_uop_mem_cmd;
  wire [1:0]  _slots_8_io_uop_mem_size;
  wire        _slots_8_io_uop_mem_signed;
  wire        _slots_8_io_uop_is_fence;
  wire        _slots_8_io_uop_is_fencei;
  wire        _slots_8_io_uop_is_amo;
  wire        _slots_8_io_uop_uses_ldq;
  wire        _slots_8_io_uop_uses_stq;
  wire        _slots_8_io_uop_is_sys_pc2epc;
  wire        _slots_8_io_uop_is_unique;
  wire        _slots_8_io_uop_flush_on_commit;
  wire        _slots_8_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_8_io_uop_ldst;
  wire [5:0]  _slots_8_io_uop_lrs1;
  wire [5:0]  _slots_8_io_uop_lrs2;
  wire [5:0]  _slots_8_io_uop_lrs3;
  wire        _slots_8_io_uop_ldst_val;
  wire [1:0]  _slots_8_io_uop_dst_rtype;
  wire [1:0]  _slots_8_io_uop_lrs1_rtype;
  wire [1:0]  _slots_8_io_uop_lrs2_rtype;
  wire        _slots_8_io_uop_frs3_en;
  wire        _slots_8_io_uop_fp_val;
  wire        _slots_8_io_uop_fp_single;
  wire        _slots_8_io_uop_xcpt_pf_if;
  wire        _slots_8_io_uop_xcpt_ae_if;
  wire        _slots_8_io_uop_xcpt_ma_if;
  wire        _slots_8_io_uop_bp_debug_if;
  wire        _slots_8_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_8_io_uop_debug_fsrc;
  wire [1:0]  _slots_8_io_uop_debug_tsrc;
  wire        _slots_7_io_valid;
  wire        _slots_7_io_will_be_valid;
  wire        _slots_7_io_request;
  wire [6:0]  _slots_7_io_out_uop_uopc;
  wire [31:0] _slots_7_io_out_uop_inst;
  wire [31:0] _slots_7_io_out_uop_debug_inst;
  wire        _slots_7_io_out_uop_is_rvc;
  wire [39:0] _slots_7_io_out_uop_debug_pc;
  wire [2:0]  _slots_7_io_out_uop_iq_type;
  wire [9:0]  _slots_7_io_out_uop_fu_code;
  wire [1:0]  _slots_7_io_out_uop_iw_state;
  wire        _slots_7_io_out_uop_iw_p1_poisoned;
  wire        _slots_7_io_out_uop_iw_p2_poisoned;
  wire        _slots_7_io_out_uop_is_br;
  wire        _slots_7_io_out_uop_is_jalr;
  wire        _slots_7_io_out_uop_is_jal;
  wire        _slots_7_io_out_uop_is_sfb;
  wire [19:0] _slots_7_io_out_uop_br_mask;
  wire [4:0]  _slots_7_io_out_uop_br_tag;
  wire [5:0]  _slots_7_io_out_uop_ftq_idx;
  wire        _slots_7_io_out_uop_edge_inst;
  wire [5:0]  _slots_7_io_out_uop_pc_lob;
  wire        _slots_7_io_out_uop_taken;
  wire [19:0] _slots_7_io_out_uop_imm_packed;
  wire [11:0] _slots_7_io_out_uop_csr_addr;
  wire [6:0]  _slots_7_io_out_uop_rob_idx;
  wire [4:0]  _slots_7_io_out_uop_ldq_idx;
  wire [4:0]  _slots_7_io_out_uop_stq_idx;
  wire [1:0]  _slots_7_io_out_uop_rxq_idx;
  wire [6:0]  _slots_7_io_out_uop_pdst;
  wire [6:0]  _slots_7_io_out_uop_prs1;
  wire [6:0]  _slots_7_io_out_uop_prs2;
  wire [6:0]  _slots_7_io_out_uop_prs3;
  wire [5:0]  _slots_7_io_out_uop_ppred;
  wire        _slots_7_io_out_uop_prs1_busy;
  wire        _slots_7_io_out_uop_prs2_busy;
  wire        _slots_7_io_out_uop_prs3_busy;
  wire        _slots_7_io_out_uop_ppred_busy;
  wire [6:0]  _slots_7_io_out_uop_stale_pdst;
  wire        _slots_7_io_out_uop_exception;
  wire [63:0] _slots_7_io_out_uop_exc_cause;
  wire        _slots_7_io_out_uop_bypassable;
  wire [4:0]  _slots_7_io_out_uop_mem_cmd;
  wire [1:0]  _slots_7_io_out_uop_mem_size;
  wire        _slots_7_io_out_uop_mem_signed;
  wire        _slots_7_io_out_uop_is_fence;
  wire        _slots_7_io_out_uop_is_fencei;
  wire        _slots_7_io_out_uop_is_amo;
  wire        _slots_7_io_out_uop_uses_ldq;
  wire        _slots_7_io_out_uop_uses_stq;
  wire        _slots_7_io_out_uop_is_sys_pc2epc;
  wire        _slots_7_io_out_uop_is_unique;
  wire        _slots_7_io_out_uop_flush_on_commit;
  wire        _slots_7_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_7_io_out_uop_ldst;
  wire [5:0]  _slots_7_io_out_uop_lrs1;
  wire [5:0]  _slots_7_io_out_uop_lrs2;
  wire [5:0]  _slots_7_io_out_uop_lrs3;
  wire        _slots_7_io_out_uop_ldst_val;
  wire [1:0]  _slots_7_io_out_uop_dst_rtype;
  wire [1:0]  _slots_7_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_7_io_out_uop_lrs2_rtype;
  wire        _slots_7_io_out_uop_frs3_en;
  wire        _slots_7_io_out_uop_fp_val;
  wire        _slots_7_io_out_uop_fp_single;
  wire        _slots_7_io_out_uop_xcpt_pf_if;
  wire        _slots_7_io_out_uop_xcpt_ae_if;
  wire        _slots_7_io_out_uop_xcpt_ma_if;
  wire        _slots_7_io_out_uop_bp_debug_if;
  wire        _slots_7_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_7_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_7_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_7_io_uop_uopc;
  wire [31:0] _slots_7_io_uop_inst;
  wire [31:0] _slots_7_io_uop_debug_inst;
  wire        _slots_7_io_uop_is_rvc;
  wire [39:0] _slots_7_io_uop_debug_pc;
  wire [2:0]  _slots_7_io_uop_iq_type;
  wire [9:0]  _slots_7_io_uop_fu_code;
  wire [1:0]  _slots_7_io_uop_iw_state;
  wire        _slots_7_io_uop_iw_p1_poisoned;
  wire        _slots_7_io_uop_iw_p2_poisoned;
  wire        _slots_7_io_uop_is_br;
  wire        _slots_7_io_uop_is_jalr;
  wire        _slots_7_io_uop_is_jal;
  wire        _slots_7_io_uop_is_sfb;
  wire [19:0] _slots_7_io_uop_br_mask;
  wire [4:0]  _slots_7_io_uop_br_tag;
  wire [5:0]  _slots_7_io_uop_ftq_idx;
  wire        _slots_7_io_uop_edge_inst;
  wire [5:0]  _slots_7_io_uop_pc_lob;
  wire        _slots_7_io_uop_taken;
  wire [19:0] _slots_7_io_uop_imm_packed;
  wire [11:0] _slots_7_io_uop_csr_addr;
  wire [6:0]  _slots_7_io_uop_rob_idx;
  wire [4:0]  _slots_7_io_uop_ldq_idx;
  wire [4:0]  _slots_7_io_uop_stq_idx;
  wire [1:0]  _slots_7_io_uop_rxq_idx;
  wire [6:0]  _slots_7_io_uop_pdst;
  wire [6:0]  _slots_7_io_uop_prs1;
  wire [6:0]  _slots_7_io_uop_prs2;
  wire [6:0]  _slots_7_io_uop_prs3;
  wire [5:0]  _slots_7_io_uop_ppred;
  wire        _slots_7_io_uop_prs1_busy;
  wire        _slots_7_io_uop_prs2_busy;
  wire        _slots_7_io_uop_prs3_busy;
  wire        _slots_7_io_uop_ppred_busy;
  wire [6:0]  _slots_7_io_uop_stale_pdst;
  wire        _slots_7_io_uop_exception;
  wire [63:0] _slots_7_io_uop_exc_cause;
  wire        _slots_7_io_uop_bypassable;
  wire [4:0]  _slots_7_io_uop_mem_cmd;
  wire [1:0]  _slots_7_io_uop_mem_size;
  wire        _slots_7_io_uop_mem_signed;
  wire        _slots_7_io_uop_is_fence;
  wire        _slots_7_io_uop_is_fencei;
  wire        _slots_7_io_uop_is_amo;
  wire        _slots_7_io_uop_uses_ldq;
  wire        _slots_7_io_uop_uses_stq;
  wire        _slots_7_io_uop_is_sys_pc2epc;
  wire        _slots_7_io_uop_is_unique;
  wire        _slots_7_io_uop_flush_on_commit;
  wire        _slots_7_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_7_io_uop_ldst;
  wire [5:0]  _slots_7_io_uop_lrs1;
  wire [5:0]  _slots_7_io_uop_lrs2;
  wire [5:0]  _slots_7_io_uop_lrs3;
  wire        _slots_7_io_uop_ldst_val;
  wire [1:0]  _slots_7_io_uop_dst_rtype;
  wire [1:0]  _slots_7_io_uop_lrs1_rtype;
  wire [1:0]  _slots_7_io_uop_lrs2_rtype;
  wire        _slots_7_io_uop_frs3_en;
  wire        _slots_7_io_uop_fp_val;
  wire        _slots_7_io_uop_fp_single;
  wire        _slots_7_io_uop_xcpt_pf_if;
  wire        _slots_7_io_uop_xcpt_ae_if;
  wire        _slots_7_io_uop_xcpt_ma_if;
  wire        _slots_7_io_uop_bp_debug_if;
  wire        _slots_7_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_7_io_uop_debug_fsrc;
  wire [1:0]  _slots_7_io_uop_debug_tsrc;
  wire        _slots_6_io_valid;
  wire        _slots_6_io_will_be_valid;
  wire        _slots_6_io_request;
  wire [6:0]  _slots_6_io_out_uop_uopc;
  wire [31:0] _slots_6_io_out_uop_inst;
  wire [31:0] _slots_6_io_out_uop_debug_inst;
  wire        _slots_6_io_out_uop_is_rvc;
  wire [39:0] _slots_6_io_out_uop_debug_pc;
  wire [2:0]  _slots_6_io_out_uop_iq_type;
  wire [9:0]  _slots_6_io_out_uop_fu_code;
  wire [1:0]  _slots_6_io_out_uop_iw_state;
  wire        _slots_6_io_out_uop_iw_p1_poisoned;
  wire        _slots_6_io_out_uop_iw_p2_poisoned;
  wire        _slots_6_io_out_uop_is_br;
  wire        _slots_6_io_out_uop_is_jalr;
  wire        _slots_6_io_out_uop_is_jal;
  wire        _slots_6_io_out_uop_is_sfb;
  wire [19:0] _slots_6_io_out_uop_br_mask;
  wire [4:0]  _slots_6_io_out_uop_br_tag;
  wire [5:0]  _slots_6_io_out_uop_ftq_idx;
  wire        _slots_6_io_out_uop_edge_inst;
  wire [5:0]  _slots_6_io_out_uop_pc_lob;
  wire        _slots_6_io_out_uop_taken;
  wire [19:0] _slots_6_io_out_uop_imm_packed;
  wire [11:0] _slots_6_io_out_uop_csr_addr;
  wire [6:0]  _slots_6_io_out_uop_rob_idx;
  wire [4:0]  _slots_6_io_out_uop_ldq_idx;
  wire [4:0]  _slots_6_io_out_uop_stq_idx;
  wire [1:0]  _slots_6_io_out_uop_rxq_idx;
  wire [6:0]  _slots_6_io_out_uop_pdst;
  wire [6:0]  _slots_6_io_out_uop_prs1;
  wire [6:0]  _slots_6_io_out_uop_prs2;
  wire [6:0]  _slots_6_io_out_uop_prs3;
  wire [5:0]  _slots_6_io_out_uop_ppred;
  wire        _slots_6_io_out_uop_prs1_busy;
  wire        _slots_6_io_out_uop_prs2_busy;
  wire        _slots_6_io_out_uop_prs3_busy;
  wire        _slots_6_io_out_uop_ppred_busy;
  wire [6:0]  _slots_6_io_out_uop_stale_pdst;
  wire        _slots_6_io_out_uop_exception;
  wire [63:0] _slots_6_io_out_uop_exc_cause;
  wire        _slots_6_io_out_uop_bypassable;
  wire [4:0]  _slots_6_io_out_uop_mem_cmd;
  wire [1:0]  _slots_6_io_out_uop_mem_size;
  wire        _slots_6_io_out_uop_mem_signed;
  wire        _slots_6_io_out_uop_is_fence;
  wire        _slots_6_io_out_uop_is_fencei;
  wire        _slots_6_io_out_uop_is_amo;
  wire        _slots_6_io_out_uop_uses_ldq;
  wire        _slots_6_io_out_uop_uses_stq;
  wire        _slots_6_io_out_uop_is_sys_pc2epc;
  wire        _slots_6_io_out_uop_is_unique;
  wire        _slots_6_io_out_uop_flush_on_commit;
  wire        _slots_6_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_6_io_out_uop_ldst;
  wire [5:0]  _slots_6_io_out_uop_lrs1;
  wire [5:0]  _slots_6_io_out_uop_lrs2;
  wire [5:0]  _slots_6_io_out_uop_lrs3;
  wire        _slots_6_io_out_uop_ldst_val;
  wire [1:0]  _slots_6_io_out_uop_dst_rtype;
  wire [1:0]  _slots_6_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_6_io_out_uop_lrs2_rtype;
  wire        _slots_6_io_out_uop_frs3_en;
  wire        _slots_6_io_out_uop_fp_val;
  wire        _slots_6_io_out_uop_fp_single;
  wire        _slots_6_io_out_uop_xcpt_pf_if;
  wire        _slots_6_io_out_uop_xcpt_ae_if;
  wire        _slots_6_io_out_uop_xcpt_ma_if;
  wire        _slots_6_io_out_uop_bp_debug_if;
  wire        _slots_6_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_6_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_6_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_6_io_uop_uopc;
  wire [31:0] _slots_6_io_uop_inst;
  wire [31:0] _slots_6_io_uop_debug_inst;
  wire        _slots_6_io_uop_is_rvc;
  wire [39:0] _slots_6_io_uop_debug_pc;
  wire [2:0]  _slots_6_io_uop_iq_type;
  wire [9:0]  _slots_6_io_uop_fu_code;
  wire [1:0]  _slots_6_io_uop_iw_state;
  wire        _slots_6_io_uop_iw_p1_poisoned;
  wire        _slots_6_io_uop_iw_p2_poisoned;
  wire        _slots_6_io_uop_is_br;
  wire        _slots_6_io_uop_is_jalr;
  wire        _slots_6_io_uop_is_jal;
  wire        _slots_6_io_uop_is_sfb;
  wire [19:0] _slots_6_io_uop_br_mask;
  wire [4:0]  _slots_6_io_uop_br_tag;
  wire [5:0]  _slots_6_io_uop_ftq_idx;
  wire        _slots_6_io_uop_edge_inst;
  wire [5:0]  _slots_6_io_uop_pc_lob;
  wire        _slots_6_io_uop_taken;
  wire [19:0] _slots_6_io_uop_imm_packed;
  wire [11:0] _slots_6_io_uop_csr_addr;
  wire [6:0]  _slots_6_io_uop_rob_idx;
  wire [4:0]  _slots_6_io_uop_ldq_idx;
  wire [4:0]  _slots_6_io_uop_stq_idx;
  wire [1:0]  _slots_6_io_uop_rxq_idx;
  wire [6:0]  _slots_6_io_uop_pdst;
  wire [6:0]  _slots_6_io_uop_prs1;
  wire [6:0]  _slots_6_io_uop_prs2;
  wire [6:0]  _slots_6_io_uop_prs3;
  wire [5:0]  _slots_6_io_uop_ppred;
  wire        _slots_6_io_uop_prs1_busy;
  wire        _slots_6_io_uop_prs2_busy;
  wire        _slots_6_io_uop_prs3_busy;
  wire        _slots_6_io_uop_ppred_busy;
  wire [6:0]  _slots_6_io_uop_stale_pdst;
  wire        _slots_6_io_uop_exception;
  wire [63:0] _slots_6_io_uop_exc_cause;
  wire        _slots_6_io_uop_bypassable;
  wire [4:0]  _slots_6_io_uop_mem_cmd;
  wire [1:0]  _slots_6_io_uop_mem_size;
  wire        _slots_6_io_uop_mem_signed;
  wire        _slots_6_io_uop_is_fence;
  wire        _slots_6_io_uop_is_fencei;
  wire        _slots_6_io_uop_is_amo;
  wire        _slots_6_io_uop_uses_ldq;
  wire        _slots_6_io_uop_uses_stq;
  wire        _slots_6_io_uop_is_sys_pc2epc;
  wire        _slots_6_io_uop_is_unique;
  wire        _slots_6_io_uop_flush_on_commit;
  wire        _slots_6_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_6_io_uop_ldst;
  wire [5:0]  _slots_6_io_uop_lrs1;
  wire [5:0]  _slots_6_io_uop_lrs2;
  wire [5:0]  _slots_6_io_uop_lrs3;
  wire        _slots_6_io_uop_ldst_val;
  wire [1:0]  _slots_6_io_uop_dst_rtype;
  wire [1:0]  _slots_6_io_uop_lrs1_rtype;
  wire [1:0]  _slots_6_io_uop_lrs2_rtype;
  wire        _slots_6_io_uop_frs3_en;
  wire        _slots_6_io_uop_fp_val;
  wire        _slots_6_io_uop_fp_single;
  wire        _slots_6_io_uop_xcpt_pf_if;
  wire        _slots_6_io_uop_xcpt_ae_if;
  wire        _slots_6_io_uop_xcpt_ma_if;
  wire        _slots_6_io_uop_bp_debug_if;
  wire        _slots_6_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_6_io_uop_debug_fsrc;
  wire [1:0]  _slots_6_io_uop_debug_tsrc;
  wire        _slots_5_io_valid;
  wire        _slots_5_io_will_be_valid;
  wire        _slots_5_io_request;
  wire [6:0]  _slots_5_io_out_uop_uopc;
  wire [31:0] _slots_5_io_out_uop_inst;
  wire [31:0] _slots_5_io_out_uop_debug_inst;
  wire        _slots_5_io_out_uop_is_rvc;
  wire [39:0] _slots_5_io_out_uop_debug_pc;
  wire [2:0]  _slots_5_io_out_uop_iq_type;
  wire [9:0]  _slots_5_io_out_uop_fu_code;
  wire [1:0]  _slots_5_io_out_uop_iw_state;
  wire        _slots_5_io_out_uop_iw_p1_poisoned;
  wire        _slots_5_io_out_uop_iw_p2_poisoned;
  wire        _slots_5_io_out_uop_is_br;
  wire        _slots_5_io_out_uop_is_jalr;
  wire        _slots_5_io_out_uop_is_jal;
  wire        _slots_5_io_out_uop_is_sfb;
  wire [19:0] _slots_5_io_out_uop_br_mask;
  wire [4:0]  _slots_5_io_out_uop_br_tag;
  wire [5:0]  _slots_5_io_out_uop_ftq_idx;
  wire        _slots_5_io_out_uop_edge_inst;
  wire [5:0]  _slots_5_io_out_uop_pc_lob;
  wire        _slots_5_io_out_uop_taken;
  wire [19:0] _slots_5_io_out_uop_imm_packed;
  wire [11:0] _slots_5_io_out_uop_csr_addr;
  wire [6:0]  _slots_5_io_out_uop_rob_idx;
  wire [4:0]  _slots_5_io_out_uop_ldq_idx;
  wire [4:0]  _slots_5_io_out_uop_stq_idx;
  wire [1:0]  _slots_5_io_out_uop_rxq_idx;
  wire [6:0]  _slots_5_io_out_uop_pdst;
  wire [6:0]  _slots_5_io_out_uop_prs1;
  wire [6:0]  _slots_5_io_out_uop_prs2;
  wire [6:0]  _slots_5_io_out_uop_prs3;
  wire [5:0]  _slots_5_io_out_uop_ppred;
  wire        _slots_5_io_out_uop_prs1_busy;
  wire        _slots_5_io_out_uop_prs2_busy;
  wire        _slots_5_io_out_uop_prs3_busy;
  wire        _slots_5_io_out_uop_ppred_busy;
  wire [6:0]  _slots_5_io_out_uop_stale_pdst;
  wire        _slots_5_io_out_uop_exception;
  wire [63:0] _slots_5_io_out_uop_exc_cause;
  wire        _slots_5_io_out_uop_bypassable;
  wire [4:0]  _slots_5_io_out_uop_mem_cmd;
  wire [1:0]  _slots_5_io_out_uop_mem_size;
  wire        _slots_5_io_out_uop_mem_signed;
  wire        _slots_5_io_out_uop_is_fence;
  wire        _slots_5_io_out_uop_is_fencei;
  wire        _slots_5_io_out_uop_is_amo;
  wire        _slots_5_io_out_uop_uses_ldq;
  wire        _slots_5_io_out_uop_uses_stq;
  wire        _slots_5_io_out_uop_is_sys_pc2epc;
  wire        _slots_5_io_out_uop_is_unique;
  wire        _slots_5_io_out_uop_flush_on_commit;
  wire        _slots_5_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_5_io_out_uop_ldst;
  wire [5:0]  _slots_5_io_out_uop_lrs1;
  wire [5:0]  _slots_5_io_out_uop_lrs2;
  wire [5:0]  _slots_5_io_out_uop_lrs3;
  wire        _slots_5_io_out_uop_ldst_val;
  wire [1:0]  _slots_5_io_out_uop_dst_rtype;
  wire [1:0]  _slots_5_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_5_io_out_uop_lrs2_rtype;
  wire        _slots_5_io_out_uop_frs3_en;
  wire        _slots_5_io_out_uop_fp_val;
  wire        _slots_5_io_out_uop_fp_single;
  wire        _slots_5_io_out_uop_xcpt_pf_if;
  wire        _slots_5_io_out_uop_xcpt_ae_if;
  wire        _slots_5_io_out_uop_xcpt_ma_if;
  wire        _slots_5_io_out_uop_bp_debug_if;
  wire        _slots_5_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_5_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_5_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_5_io_uop_uopc;
  wire [31:0] _slots_5_io_uop_inst;
  wire [31:0] _slots_5_io_uop_debug_inst;
  wire        _slots_5_io_uop_is_rvc;
  wire [39:0] _slots_5_io_uop_debug_pc;
  wire [2:0]  _slots_5_io_uop_iq_type;
  wire [9:0]  _slots_5_io_uop_fu_code;
  wire [1:0]  _slots_5_io_uop_iw_state;
  wire        _slots_5_io_uop_iw_p1_poisoned;
  wire        _slots_5_io_uop_iw_p2_poisoned;
  wire        _slots_5_io_uop_is_br;
  wire        _slots_5_io_uop_is_jalr;
  wire        _slots_5_io_uop_is_jal;
  wire        _slots_5_io_uop_is_sfb;
  wire [19:0] _slots_5_io_uop_br_mask;
  wire [4:0]  _slots_5_io_uop_br_tag;
  wire [5:0]  _slots_5_io_uop_ftq_idx;
  wire        _slots_5_io_uop_edge_inst;
  wire [5:0]  _slots_5_io_uop_pc_lob;
  wire        _slots_5_io_uop_taken;
  wire [19:0] _slots_5_io_uop_imm_packed;
  wire [11:0] _slots_5_io_uop_csr_addr;
  wire [6:0]  _slots_5_io_uop_rob_idx;
  wire [4:0]  _slots_5_io_uop_ldq_idx;
  wire [4:0]  _slots_5_io_uop_stq_idx;
  wire [1:0]  _slots_5_io_uop_rxq_idx;
  wire [6:0]  _slots_5_io_uop_pdst;
  wire [6:0]  _slots_5_io_uop_prs1;
  wire [6:0]  _slots_5_io_uop_prs2;
  wire [6:0]  _slots_5_io_uop_prs3;
  wire [5:0]  _slots_5_io_uop_ppred;
  wire        _slots_5_io_uop_prs1_busy;
  wire        _slots_5_io_uop_prs2_busy;
  wire        _slots_5_io_uop_prs3_busy;
  wire        _slots_5_io_uop_ppred_busy;
  wire [6:0]  _slots_5_io_uop_stale_pdst;
  wire        _slots_5_io_uop_exception;
  wire [63:0] _slots_5_io_uop_exc_cause;
  wire        _slots_5_io_uop_bypassable;
  wire [4:0]  _slots_5_io_uop_mem_cmd;
  wire [1:0]  _slots_5_io_uop_mem_size;
  wire        _slots_5_io_uop_mem_signed;
  wire        _slots_5_io_uop_is_fence;
  wire        _slots_5_io_uop_is_fencei;
  wire        _slots_5_io_uop_is_amo;
  wire        _slots_5_io_uop_uses_ldq;
  wire        _slots_5_io_uop_uses_stq;
  wire        _slots_5_io_uop_is_sys_pc2epc;
  wire        _slots_5_io_uop_is_unique;
  wire        _slots_5_io_uop_flush_on_commit;
  wire        _slots_5_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_5_io_uop_ldst;
  wire [5:0]  _slots_5_io_uop_lrs1;
  wire [5:0]  _slots_5_io_uop_lrs2;
  wire [5:0]  _slots_5_io_uop_lrs3;
  wire        _slots_5_io_uop_ldst_val;
  wire [1:0]  _slots_5_io_uop_dst_rtype;
  wire [1:0]  _slots_5_io_uop_lrs1_rtype;
  wire [1:0]  _slots_5_io_uop_lrs2_rtype;
  wire        _slots_5_io_uop_frs3_en;
  wire        _slots_5_io_uop_fp_val;
  wire        _slots_5_io_uop_fp_single;
  wire        _slots_5_io_uop_xcpt_pf_if;
  wire        _slots_5_io_uop_xcpt_ae_if;
  wire        _slots_5_io_uop_xcpt_ma_if;
  wire        _slots_5_io_uop_bp_debug_if;
  wire        _slots_5_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_5_io_uop_debug_fsrc;
  wire [1:0]  _slots_5_io_uop_debug_tsrc;
  wire        _slots_4_io_valid;
  wire        _slots_4_io_will_be_valid;
  wire        _slots_4_io_request;
  wire [6:0]  _slots_4_io_out_uop_uopc;
  wire [31:0] _slots_4_io_out_uop_inst;
  wire [31:0] _slots_4_io_out_uop_debug_inst;
  wire        _slots_4_io_out_uop_is_rvc;
  wire [39:0] _slots_4_io_out_uop_debug_pc;
  wire [2:0]  _slots_4_io_out_uop_iq_type;
  wire [9:0]  _slots_4_io_out_uop_fu_code;
  wire [1:0]  _slots_4_io_out_uop_iw_state;
  wire        _slots_4_io_out_uop_iw_p1_poisoned;
  wire        _slots_4_io_out_uop_iw_p2_poisoned;
  wire        _slots_4_io_out_uop_is_br;
  wire        _slots_4_io_out_uop_is_jalr;
  wire        _slots_4_io_out_uop_is_jal;
  wire        _slots_4_io_out_uop_is_sfb;
  wire [19:0] _slots_4_io_out_uop_br_mask;
  wire [4:0]  _slots_4_io_out_uop_br_tag;
  wire [5:0]  _slots_4_io_out_uop_ftq_idx;
  wire        _slots_4_io_out_uop_edge_inst;
  wire [5:0]  _slots_4_io_out_uop_pc_lob;
  wire        _slots_4_io_out_uop_taken;
  wire [19:0] _slots_4_io_out_uop_imm_packed;
  wire [11:0] _slots_4_io_out_uop_csr_addr;
  wire [6:0]  _slots_4_io_out_uop_rob_idx;
  wire [4:0]  _slots_4_io_out_uop_ldq_idx;
  wire [4:0]  _slots_4_io_out_uop_stq_idx;
  wire [1:0]  _slots_4_io_out_uop_rxq_idx;
  wire [6:0]  _slots_4_io_out_uop_pdst;
  wire [6:0]  _slots_4_io_out_uop_prs1;
  wire [6:0]  _slots_4_io_out_uop_prs2;
  wire [6:0]  _slots_4_io_out_uop_prs3;
  wire [5:0]  _slots_4_io_out_uop_ppred;
  wire        _slots_4_io_out_uop_prs1_busy;
  wire        _slots_4_io_out_uop_prs2_busy;
  wire        _slots_4_io_out_uop_prs3_busy;
  wire        _slots_4_io_out_uop_ppred_busy;
  wire [6:0]  _slots_4_io_out_uop_stale_pdst;
  wire        _slots_4_io_out_uop_exception;
  wire [63:0] _slots_4_io_out_uop_exc_cause;
  wire        _slots_4_io_out_uop_bypassable;
  wire [4:0]  _slots_4_io_out_uop_mem_cmd;
  wire [1:0]  _slots_4_io_out_uop_mem_size;
  wire        _slots_4_io_out_uop_mem_signed;
  wire        _slots_4_io_out_uop_is_fence;
  wire        _slots_4_io_out_uop_is_fencei;
  wire        _slots_4_io_out_uop_is_amo;
  wire        _slots_4_io_out_uop_uses_ldq;
  wire        _slots_4_io_out_uop_uses_stq;
  wire        _slots_4_io_out_uop_is_sys_pc2epc;
  wire        _slots_4_io_out_uop_is_unique;
  wire        _slots_4_io_out_uop_flush_on_commit;
  wire        _slots_4_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_4_io_out_uop_ldst;
  wire [5:0]  _slots_4_io_out_uop_lrs1;
  wire [5:0]  _slots_4_io_out_uop_lrs2;
  wire [5:0]  _slots_4_io_out_uop_lrs3;
  wire        _slots_4_io_out_uop_ldst_val;
  wire [1:0]  _slots_4_io_out_uop_dst_rtype;
  wire [1:0]  _slots_4_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_4_io_out_uop_lrs2_rtype;
  wire        _slots_4_io_out_uop_frs3_en;
  wire        _slots_4_io_out_uop_fp_val;
  wire        _slots_4_io_out_uop_fp_single;
  wire        _slots_4_io_out_uop_xcpt_pf_if;
  wire        _slots_4_io_out_uop_xcpt_ae_if;
  wire        _slots_4_io_out_uop_xcpt_ma_if;
  wire        _slots_4_io_out_uop_bp_debug_if;
  wire        _slots_4_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_4_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_4_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_4_io_uop_uopc;
  wire [31:0] _slots_4_io_uop_inst;
  wire [31:0] _slots_4_io_uop_debug_inst;
  wire        _slots_4_io_uop_is_rvc;
  wire [39:0] _slots_4_io_uop_debug_pc;
  wire [2:0]  _slots_4_io_uop_iq_type;
  wire [9:0]  _slots_4_io_uop_fu_code;
  wire [1:0]  _slots_4_io_uop_iw_state;
  wire        _slots_4_io_uop_iw_p1_poisoned;
  wire        _slots_4_io_uop_iw_p2_poisoned;
  wire        _slots_4_io_uop_is_br;
  wire        _slots_4_io_uop_is_jalr;
  wire        _slots_4_io_uop_is_jal;
  wire        _slots_4_io_uop_is_sfb;
  wire [19:0] _slots_4_io_uop_br_mask;
  wire [4:0]  _slots_4_io_uop_br_tag;
  wire [5:0]  _slots_4_io_uop_ftq_idx;
  wire        _slots_4_io_uop_edge_inst;
  wire [5:0]  _slots_4_io_uop_pc_lob;
  wire        _slots_4_io_uop_taken;
  wire [19:0] _slots_4_io_uop_imm_packed;
  wire [11:0] _slots_4_io_uop_csr_addr;
  wire [6:0]  _slots_4_io_uop_rob_idx;
  wire [4:0]  _slots_4_io_uop_ldq_idx;
  wire [4:0]  _slots_4_io_uop_stq_idx;
  wire [1:0]  _slots_4_io_uop_rxq_idx;
  wire [6:0]  _slots_4_io_uop_pdst;
  wire [6:0]  _slots_4_io_uop_prs1;
  wire [6:0]  _slots_4_io_uop_prs2;
  wire [6:0]  _slots_4_io_uop_prs3;
  wire [5:0]  _slots_4_io_uop_ppred;
  wire        _slots_4_io_uop_prs1_busy;
  wire        _slots_4_io_uop_prs2_busy;
  wire        _slots_4_io_uop_prs3_busy;
  wire        _slots_4_io_uop_ppred_busy;
  wire [6:0]  _slots_4_io_uop_stale_pdst;
  wire        _slots_4_io_uop_exception;
  wire [63:0] _slots_4_io_uop_exc_cause;
  wire        _slots_4_io_uop_bypassable;
  wire [4:0]  _slots_4_io_uop_mem_cmd;
  wire [1:0]  _slots_4_io_uop_mem_size;
  wire        _slots_4_io_uop_mem_signed;
  wire        _slots_4_io_uop_is_fence;
  wire        _slots_4_io_uop_is_fencei;
  wire        _slots_4_io_uop_is_amo;
  wire        _slots_4_io_uop_uses_ldq;
  wire        _slots_4_io_uop_uses_stq;
  wire        _slots_4_io_uop_is_sys_pc2epc;
  wire        _slots_4_io_uop_is_unique;
  wire        _slots_4_io_uop_flush_on_commit;
  wire        _slots_4_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_4_io_uop_ldst;
  wire [5:0]  _slots_4_io_uop_lrs1;
  wire [5:0]  _slots_4_io_uop_lrs2;
  wire [5:0]  _slots_4_io_uop_lrs3;
  wire        _slots_4_io_uop_ldst_val;
  wire [1:0]  _slots_4_io_uop_dst_rtype;
  wire [1:0]  _slots_4_io_uop_lrs1_rtype;
  wire [1:0]  _slots_4_io_uop_lrs2_rtype;
  wire        _slots_4_io_uop_frs3_en;
  wire        _slots_4_io_uop_fp_val;
  wire        _slots_4_io_uop_fp_single;
  wire        _slots_4_io_uop_xcpt_pf_if;
  wire        _slots_4_io_uop_xcpt_ae_if;
  wire        _slots_4_io_uop_xcpt_ma_if;
  wire        _slots_4_io_uop_bp_debug_if;
  wire        _slots_4_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_4_io_uop_debug_fsrc;
  wire [1:0]  _slots_4_io_uop_debug_tsrc;
  wire        _slots_3_io_valid;
  wire        _slots_3_io_will_be_valid;
  wire        _slots_3_io_request;
  wire [6:0]  _slots_3_io_out_uop_uopc;
  wire [31:0] _slots_3_io_out_uop_inst;
  wire [31:0] _slots_3_io_out_uop_debug_inst;
  wire        _slots_3_io_out_uop_is_rvc;
  wire [39:0] _slots_3_io_out_uop_debug_pc;
  wire [2:0]  _slots_3_io_out_uop_iq_type;
  wire [9:0]  _slots_3_io_out_uop_fu_code;
  wire [1:0]  _slots_3_io_out_uop_iw_state;
  wire        _slots_3_io_out_uop_iw_p1_poisoned;
  wire        _slots_3_io_out_uop_iw_p2_poisoned;
  wire        _slots_3_io_out_uop_is_br;
  wire        _slots_3_io_out_uop_is_jalr;
  wire        _slots_3_io_out_uop_is_jal;
  wire        _slots_3_io_out_uop_is_sfb;
  wire [19:0] _slots_3_io_out_uop_br_mask;
  wire [4:0]  _slots_3_io_out_uop_br_tag;
  wire [5:0]  _slots_3_io_out_uop_ftq_idx;
  wire        _slots_3_io_out_uop_edge_inst;
  wire [5:0]  _slots_3_io_out_uop_pc_lob;
  wire        _slots_3_io_out_uop_taken;
  wire [19:0] _slots_3_io_out_uop_imm_packed;
  wire [11:0] _slots_3_io_out_uop_csr_addr;
  wire [6:0]  _slots_3_io_out_uop_rob_idx;
  wire [4:0]  _slots_3_io_out_uop_ldq_idx;
  wire [4:0]  _slots_3_io_out_uop_stq_idx;
  wire [1:0]  _slots_3_io_out_uop_rxq_idx;
  wire [6:0]  _slots_3_io_out_uop_pdst;
  wire [6:0]  _slots_3_io_out_uop_prs1;
  wire [6:0]  _slots_3_io_out_uop_prs2;
  wire [6:0]  _slots_3_io_out_uop_prs3;
  wire [5:0]  _slots_3_io_out_uop_ppred;
  wire        _slots_3_io_out_uop_prs1_busy;
  wire        _slots_3_io_out_uop_prs2_busy;
  wire        _slots_3_io_out_uop_prs3_busy;
  wire        _slots_3_io_out_uop_ppred_busy;
  wire [6:0]  _slots_3_io_out_uop_stale_pdst;
  wire        _slots_3_io_out_uop_exception;
  wire [63:0] _slots_3_io_out_uop_exc_cause;
  wire        _slots_3_io_out_uop_bypassable;
  wire [4:0]  _slots_3_io_out_uop_mem_cmd;
  wire [1:0]  _slots_3_io_out_uop_mem_size;
  wire        _slots_3_io_out_uop_mem_signed;
  wire        _slots_3_io_out_uop_is_fence;
  wire        _slots_3_io_out_uop_is_fencei;
  wire        _slots_3_io_out_uop_is_amo;
  wire        _slots_3_io_out_uop_uses_ldq;
  wire        _slots_3_io_out_uop_uses_stq;
  wire        _slots_3_io_out_uop_is_sys_pc2epc;
  wire        _slots_3_io_out_uop_is_unique;
  wire        _slots_3_io_out_uop_flush_on_commit;
  wire        _slots_3_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_3_io_out_uop_ldst;
  wire [5:0]  _slots_3_io_out_uop_lrs1;
  wire [5:0]  _slots_3_io_out_uop_lrs2;
  wire [5:0]  _slots_3_io_out_uop_lrs3;
  wire        _slots_3_io_out_uop_ldst_val;
  wire [1:0]  _slots_3_io_out_uop_dst_rtype;
  wire [1:0]  _slots_3_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_3_io_out_uop_lrs2_rtype;
  wire        _slots_3_io_out_uop_frs3_en;
  wire        _slots_3_io_out_uop_fp_val;
  wire        _slots_3_io_out_uop_fp_single;
  wire        _slots_3_io_out_uop_xcpt_pf_if;
  wire        _slots_3_io_out_uop_xcpt_ae_if;
  wire        _slots_3_io_out_uop_xcpt_ma_if;
  wire        _slots_3_io_out_uop_bp_debug_if;
  wire        _slots_3_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_3_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_3_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_3_io_uop_uopc;
  wire [31:0] _slots_3_io_uop_inst;
  wire [31:0] _slots_3_io_uop_debug_inst;
  wire        _slots_3_io_uop_is_rvc;
  wire [39:0] _slots_3_io_uop_debug_pc;
  wire [2:0]  _slots_3_io_uop_iq_type;
  wire [9:0]  _slots_3_io_uop_fu_code;
  wire [1:0]  _slots_3_io_uop_iw_state;
  wire        _slots_3_io_uop_iw_p1_poisoned;
  wire        _slots_3_io_uop_iw_p2_poisoned;
  wire        _slots_3_io_uop_is_br;
  wire        _slots_3_io_uop_is_jalr;
  wire        _slots_3_io_uop_is_jal;
  wire        _slots_3_io_uop_is_sfb;
  wire [19:0] _slots_3_io_uop_br_mask;
  wire [4:0]  _slots_3_io_uop_br_tag;
  wire [5:0]  _slots_3_io_uop_ftq_idx;
  wire        _slots_3_io_uop_edge_inst;
  wire [5:0]  _slots_3_io_uop_pc_lob;
  wire        _slots_3_io_uop_taken;
  wire [19:0] _slots_3_io_uop_imm_packed;
  wire [11:0] _slots_3_io_uop_csr_addr;
  wire [6:0]  _slots_3_io_uop_rob_idx;
  wire [4:0]  _slots_3_io_uop_ldq_idx;
  wire [4:0]  _slots_3_io_uop_stq_idx;
  wire [1:0]  _slots_3_io_uop_rxq_idx;
  wire [6:0]  _slots_3_io_uop_pdst;
  wire [6:0]  _slots_3_io_uop_prs1;
  wire [6:0]  _slots_3_io_uop_prs2;
  wire [6:0]  _slots_3_io_uop_prs3;
  wire [5:0]  _slots_3_io_uop_ppred;
  wire        _slots_3_io_uop_prs1_busy;
  wire        _slots_3_io_uop_prs2_busy;
  wire        _slots_3_io_uop_prs3_busy;
  wire        _slots_3_io_uop_ppred_busy;
  wire [6:0]  _slots_3_io_uop_stale_pdst;
  wire        _slots_3_io_uop_exception;
  wire [63:0] _slots_3_io_uop_exc_cause;
  wire        _slots_3_io_uop_bypassable;
  wire [4:0]  _slots_3_io_uop_mem_cmd;
  wire [1:0]  _slots_3_io_uop_mem_size;
  wire        _slots_3_io_uop_mem_signed;
  wire        _slots_3_io_uop_is_fence;
  wire        _slots_3_io_uop_is_fencei;
  wire        _slots_3_io_uop_is_amo;
  wire        _slots_3_io_uop_uses_ldq;
  wire        _slots_3_io_uop_uses_stq;
  wire        _slots_3_io_uop_is_sys_pc2epc;
  wire        _slots_3_io_uop_is_unique;
  wire        _slots_3_io_uop_flush_on_commit;
  wire        _slots_3_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_3_io_uop_ldst;
  wire [5:0]  _slots_3_io_uop_lrs1;
  wire [5:0]  _slots_3_io_uop_lrs2;
  wire [5:0]  _slots_3_io_uop_lrs3;
  wire        _slots_3_io_uop_ldst_val;
  wire [1:0]  _slots_3_io_uop_dst_rtype;
  wire [1:0]  _slots_3_io_uop_lrs1_rtype;
  wire [1:0]  _slots_3_io_uop_lrs2_rtype;
  wire        _slots_3_io_uop_frs3_en;
  wire        _slots_3_io_uop_fp_val;
  wire        _slots_3_io_uop_fp_single;
  wire        _slots_3_io_uop_xcpt_pf_if;
  wire        _slots_3_io_uop_xcpt_ae_if;
  wire        _slots_3_io_uop_xcpt_ma_if;
  wire        _slots_3_io_uop_bp_debug_if;
  wire        _slots_3_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_3_io_uop_debug_fsrc;
  wire [1:0]  _slots_3_io_uop_debug_tsrc;
  wire        _slots_2_io_valid;
  wire        _slots_2_io_will_be_valid;
  wire        _slots_2_io_request;
  wire [6:0]  _slots_2_io_out_uop_uopc;
  wire [31:0] _slots_2_io_out_uop_inst;
  wire [31:0] _slots_2_io_out_uop_debug_inst;
  wire        _slots_2_io_out_uop_is_rvc;
  wire [39:0] _slots_2_io_out_uop_debug_pc;
  wire [2:0]  _slots_2_io_out_uop_iq_type;
  wire [9:0]  _slots_2_io_out_uop_fu_code;
  wire [1:0]  _slots_2_io_out_uop_iw_state;
  wire        _slots_2_io_out_uop_iw_p1_poisoned;
  wire        _slots_2_io_out_uop_iw_p2_poisoned;
  wire        _slots_2_io_out_uop_is_br;
  wire        _slots_2_io_out_uop_is_jalr;
  wire        _slots_2_io_out_uop_is_jal;
  wire        _slots_2_io_out_uop_is_sfb;
  wire [19:0] _slots_2_io_out_uop_br_mask;
  wire [4:0]  _slots_2_io_out_uop_br_tag;
  wire [5:0]  _slots_2_io_out_uop_ftq_idx;
  wire        _slots_2_io_out_uop_edge_inst;
  wire [5:0]  _slots_2_io_out_uop_pc_lob;
  wire        _slots_2_io_out_uop_taken;
  wire [19:0] _slots_2_io_out_uop_imm_packed;
  wire [11:0] _slots_2_io_out_uop_csr_addr;
  wire [6:0]  _slots_2_io_out_uop_rob_idx;
  wire [4:0]  _slots_2_io_out_uop_ldq_idx;
  wire [4:0]  _slots_2_io_out_uop_stq_idx;
  wire [1:0]  _slots_2_io_out_uop_rxq_idx;
  wire [6:0]  _slots_2_io_out_uop_pdst;
  wire [6:0]  _slots_2_io_out_uop_prs1;
  wire [6:0]  _slots_2_io_out_uop_prs2;
  wire [6:0]  _slots_2_io_out_uop_prs3;
  wire [5:0]  _slots_2_io_out_uop_ppred;
  wire        _slots_2_io_out_uop_prs1_busy;
  wire        _slots_2_io_out_uop_prs2_busy;
  wire        _slots_2_io_out_uop_prs3_busy;
  wire        _slots_2_io_out_uop_ppred_busy;
  wire [6:0]  _slots_2_io_out_uop_stale_pdst;
  wire        _slots_2_io_out_uop_exception;
  wire [63:0] _slots_2_io_out_uop_exc_cause;
  wire        _slots_2_io_out_uop_bypassable;
  wire [4:0]  _slots_2_io_out_uop_mem_cmd;
  wire [1:0]  _slots_2_io_out_uop_mem_size;
  wire        _slots_2_io_out_uop_mem_signed;
  wire        _slots_2_io_out_uop_is_fence;
  wire        _slots_2_io_out_uop_is_fencei;
  wire        _slots_2_io_out_uop_is_amo;
  wire        _slots_2_io_out_uop_uses_ldq;
  wire        _slots_2_io_out_uop_uses_stq;
  wire        _slots_2_io_out_uop_is_sys_pc2epc;
  wire        _slots_2_io_out_uop_is_unique;
  wire        _slots_2_io_out_uop_flush_on_commit;
  wire        _slots_2_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_2_io_out_uop_ldst;
  wire [5:0]  _slots_2_io_out_uop_lrs1;
  wire [5:0]  _slots_2_io_out_uop_lrs2;
  wire [5:0]  _slots_2_io_out_uop_lrs3;
  wire        _slots_2_io_out_uop_ldst_val;
  wire [1:0]  _slots_2_io_out_uop_dst_rtype;
  wire [1:0]  _slots_2_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_2_io_out_uop_lrs2_rtype;
  wire        _slots_2_io_out_uop_frs3_en;
  wire        _slots_2_io_out_uop_fp_val;
  wire        _slots_2_io_out_uop_fp_single;
  wire        _slots_2_io_out_uop_xcpt_pf_if;
  wire        _slots_2_io_out_uop_xcpt_ae_if;
  wire        _slots_2_io_out_uop_xcpt_ma_if;
  wire        _slots_2_io_out_uop_bp_debug_if;
  wire        _slots_2_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_2_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_2_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_2_io_uop_uopc;
  wire [31:0] _slots_2_io_uop_inst;
  wire [31:0] _slots_2_io_uop_debug_inst;
  wire        _slots_2_io_uop_is_rvc;
  wire [39:0] _slots_2_io_uop_debug_pc;
  wire [2:0]  _slots_2_io_uop_iq_type;
  wire [9:0]  _slots_2_io_uop_fu_code;
  wire [1:0]  _slots_2_io_uop_iw_state;
  wire        _slots_2_io_uop_iw_p1_poisoned;
  wire        _slots_2_io_uop_iw_p2_poisoned;
  wire        _slots_2_io_uop_is_br;
  wire        _slots_2_io_uop_is_jalr;
  wire        _slots_2_io_uop_is_jal;
  wire        _slots_2_io_uop_is_sfb;
  wire [19:0] _slots_2_io_uop_br_mask;
  wire [4:0]  _slots_2_io_uop_br_tag;
  wire [5:0]  _slots_2_io_uop_ftq_idx;
  wire        _slots_2_io_uop_edge_inst;
  wire [5:0]  _slots_2_io_uop_pc_lob;
  wire        _slots_2_io_uop_taken;
  wire [19:0] _slots_2_io_uop_imm_packed;
  wire [11:0] _slots_2_io_uop_csr_addr;
  wire [6:0]  _slots_2_io_uop_rob_idx;
  wire [4:0]  _slots_2_io_uop_ldq_idx;
  wire [4:0]  _slots_2_io_uop_stq_idx;
  wire [1:0]  _slots_2_io_uop_rxq_idx;
  wire [6:0]  _slots_2_io_uop_pdst;
  wire [6:0]  _slots_2_io_uop_prs1;
  wire [6:0]  _slots_2_io_uop_prs2;
  wire [6:0]  _slots_2_io_uop_prs3;
  wire [5:0]  _slots_2_io_uop_ppred;
  wire        _slots_2_io_uop_prs1_busy;
  wire        _slots_2_io_uop_prs2_busy;
  wire        _slots_2_io_uop_prs3_busy;
  wire        _slots_2_io_uop_ppred_busy;
  wire [6:0]  _slots_2_io_uop_stale_pdst;
  wire        _slots_2_io_uop_exception;
  wire [63:0] _slots_2_io_uop_exc_cause;
  wire        _slots_2_io_uop_bypassable;
  wire [4:0]  _slots_2_io_uop_mem_cmd;
  wire [1:0]  _slots_2_io_uop_mem_size;
  wire        _slots_2_io_uop_mem_signed;
  wire        _slots_2_io_uop_is_fence;
  wire        _slots_2_io_uop_is_fencei;
  wire        _slots_2_io_uop_is_amo;
  wire        _slots_2_io_uop_uses_ldq;
  wire        _slots_2_io_uop_uses_stq;
  wire        _slots_2_io_uop_is_sys_pc2epc;
  wire        _slots_2_io_uop_is_unique;
  wire        _slots_2_io_uop_flush_on_commit;
  wire        _slots_2_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_2_io_uop_ldst;
  wire [5:0]  _slots_2_io_uop_lrs1;
  wire [5:0]  _slots_2_io_uop_lrs2;
  wire [5:0]  _slots_2_io_uop_lrs3;
  wire        _slots_2_io_uop_ldst_val;
  wire [1:0]  _slots_2_io_uop_dst_rtype;
  wire [1:0]  _slots_2_io_uop_lrs1_rtype;
  wire [1:0]  _slots_2_io_uop_lrs2_rtype;
  wire        _slots_2_io_uop_frs3_en;
  wire        _slots_2_io_uop_fp_val;
  wire        _slots_2_io_uop_fp_single;
  wire        _slots_2_io_uop_xcpt_pf_if;
  wire        _slots_2_io_uop_xcpt_ae_if;
  wire        _slots_2_io_uop_xcpt_ma_if;
  wire        _slots_2_io_uop_bp_debug_if;
  wire        _slots_2_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_2_io_uop_debug_fsrc;
  wire [1:0]  _slots_2_io_uop_debug_tsrc;
  wire        _slots_1_io_valid;
  wire        _slots_1_io_will_be_valid;
  wire        _slots_1_io_request;
  wire [6:0]  _slots_1_io_out_uop_uopc;
  wire [31:0] _slots_1_io_out_uop_inst;
  wire [31:0] _slots_1_io_out_uop_debug_inst;
  wire        _slots_1_io_out_uop_is_rvc;
  wire [39:0] _slots_1_io_out_uop_debug_pc;
  wire [2:0]  _slots_1_io_out_uop_iq_type;
  wire [9:0]  _slots_1_io_out_uop_fu_code;
  wire [1:0]  _slots_1_io_out_uop_iw_state;
  wire        _slots_1_io_out_uop_iw_p1_poisoned;
  wire        _slots_1_io_out_uop_iw_p2_poisoned;
  wire        _slots_1_io_out_uop_is_br;
  wire        _slots_1_io_out_uop_is_jalr;
  wire        _slots_1_io_out_uop_is_jal;
  wire        _slots_1_io_out_uop_is_sfb;
  wire [19:0] _slots_1_io_out_uop_br_mask;
  wire [4:0]  _slots_1_io_out_uop_br_tag;
  wire [5:0]  _slots_1_io_out_uop_ftq_idx;
  wire        _slots_1_io_out_uop_edge_inst;
  wire [5:0]  _slots_1_io_out_uop_pc_lob;
  wire        _slots_1_io_out_uop_taken;
  wire [19:0] _slots_1_io_out_uop_imm_packed;
  wire [11:0] _slots_1_io_out_uop_csr_addr;
  wire [6:0]  _slots_1_io_out_uop_rob_idx;
  wire [4:0]  _slots_1_io_out_uop_ldq_idx;
  wire [4:0]  _slots_1_io_out_uop_stq_idx;
  wire [1:0]  _slots_1_io_out_uop_rxq_idx;
  wire [6:0]  _slots_1_io_out_uop_pdst;
  wire [6:0]  _slots_1_io_out_uop_prs1;
  wire [6:0]  _slots_1_io_out_uop_prs2;
  wire [6:0]  _slots_1_io_out_uop_prs3;
  wire [5:0]  _slots_1_io_out_uop_ppred;
  wire        _slots_1_io_out_uop_prs1_busy;
  wire        _slots_1_io_out_uop_prs2_busy;
  wire        _slots_1_io_out_uop_prs3_busy;
  wire        _slots_1_io_out_uop_ppred_busy;
  wire [6:0]  _slots_1_io_out_uop_stale_pdst;
  wire        _slots_1_io_out_uop_exception;
  wire [63:0] _slots_1_io_out_uop_exc_cause;
  wire        _slots_1_io_out_uop_bypassable;
  wire [4:0]  _slots_1_io_out_uop_mem_cmd;
  wire [1:0]  _slots_1_io_out_uop_mem_size;
  wire        _slots_1_io_out_uop_mem_signed;
  wire        _slots_1_io_out_uop_is_fence;
  wire        _slots_1_io_out_uop_is_fencei;
  wire        _slots_1_io_out_uop_is_amo;
  wire        _slots_1_io_out_uop_uses_ldq;
  wire        _slots_1_io_out_uop_uses_stq;
  wire        _slots_1_io_out_uop_is_sys_pc2epc;
  wire        _slots_1_io_out_uop_is_unique;
  wire        _slots_1_io_out_uop_flush_on_commit;
  wire        _slots_1_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_1_io_out_uop_ldst;
  wire [5:0]  _slots_1_io_out_uop_lrs1;
  wire [5:0]  _slots_1_io_out_uop_lrs2;
  wire [5:0]  _slots_1_io_out_uop_lrs3;
  wire        _slots_1_io_out_uop_ldst_val;
  wire [1:0]  _slots_1_io_out_uop_dst_rtype;
  wire [1:0]  _slots_1_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_1_io_out_uop_lrs2_rtype;
  wire        _slots_1_io_out_uop_frs3_en;
  wire        _slots_1_io_out_uop_fp_val;
  wire        _slots_1_io_out_uop_fp_single;
  wire        _slots_1_io_out_uop_xcpt_pf_if;
  wire        _slots_1_io_out_uop_xcpt_ae_if;
  wire        _slots_1_io_out_uop_xcpt_ma_if;
  wire        _slots_1_io_out_uop_bp_debug_if;
  wire        _slots_1_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_1_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_1_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_1_io_uop_uopc;
  wire [31:0] _slots_1_io_uop_inst;
  wire [31:0] _slots_1_io_uop_debug_inst;
  wire        _slots_1_io_uop_is_rvc;
  wire [39:0] _slots_1_io_uop_debug_pc;
  wire [2:0]  _slots_1_io_uop_iq_type;
  wire [9:0]  _slots_1_io_uop_fu_code;
  wire [1:0]  _slots_1_io_uop_iw_state;
  wire        _slots_1_io_uop_iw_p1_poisoned;
  wire        _slots_1_io_uop_iw_p2_poisoned;
  wire        _slots_1_io_uop_is_br;
  wire        _slots_1_io_uop_is_jalr;
  wire        _slots_1_io_uop_is_jal;
  wire        _slots_1_io_uop_is_sfb;
  wire [19:0] _slots_1_io_uop_br_mask;
  wire [4:0]  _slots_1_io_uop_br_tag;
  wire [5:0]  _slots_1_io_uop_ftq_idx;
  wire        _slots_1_io_uop_edge_inst;
  wire [5:0]  _slots_1_io_uop_pc_lob;
  wire        _slots_1_io_uop_taken;
  wire [19:0] _slots_1_io_uop_imm_packed;
  wire [11:0] _slots_1_io_uop_csr_addr;
  wire [6:0]  _slots_1_io_uop_rob_idx;
  wire [4:0]  _slots_1_io_uop_ldq_idx;
  wire [4:0]  _slots_1_io_uop_stq_idx;
  wire [1:0]  _slots_1_io_uop_rxq_idx;
  wire [6:0]  _slots_1_io_uop_pdst;
  wire [6:0]  _slots_1_io_uop_prs1;
  wire [6:0]  _slots_1_io_uop_prs2;
  wire [6:0]  _slots_1_io_uop_prs3;
  wire [5:0]  _slots_1_io_uop_ppred;
  wire        _slots_1_io_uop_prs1_busy;
  wire        _slots_1_io_uop_prs2_busy;
  wire        _slots_1_io_uop_prs3_busy;
  wire        _slots_1_io_uop_ppred_busy;
  wire [6:0]  _slots_1_io_uop_stale_pdst;
  wire        _slots_1_io_uop_exception;
  wire [63:0] _slots_1_io_uop_exc_cause;
  wire        _slots_1_io_uop_bypassable;
  wire [4:0]  _slots_1_io_uop_mem_cmd;
  wire [1:0]  _slots_1_io_uop_mem_size;
  wire        _slots_1_io_uop_mem_signed;
  wire        _slots_1_io_uop_is_fence;
  wire        _slots_1_io_uop_is_fencei;
  wire        _slots_1_io_uop_is_amo;
  wire        _slots_1_io_uop_uses_ldq;
  wire        _slots_1_io_uop_uses_stq;
  wire        _slots_1_io_uop_is_sys_pc2epc;
  wire        _slots_1_io_uop_is_unique;
  wire        _slots_1_io_uop_flush_on_commit;
  wire        _slots_1_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_1_io_uop_ldst;
  wire [5:0]  _slots_1_io_uop_lrs1;
  wire [5:0]  _slots_1_io_uop_lrs2;
  wire [5:0]  _slots_1_io_uop_lrs3;
  wire        _slots_1_io_uop_ldst_val;
  wire [1:0]  _slots_1_io_uop_dst_rtype;
  wire [1:0]  _slots_1_io_uop_lrs1_rtype;
  wire [1:0]  _slots_1_io_uop_lrs2_rtype;
  wire        _slots_1_io_uop_frs3_en;
  wire        _slots_1_io_uop_fp_val;
  wire        _slots_1_io_uop_fp_single;
  wire        _slots_1_io_uop_xcpt_pf_if;
  wire        _slots_1_io_uop_xcpt_ae_if;
  wire        _slots_1_io_uop_xcpt_ma_if;
  wire        _slots_1_io_uop_bp_debug_if;
  wire        _slots_1_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_1_io_uop_debug_fsrc;
  wire [1:0]  _slots_1_io_uop_debug_tsrc;
  wire        _slots_0_io_valid;
  wire        _slots_0_io_will_be_valid;
  wire        _slots_0_io_request;
  wire [6:0]  _slots_0_io_uop_uopc;
  wire [31:0] _slots_0_io_uop_inst;
  wire [31:0] _slots_0_io_uop_debug_inst;
  wire        _slots_0_io_uop_is_rvc;
  wire [39:0] _slots_0_io_uop_debug_pc;
  wire [2:0]  _slots_0_io_uop_iq_type;
  wire [9:0]  _slots_0_io_uop_fu_code;
  wire [1:0]  _slots_0_io_uop_iw_state;
  wire        _slots_0_io_uop_iw_p1_poisoned;
  wire        _slots_0_io_uop_iw_p2_poisoned;
  wire        _slots_0_io_uop_is_br;
  wire        _slots_0_io_uop_is_jalr;
  wire        _slots_0_io_uop_is_jal;
  wire        _slots_0_io_uop_is_sfb;
  wire [19:0] _slots_0_io_uop_br_mask;
  wire [4:0]  _slots_0_io_uop_br_tag;
  wire [5:0]  _slots_0_io_uop_ftq_idx;
  wire        _slots_0_io_uop_edge_inst;
  wire [5:0]  _slots_0_io_uop_pc_lob;
  wire        _slots_0_io_uop_taken;
  wire [19:0] _slots_0_io_uop_imm_packed;
  wire [11:0] _slots_0_io_uop_csr_addr;
  wire [6:0]  _slots_0_io_uop_rob_idx;
  wire [4:0]  _slots_0_io_uop_ldq_idx;
  wire [4:0]  _slots_0_io_uop_stq_idx;
  wire [1:0]  _slots_0_io_uop_rxq_idx;
  wire [6:0]  _slots_0_io_uop_pdst;
  wire [6:0]  _slots_0_io_uop_prs1;
  wire [6:0]  _slots_0_io_uop_prs2;
  wire [6:0]  _slots_0_io_uop_prs3;
  wire [5:0]  _slots_0_io_uop_ppred;
  wire        _slots_0_io_uop_prs1_busy;
  wire        _slots_0_io_uop_prs2_busy;
  wire        _slots_0_io_uop_prs3_busy;
  wire        _slots_0_io_uop_ppred_busy;
  wire [6:0]  _slots_0_io_uop_stale_pdst;
  wire        _slots_0_io_uop_exception;
  wire [63:0] _slots_0_io_uop_exc_cause;
  wire        _slots_0_io_uop_bypassable;
  wire [4:0]  _slots_0_io_uop_mem_cmd;
  wire [1:0]  _slots_0_io_uop_mem_size;
  wire        _slots_0_io_uop_mem_signed;
  wire        _slots_0_io_uop_is_fence;
  wire        _slots_0_io_uop_is_fencei;
  wire        _slots_0_io_uop_is_amo;
  wire        _slots_0_io_uop_uses_ldq;
  wire        _slots_0_io_uop_uses_stq;
  wire        _slots_0_io_uop_is_sys_pc2epc;
  wire        _slots_0_io_uop_is_unique;
  wire        _slots_0_io_uop_flush_on_commit;
  wire        _slots_0_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_0_io_uop_ldst;
  wire [5:0]  _slots_0_io_uop_lrs1;
  wire [5:0]  _slots_0_io_uop_lrs2;
  wire [5:0]  _slots_0_io_uop_lrs3;
  wire        _slots_0_io_uop_ldst_val;
  wire [1:0]  _slots_0_io_uop_dst_rtype;
  wire [1:0]  _slots_0_io_uop_lrs1_rtype;
  wire [1:0]  _slots_0_io_uop_lrs2_rtype;
  wire        _slots_0_io_uop_frs3_en;
  wire        _slots_0_io_uop_fp_val;
  wire        _slots_0_io_uop_fp_single;
  wire        _slots_0_io_uop_xcpt_pf_if;
  wire        _slots_0_io_uop_xcpt_ae_if;
  wire        _slots_0_io_uop_xcpt_ma_if;
  wire        _slots_0_io_uop_bp_debug_if;
  wire        _slots_0_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_0_io_uop_debug_fsrc;
  wire [1:0]  _slots_0_io_uop_debug_tsrc;
  wire        _GEN = io_dis_uops_0_bits_uopc == 7'h2;
  wire        _GEN_0 = _GEN & ~(|io_dis_uops_0_bits_lrs2_rtype) | io_dis_uops_0_bits_uopc == 7'h43;
  wire [1:0]  _GEN_1 = _GEN_0 ? 2'h2 : 2'h1;
  wire        _GEN_2 = _GEN_0 | ~(_GEN & (|io_dis_uops_0_bits_lrs2_rtype));
  wire [1:0]  _GEN_3 = _GEN_2 ? io_dis_uops_0_bits_lrs2_rtype : 2'h2;
  wire        _GEN_4 = _GEN_2 & io_dis_uops_0_bits_prs2_busy;
  wire        _GEN_5 = io_dis_uops_1_bits_uopc == 7'h2;
  wire        _GEN_6 = _GEN_5 & ~(|io_dis_uops_1_bits_lrs2_rtype) | io_dis_uops_1_bits_uopc == 7'h43;
  wire [1:0]  _GEN_7 = _GEN_6 ? 2'h2 : 2'h1;
  wire        _GEN_8 = _GEN_6 | ~(_GEN_5 & (|io_dis_uops_1_bits_lrs2_rtype));
  wire [1:0]  _GEN_9 = _GEN_8 ? io_dis_uops_1_bits_lrs2_rtype : 2'h2;
  wire        _GEN_10 = _GEN_8 & io_dis_uops_1_bits_prs2_busy;
  wire        _GEN_11 = io_dis_uops_2_bits_uopc == 7'h2;
  wire        _GEN_12 = _GEN_11 & ~(|io_dis_uops_2_bits_lrs2_rtype) | io_dis_uops_2_bits_uopc == 7'h43;
  wire        _GEN_13 = _GEN_12 | ~(_GEN_11 & (|io_dis_uops_2_bits_lrs2_rtype));
  wire [1:0]  _GEN_14 = _GEN_13 ? io_dis_uops_2_bits_lrs2_rtype : 2'h2;
  wire        _GEN_15 = _GEN_13 & io_dis_uops_2_bits_prs2_busy;
  wire        _GEN_16 = io_dis_uops_3_bits_uopc == 7'h2;
  wire        _GEN_17 = _GEN_16 & ~(|io_dis_uops_3_bits_lrs2_rtype) | io_dis_uops_3_bits_uopc == 7'h43;
  wire        _GEN_18 = _GEN_17 | ~(_GEN_16 & (|io_dis_uops_3_bits_lrs2_rtype));
  wire [4:0]  count = {1'h0, {1'h0, {1'h0, {1'h0, _slots_0_io_valid} + {1'h0, _slots_1_io_valid} + {1'h0, _slots_2_io_valid}} + {1'h0, {1'h0, _slots_3_io_valid} + {1'h0, _slots_4_io_valid} + {1'h0, _slots_5_io_valid}}} + {1'h0, {1'h0, {1'h0, _slots_6_io_valid} + {1'h0, _slots_7_io_valid} + {1'h0, _slots_8_io_valid}} + {1'h0, {1'h0, _slots_9_io_valid} + {1'h0, _slots_10_io_valid} + {1'h0, _slots_11_io_valid}}}} + {1'h0, {1'h0, {1'h0, {1'h0, _slots_12_io_valid} + {1'h0, _slots_13_io_valid} + {1'h0, _slots_14_io_valid}} + {1'h0, {1'h0, _slots_15_io_valid} + {1'h0, _slots_16_io_valid} + {1'h0, _slots_17_io_valid}}} + {1'h0, {1'h0, {1'h0, _slots_18_io_valid} + {1'h0, _slots_19_io_valid} + {1'h0, _slots_20_io_valid}} + {1'h0, {1'h0, _slots_21_io_valid} + {1'h0, _slots_22_io_valid} + {1'h0, _slots_23_io_valid}}}};
  `ifndef SYNTHESIS
    always @(posedge clock) begin
      if (~reset & {1'h0, {1'h0, {1'h0, {1'h0, issue_slots_0_grant} + {1'h0, issue_slots_1_grant} + {1'h0, issue_slots_2_grant}} + {1'h0, {1'h0, issue_slots_3_grant} + {1'h0, issue_slots_4_grant} + {1'h0, issue_slots_5_grant}}} + {1'h0, {1'h0, {1'h0, issue_slots_6_grant} + {1'h0, issue_slots_7_grant} + {1'h0, issue_slots_8_grant}} + {1'h0, {1'h0, issue_slots_9_grant} + {1'h0, issue_slots_10_grant} + {1'h0, issue_slots_11_grant}}}} + {1'h0, {1'h0, {1'h0, {1'h0, issue_slots_12_grant} + {1'h0, issue_slots_13_grant} + {1'h0, issue_slots_14_grant}} + {1'h0, {1'h0, issue_slots_15_grant} + {1'h0, issue_slots_16_grant} + {1'h0, issue_slots_17_grant}}} + {1'h0, {1'h0, {1'h0, issue_slots_18_grant} + {1'h0, issue_slots_19_grant} + {1'h0, issue_slots_20_grant}} + {1'h0, {1'h0, issue_slots_21_grant} + {1'h0, issue_slots_22_grant} + {1'h0, issue_slots_23_grant}}}} > 5'h2) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [issue] window giving out too many grants.\n    at issue-unit.scala:172 assert (PopCount(issue_slots.map(s => s.grant)) <= issueWidth.U, \"[issue] window giving out too many grants.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire [3:0]  next_1 = _slots_0_io_valid & ~_slots_1_io_valid ? 4'h1 : _slots_1_io_valid ? {3'h0, ~_slots_0_io_valid} : {2'h0, ~_slots_0_io_valid, 1'h0};
  assign _next_1_1to0 = next_1[1:0];
  assign next_2 = _next_1_1to0 == 2'h0 & ~_slots_2_io_valid ? 4'h1 : next_1[3] | _slots_2_io_valid ? next_1 : {next_1[2:0], 1'h0};
  assign next_3 = next_2 == 4'h0 & ~_slots_3_io_valid ? 4'h1 : next_2[3] | _slots_3_io_valid ? next_2 : {next_2[2:0], 1'h0};
  assign next_4 = next_3 == 4'h0 & ~_slots_4_io_valid ? 4'h1 : next_3[3] | _slots_4_io_valid ? next_3 : {next_3[2:0], 1'h0};
  assign next_5 = next_4 == 4'h0 & ~_slots_5_io_valid ? 4'h1 : next_4[3] | _slots_5_io_valid ? next_4 : {next_4[2:0], 1'h0};
  assign next_6 = next_5 == 4'h0 & ~_slots_6_io_valid ? 4'h1 : next_5[3] | _slots_6_io_valid ? next_5 : {next_5[2:0], 1'h0};
  assign next_7 = next_6 == 4'h0 & ~_slots_7_io_valid ? 4'h1 : next_6[3] | _slots_7_io_valid ? next_6 : {next_6[2:0], 1'h0};
  assign next_8 = next_7 == 4'h0 & ~_slots_8_io_valid ? 4'h1 : next_7[3] | _slots_8_io_valid ? next_7 : {next_7[2:0], 1'h0};
  assign next_9 = next_8 == 4'h0 & ~_slots_9_io_valid ? 4'h1 : next_8[3] | _slots_9_io_valid ? next_8 : {next_8[2:0], 1'h0};
  assign next_10 = next_9 == 4'h0 & ~_slots_10_io_valid ? 4'h1 : next_9[3] | _slots_10_io_valid ? next_9 : {next_9[2:0], 1'h0};
  assign next_11 = next_10 == 4'h0 & ~_slots_11_io_valid ? 4'h1 : next_10[3] | _slots_11_io_valid ? next_10 : {next_10[2:0], 1'h0};
  assign next_12 = next_11 == 4'h0 & ~_slots_12_io_valid ? 4'h1 : next_11[3] | _slots_12_io_valid ? next_11 : {next_11[2:0], 1'h0};
  assign next_13 = next_12 == 4'h0 & ~_slots_13_io_valid ? 4'h1 : next_12[3] | _slots_13_io_valid ? next_12 : {next_12[2:0], 1'h0};
  assign next_14 = next_13 == 4'h0 & ~_slots_14_io_valid ? 4'h1 : next_13[3] | _slots_14_io_valid ? next_13 : {next_13[2:0], 1'h0};
  assign next_15 = next_14 == 4'h0 & ~_slots_15_io_valid ? 4'h1 : next_14[3] | _slots_15_io_valid ? next_14 : {next_14[2:0], 1'h0};
  assign next_16 = next_15 == 4'h0 & ~_slots_16_io_valid ? 4'h1 : next_15[3] | _slots_16_io_valid ? next_15 : {next_15[2:0], 1'h0};
  assign next_17 = next_16 == 4'h0 & ~_slots_17_io_valid ? 4'h1 : next_16[3] | _slots_17_io_valid ? next_16 : {next_16[2:0], 1'h0};
  assign next_18 = next_17 == 4'h0 & ~_slots_18_io_valid ? 4'h1 : next_17[3] | _slots_18_io_valid ? next_17 : {next_17[2:0], 1'h0};
  assign next_19 = next_18 == 4'h0 & ~_slots_19_io_valid ? 4'h1 : next_18[3] | _slots_19_io_valid ? next_18 : {next_18[2:0], 1'h0};
  assign next_20 = next_19 == 4'h0 & ~_slots_20_io_valid ? 4'h1 : next_19[3] | _slots_20_io_valid ? next_19 : {next_19[2:0], 1'h0};
  assign next_21 = next_20 == 4'h0 & ~_slots_21_io_valid ? 4'h1 : next_20[3] | _slots_21_io_valid ? next_20 : {next_20[2:0], 1'h0};
  assign next_22 = next_21 == 4'h0 & ~_slots_22_io_valid ? 4'h1 : next_21[3] | _slots_22_io_valid ? next_21 : {next_21[2:0], 1'h0};
  wire [3:0]  next_23 = next_22 == 4'h0 & ~_slots_23_io_valid ? 4'h1 : next_22[3] | _slots_23_io_valid ? next_22 : {next_22[2:0], 1'h0};
  wire [3:0]  next_24 = next_23 == 4'h0 & ~io_dis_uops_0_valid ? 4'h1 : next_23[3] | io_dis_uops_0_valid ? next_23 : {next_23[2:0], 1'h0};
  wire [3:0]  next_25 = next_24 == 4'h0 & ~io_dis_uops_1_valid ? 4'h1 : next_24[3] | io_dis_uops_1_valid ? next_24 : {next_24[2:0], 1'h0};
  wire        will_be_valid_24 = io_dis_uops_0_valid & ~io_dis_uops_0_bits_exception & ~io_dis_uops_0_bits_is_fence & ~io_dis_uops_0_bits_is_fencei;
  wire        will_be_valid_25 = io_dis_uops_1_valid & ~io_dis_uops_1_bits_exception & ~io_dis_uops_1_bits_is_fence & ~io_dis_uops_1_bits_is_fencei;
  wire        will_be_valid_26 = io_dis_uops_2_valid & ~io_dis_uops_2_bits_exception & ~io_dis_uops_2_bits_is_fence & ~io_dis_uops_2_bits_is_fencei;
  wire        _GEN_19 = _next_1_1to0 == 2'h2;
  wire        _GEN_20 = next_2 == 4'h4;
  wire        _GEN_21 = next_3 == 4'h8;
  wire        issue_slots_0_in_uop_valid = _GEN_21 ? _slots_4_io_will_be_valid : _GEN_20 ? _slots_3_io_will_be_valid : _GEN_19 ? _slots_2_io_will_be_valid : ~_slots_0_io_valid & _slots_1_io_will_be_valid;
  wire        _GEN_22 = next_2 == 4'h2;
  wire        _GEN_23 = next_3 == 4'h4;
  wire        _GEN_24 = next_4 == 4'h8;
  wire        issue_slots_1_in_uop_valid = _GEN_24 ? _slots_5_io_will_be_valid : _GEN_23 ? _slots_4_io_will_be_valid : _GEN_22 ? _slots_3_io_will_be_valid : _next_1_1to0 == 2'h1 & _slots_2_io_will_be_valid;
  wire        _GEN_25 = next_3 == 4'h2;
  wire        _GEN_26 = next_4 == 4'h4;
  wire        _GEN_27 = next_5 == 4'h8;
  wire        issue_slots_2_in_uop_valid = _GEN_27 ? _slots_6_io_will_be_valid : _GEN_26 ? _slots_5_io_will_be_valid : _GEN_25 ? _slots_4_io_will_be_valid : next_2 == 4'h1 & _slots_3_io_will_be_valid;
  wire        _GEN_28 = next_4 == 4'h2;
  wire        _GEN_29 = next_5 == 4'h4;
  wire        _GEN_30 = next_6 == 4'h8;
  wire        issue_slots_3_in_uop_valid = _GEN_30 ? _slots_7_io_will_be_valid : _GEN_29 ? _slots_6_io_will_be_valid : _GEN_28 ? _slots_5_io_will_be_valid : next_3 == 4'h1 & _slots_4_io_will_be_valid;
  wire        _GEN_31 = next_5 == 4'h2;
  wire        _GEN_32 = next_6 == 4'h4;
  wire        _GEN_33 = next_7 == 4'h8;
  wire        issue_slots_4_in_uop_valid = _GEN_33 ? _slots_8_io_will_be_valid : _GEN_32 ? _slots_7_io_will_be_valid : _GEN_31 ? _slots_6_io_will_be_valid : next_4 == 4'h1 & _slots_5_io_will_be_valid;
  wire        _GEN_34 = next_6 == 4'h2;
  wire        _GEN_35 = next_7 == 4'h4;
  wire        _GEN_36 = next_8 == 4'h8;
  wire        issue_slots_5_in_uop_valid = _GEN_36 ? _slots_9_io_will_be_valid : _GEN_35 ? _slots_8_io_will_be_valid : _GEN_34 ? _slots_7_io_will_be_valid : next_5 == 4'h1 & _slots_6_io_will_be_valid;
  wire        _GEN_37 = next_7 == 4'h2;
  wire        _GEN_38 = next_8 == 4'h4;
  wire        _GEN_39 = next_9 == 4'h8;
  wire        issue_slots_6_in_uop_valid = _GEN_39 ? _slots_10_io_will_be_valid : _GEN_38 ? _slots_9_io_will_be_valid : _GEN_37 ? _slots_8_io_will_be_valid : next_6 == 4'h1 & _slots_7_io_will_be_valid;
  wire        _GEN_40 = next_8 == 4'h2;
  wire        _GEN_41 = next_9 == 4'h4;
  wire        _GEN_42 = next_10 == 4'h8;
  wire        issue_slots_7_in_uop_valid = _GEN_42 ? _slots_11_io_will_be_valid : _GEN_41 ? _slots_10_io_will_be_valid : _GEN_40 ? _slots_9_io_will_be_valid : next_7 == 4'h1 & _slots_8_io_will_be_valid;
  wire        _GEN_43 = next_9 == 4'h2;
  wire        _GEN_44 = next_10 == 4'h4;
  wire        _GEN_45 = next_11 == 4'h8;
  wire        issue_slots_8_in_uop_valid = _GEN_45 ? _slots_12_io_will_be_valid : _GEN_44 ? _slots_11_io_will_be_valid : _GEN_43 ? _slots_10_io_will_be_valid : next_8 == 4'h1 & _slots_9_io_will_be_valid;
  wire        _GEN_46 = next_10 == 4'h2;
  wire        _GEN_47 = next_11 == 4'h4;
  wire        _GEN_48 = next_12 == 4'h8;
  wire        issue_slots_9_in_uop_valid = _GEN_48 ? _slots_13_io_will_be_valid : _GEN_47 ? _slots_12_io_will_be_valid : _GEN_46 ? _slots_11_io_will_be_valid : next_9 == 4'h1 & _slots_10_io_will_be_valid;
  wire        _GEN_49 = next_11 == 4'h2;
  wire        _GEN_50 = next_12 == 4'h4;
  wire        _GEN_51 = next_13 == 4'h8;
  wire        issue_slots_10_in_uop_valid = _GEN_51 ? _slots_14_io_will_be_valid : _GEN_50 ? _slots_13_io_will_be_valid : _GEN_49 ? _slots_12_io_will_be_valid : next_10 == 4'h1 & _slots_11_io_will_be_valid;
  wire        _GEN_52 = next_12 == 4'h2;
  wire        _GEN_53 = next_13 == 4'h4;
  wire        _GEN_54 = next_14 == 4'h8;
  wire        issue_slots_11_in_uop_valid = _GEN_54 ? _slots_15_io_will_be_valid : _GEN_53 ? _slots_14_io_will_be_valid : _GEN_52 ? _slots_13_io_will_be_valid : next_11 == 4'h1 & _slots_12_io_will_be_valid;
  wire        _GEN_55 = next_13 == 4'h2;
  wire        _GEN_56 = next_14 == 4'h4;
  wire        _GEN_57 = next_15 == 4'h8;
  wire        issue_slots_12_in_uop_valid = _GEN_57 ? _slots_16_io_will_be_valid : _GEN_56 ? _slots_15_io_will_be_valid : _GEN_55 ? _slots_14_io_will_be_valid : next_12 == 4'h1 & _slots_13_io_will_be_valid;
  wire        _GEN_58 = next_14 == 4'h2;
  wire        _GEN_59 = next_15 == 4'h4;
  wire        _GEN_60 = next_16 == 4'h8;
  wire        issue_slots_13_in_uop_valid = _GEN_60 ? _slots_17_io_will_be_valid : _GEN_59 ? _slots_16_io_will_be_valid : _GEN_58 ? _slots_15_io_will_be_valid : next_13 == 4'h1 & _slots_14_io_will_be_valid;
  wire        _GEN_61 = next_15 == 4'h2;
  wire        _GEN_62 = next_16 == 4'h4;
  wire        _GEN_63 = next_17 == 4'h8;
  wire        issue_slots_14_in_uop_valid = _GEN_63 ? _slots_18_io_will_be_valid : _GEN_62 ? _slots_17_io_will_be_valid : _GEN_61 ? _slots_16_io_will_be_valid : next_14 == 4'h1 & _slots_15_io_will_be_valid;
  wire        _GEN_64 = next_16 == 4'h2;
  wire        _GEN_65 = next_17 == 4'h4;
  wire        _GEN_66 = next_18 == 4'h8;
  wire        issue_slots_15_in_uop_valid = _GEN_66 ? _slots_19_io_will_be_valid : _GEN_65 ? _slots_18_io_will_be_valid : _GEN_64 ? _slots_17_io_will_be_valid : next_15 == 4'h1 & _slots_16_io_will_be_valid;
  wire        _GEN_67 = next_17 == 4'h2;
  wire        _GEN_68 = next_18 == 4'h4;
  wire        _GEN_69 = next_19 == 4'h8;
  wire        issue_slots_16_in_uop_valid = _GEN_69 ? _slots_20_io_will_be_valid : _GEN_68 ? _slots_19_io_will_be_valid : _GEN_67 ? _slots_18_io_will_be_valid : next_16 == 4'h1 & _slots_17_io_will_be_valid;
  wire        _GEN_70 = next_18 == 4'h2;
  wire        _GEN_71 = next_19 == 4'h4;
  wire        _GEN_72 = next_20 == 4'h8;
  wire        issue_slots_17_in_uop_valid = _GEN_72 ? _slots_21_io_will_be_valid : _GEN_71 ? _slots_20_io_will_be_valid : _GEN_70 ? _slots_19_io_will_be_valid : next_17 == 4'h1 & _slots_18_io_will_be_valid;
  wire        _GEN_73 = next_19 == 4'h2;
  wire        _GEN_74 = next_20 == 4'h4;
  wire        _GEN_75 = next_21 == 4'h8;
  wire        issue_slots_18_in_uop_valid = _GEN_75 ? _slots_22_io_will_be_valid : _GEN_74 ? _slots_21_io_will_be_valid : _GEN_73 ? _slots_20_io_will_be_valid : next_18 == 4'h1 & _slots_19_io_will_be_valid;
  wire        _GEN_76 = next_20 == 4'h2;
  wire        _GEN_77 = next_21 == 4'h4;
  wire        _GEN_78 = next_22 == 4'h8;
  wire        issue_slots_19_in_uop_valid = _GEN_78 ? _slots_23_io_will_be_valid : _GEN_77 ? _slots_22_io_will_be_valid : _GEN_76 ? _slots_21_io_will_be_valid : next_19 == 4'h1 & _slots_20_io_will_be_valid;
  wire        _GEN_79 = next_21 == 4'h2;
  wire        _GEN_80 = next_22 == 4'h4;
  wire        _GEN_81 = next_23 == 4'h8;
  wire        issue_slots_20_in_uop_valid = _GEN_81 ? will_be_valid_24 : _GEN_80 ? _slots_23_io_will_be_valid : _GEN_79 ? _slots_22_io_will_be_valid : next_20 == 4'h1 & _slots_21_io_will_be_valid;
  wire        _GEN_82 = next_22 == 4'h2;
  wire        _GEN_83 = next_23 == 4'h4;
  wire        _GEN_84 = next_24 == 4'h8;
  wire        issue_slots_21_in_uop_valid = _GEN_84 ? will_be_valid_25 : _GEN_83 ? will_be_valid_24 : _GEN_82 ? _slots_23_io_will_be_valid : next_21 == 4'h1 & _slots_22_io_will_be_valid;
  wire        _GEN_85 = _GEN_84 | _GEN_83;
  wire        _GEN_86 = next_23 == 4'h2;
  wire        _GEN_87 = next_24 == 4'h4;
  wire        _GEN_88 = next_25 == 4'h8;
  wire        issue_slots_22_in_uop_valid = _GEN_88 ? will_be_valid_26 : _GEN_87 ? will_be_valid_25 : _GEN_86 ? will_be_valid_24 : next_22 == 4'h1 & _slots_23_io_will_be_valid;
  wire        _GEN_89 = _GEN_88 | _GEN_87 | _GEN_86;
  wire        _GEN_90 = next_24 == 4'h2;
  wire        _GEN_91 = next_25 == 4'h4;
  wire        _GEN_92 = (next_25 == 4'h0 & ~io_dis_uops_2_valid ? 4'h1 : next_25[3] | io_dis_uops_2_valid ? next_25 : {next_25[2:0], 1'h0}) == 4'h8;
  wire        issue_slots_23_in_uop_valid = _GEN_92 ? io_dis_uops_3_valid & ~io_dis_uops_3_bits_exception & ~io_dis_uops_3_bits_is_fence & ~io_dis_uops_3_bits_is_fencei : _GEN_91 ? will_be_valid_26 : _GEN_90 ? will_be_valid_25 : next_23 == 4'h1 & will_be_valid_24;
  reg         io_dis_uops_0_ready_REG;
  reg         io_dis_uops_1_ready_REG;
  reg         io_dis_uops_2_ready_REG;
  reg         io_dis_uops_3_ready_REG;
  wire        _GEN_93 = _slots_0_io_request & (|(_slots_0_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_94 = _slots_0_io_request & ~_GEN_93 & (|(_slots_0_io_uop_fu_code & io_fu_types_1));
  assign issue_slots_0_grant = _GEN_94 | _GEN_93;
  wire        _GEN_95 = _slots_1_io_request & (|(_slots_1_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_96 = _GEN_95 & ~_GEN_93;
  wire        _GEN_97 = _GEN_95 | _GEN_93;
  wire        _GEN_98 = _slots_1_io_request & ~_GEN_96 & (|(_slots_1_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_99 = _GEN_98 & ~_GEN_94;
  assign issue_slots_1_grant = _GEN_99 | _GEN_96;
  wire        _GEN_100 = _GEN_98 | _GEN_94;
  wire        _GEN_101 = _slots_2_io_request & (|(_slots_2_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_102 = _GEN_101 & ~_GEN_97;
  wire        _GEN_103 = _GEN_101 | _GEN_97;
  wire        _GEN_104 = _slots_2_io_request & ~_GEN_102 & (|(_slots_2_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_105 = _GEN_104 & ~_GEN_100;
  assign issue_slots_2_grant = _GEN_105 | _GEN_102;
  wire        _GEN_106 = _GEN_104 | _GEN_100;
  wire        _GEN_107 = _slots_3_io_request & (|(_slots_3_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_108 = _GEN_107 & ~_GEN_103;
  wire        _GEN_109 = _GEN_107 | _GEN_103;
  wire        _GEN_110 = _slots_3_io_request & ~_GEN_108 & (|(_slots_3_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_111 = _GEN_110 & ~_GEN_106;
  assign issue_slots_3_grant = _GEN_111 | _GEN_108;
  wire        _GEN_112 = _GEN_110 | _GEN_106;
  wire        _GEN_113 = _slots_4_io_request & (|(_slots_4_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_114 = _GEN_113 & ~_GEN_109;
  wire        _GEN_115 = _GEN_113 | _GEN_109;
  wire        _GEN_116 = _slots_4_io_request & ~_GEN_114 & (|(_slots_4_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_117 = _GEN_116 & ~_GEN_112;
  assign issue_slots_4_grant = _GEN_117 | _GEN_114;
  wire        _GEN_118 = _GEN_116 | _GEN_112;
  wire        _GEN_119 = _slots_5_io_request & (|(_slots_5_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_120 = _GEN_119 & ~_GEN_115;
  wire        _GEN_121 = _GEN_119 | _GEN_115;
  wire        _GEN_122 = _slots_5_io_request & ~_GEN_120 & (|(_slots_5_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_123 = _GEN_122 & ~_GEN_118;
  assign issue_slots_5_grant = _GEN_123 | _GEN_120;
  wire        _GEN_124 = _GEN_122 | _GEN_118;
  wire        _GEN_125 = _slots_6_io_request & (|(_slots_6_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_126 = _GEN_125 & ~_GEN_121;
  wire        _GEN_127 = _GEN_125 | _GEN_121;
  wire        _GEN_128 = _slots_6_io_request & ~_GEN_126 & (|(_slots_6_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_129 = _GEN_128 & ~_GEN_124;
  assign issue_slots_6_grant = _GEN_129 | _GEN_126;
  wire        _GEN_130 = _GEN_128 | _GEN_124;
  wire        _GEN_131 = _slots_7_io_request & (|(_slots_7_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_132 = _GEN_131 & ~_GEN_127;
  wire        _GEN_133 = _GEN_131 | _GEN_127;
  wire        _GEN_134 = _slots_7_io_request & ~_GEN_132 & (|(_slots_7_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_135 = _GEN_134 & ~_GEN_130;
  assign issue_slots_7_grant = _GEN_135 | _GEN_132;
  wire        _GEN_136 = _GEN_134 | _GEN_130;
  wire        _GEN_137 = _slots_8_io_request & (|(_slots_8_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_138 = _GEN_137 & ~_GEN_133;
  wire        _GEN_139 = _GEN_137 | _GEN_133;
  wire        _GEN_140 = _slots_8_io_request & ~_GEN_138 & (|(_slots_8_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_141 = _GEN_140 & ~_GEN_136;
  assign issue_slots_8_grant = _GEN_141 | _GEN_138;
  wire        _GEN_142 = _GEN_140 | _GEN_136;
  wire        _GEN_143 = _slots_9_io_request & (|(_slots_9_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_144 = _GEN_143 & ~_GEN_139;
  wire        _GEN_145 = _GEN_143 | _GEN_139;
  wire        _GEN_146 = _slots_9_io_request & ~_GEN_144 & (|(_slots_9_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_147 = _GEN_146 & ~_GEN_142;
  assign issue_slots_9_grant = _GEN_147 | _GEN_144;
  wire        _GEN_148 = _GEN_146 | _GEN_142;
  wire        _GEN_149 = _slots_10_io_request & (|(_slots_10_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_150 = _GEN_149 & ~_GEN_145;
  wire        _GEN_151 = _GEN_149 | _GEN_145;
  wire        _GEN_152 = _slots_10_io_request & ~_GEN_150 & (|(_slots_10_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_153 = _GEN_152 & ~_GEN_148;
  assign issue_slots_10_grant = _GEN_153 | _GEN_150;
  wire        _GEN_154 = _GEN_152 | _GEN_148;
  wire        _GEN_155 = _slots_11_io_request & (|(_slots_11_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_156 = _GEN_155 & ~_GEN_151;
  wire        _GEN_157 = _GEN_155 | _GEN_151;
  wire        _GEN_158 = _slots_11_io_request & ~_GEN_156 & (|(_slots_11_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_159 = _GEN_158 & ~_GEN_154;
  assign issue_slots_11_grant = _GEN_159 | _GEN_156;
  wire        _GEN_160 = _GEN_158 | _GEN_154;
  wire        _GEN_161 = _slots_12_io_request & (|(_slots_12_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_162 = _GEN_161 & ~_GEN_157;
  wire        _GEN_163 = _GEN_161 | _GEN_157;
  wire        _GEN_164 = _slots_12_io_request & ~_GEN_162 & (|(_slots_12_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_165 = _GEN_164 & ~_GEN_160;
  assign issue_slots_12_grant = _GEN_165 | _GEN_162;
  wire        _GEN_166 = _GEN_164 | _GEN_160;
  wire        _GEN_167 = _slots_13_io_request & (|(_slots_13_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_168 = _GEN_167 & ~_GEN_163;
  wire        _GEN_169 = _GEN_167 | _GEN_163;
  wire        _GEN_170 = _slots_13_io_request & ~_GEN_168 & (|(_slots_13_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_171 = _GEN_170 & ~_GEN_166;
  assign issue_slots_13_grant = _GEN_171 | _GEN_168;
  wire        _GEN_172 = _GEN_170 | _GEN_166;
  wire        _GEN_173 = _slots_14_io_request & (|(_slots_14_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_174 = _GEN_173 & ~_GEN_169;
  wire        _GEN_175 = _GEN_173 | _GEN_169;
  wire        _GEN_176 = _slots_14_io_request & ~_GEN_174 & (|(_slots_14_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_177 = _GEN_176 & ~_GEN_172;
  assign issue_slots_14_grant = _GEN_177 | _GEN_174;
  wire        _GEN_178 = _GEN_176 | _GEN_172;
  wire        _GEN_179 = _slots_15_io_request & (|(_slots_15_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_180 = _GEN_179 & ~_GEN_175;
  wire        _GEN_181 = _GEN_179 | _GEN_175;
  wire        _GEN_182 = _slots_15_io_request & ~_GEN_180 & (|(_slots_15_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_183 = _GEN_182 & ~_GEN_178;
  assign issue_slots_15_grant = _GEN_183 | _GEN_180;
  wire        _GEN_184 = _GEN_182 | _GEN_178;
  wire        _GEN_185 = _slots_16_io_request & (|(_slots_16_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_186 = _GEN_185 & ~_GEN_181;
  wire        _GEN_187 = _GEN_185 | _GEN_181;
  wire        _GEN_188 = _slots_16_io_request & ~_GEN_186 & (|(_slots_16_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_189 = _GEN_188 & ~_GEN_184;
  assign issue_slots_16_grant = _GEN_189 | _GEN_186;
  wire        _GEN_190 = _GEN_188 | _GEN_184;
  wire        _GEN_191 = _slots_17_io_request & (|(_slots_17_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_192 = _GEN_191 & ~_GEN_187;
  wire        _GEN_193 = _GEN_191 | _GEN_187;
  wire        _GEN_194 = _slots_17_io_request & ~_GEN_192 & (|(_slots_17_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_195 = _GEN_194 & ~_GEN_190;
  assign issue_slots_17_grant = _GEN_195 | _GEN_192;
  wire        _GEN_196 = _GEN_194 | _GEN_190;
  wire        _GEN_197 = _slots_18_io_request & (|(_slots_18_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_198 = _GEN_197 & ~_GEN_193;
  wire        _GEN_199 = _GEN_197 | _GEN_193;
  wire        _GEN_200 = _slots_18_io_request & ~_GEN_198 & (|(_slots_18_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_201 = _GEN_200 & ~_GEN_196;
  assign issue_slots_18_grant = _GEN_201 | _GEN_198;
  wire        _GEN_202 = _GEN_200 | _GEN_196;
  wire        _GEN_203 = _slots_19_io_request & (|(_slots_19_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_204 = _GEN_203 & ~_GEN_199;
  wire        _GEN_205 = _GEN_203 | _GEN_199;
  wire        _GEN_206 = _slots_19_io_request & ~_GEN_204 & (|(_slots_19_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_207 = _GEN_206 & ~_GEN_202;
  assign issue_slots_19_grant = _GEN_207 | _GEN_204;
  wire        _GEN_208 = _GEN_206 | _GEN_202;
  wire        _GEN_209 = _slots_20_io_request & (|(_slots_20_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_210 = _GEN_209 & ~_GEN_205;
  wire        _GEN_211 = _GEN_209 | _GEN_205;
  wire        _GEN_212 = _slots_20_io_request & ~_GEN_210 & (|(_slots_20_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_213 = _GEN_212 & ~_GEN_208;
  assign issue_slots_20_grant = _GEN_213 | _GEN_210;
  wire        _GEN_214 = _GEN_212 | _GEN_208;
  wire        _GEN_215 = _slots_21_io_request & (|(_slots_21_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_216 = _GEN_215 & ~_GEN_211;
  wire        _GEN_217 = _GEN_215 | _GEN_211;
  wire        _GEN_218 = _slots_21_io_request & ~_GEN_216 & (|(_slots_21_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_219 = _GEN_218 & ~_GEN_214;
  assign issue_slots_21_grant = _GEN_219 | _GEN_216;
  wire        _GEN_220 = _GEN_218 | _GEN_214;
  wire        _GEN_221 = _slots_22_io_request & (|(_slots_22_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_222 = _GEN_221 & ~_GEN_217;
  wire        _GEN_223 = _slots_22_io_request & ~_GEN_222 & (|(_slots_22_io_uop_fu_code & io_fu_types_1));
  wire        _GEN_224 = _GEN_223 & ~_GEN_220;
  assign issue_slots_22_grant = _GEN_224 | _GEN_222;
  wire        _GEN_225 = _slots_23_io_request & (|(_slots_23_io_uop_fu_code & io_fu_types_0)) & ~(_GEN_221 | _GEN_217);
  wire        _GEN_226 = _slots_23_io_request & ~_GEN_225 & (|(_slots_23_io_uop_fu_code & io_fu_types_1)) & ~(_GEN_223 | _GEN_220);
  assign issue_slots_23_grant = _GEN_226 | _GEN_225;
  wire [4:0]  num_available =
    {1'h0, {1'h0, {1'h0, {1'h0, ~_slots_0_io_will_be_valid & ~issue_slots_0_in_uop_valid} + {1'h0, (~_slots_1_io_will_be_valid | ~_slots_0_io_valid) & ~issue_slots_1_in_uop_valid} + {1'h0, (~_slots_2_io_will_be_valid | (|_next_1_1to0)) & ~issue_slots_2_in_uop_valid}} + {1'h0, {1'h0, (~_slots_3_io_will_be_valid | (|next_2)) & ~issue_slots_3_in_uop_valid} + {1'h0, (~_slots_4_io_will_be_valid | (|next_3)) & ~issue_slots_4_in_uop_valid} + {1'h0, (~_slots_5_io_will_be_valid | (|next_4)) & ~issue_slots_5_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_6_io_will_be_valid | (|next_5)) & ~issue_slots_6_in_uop_valid} + {1'h0, (~_slots_7_io_will_be_valid | (|next_6)) & ~issue_slots_7_in_uop_valid} + {1'h0, (~_slots_8_io_will_be_valid | (|next_7)) & ~issue_slots_8_in_uop_valid}} + {1'h0, {1'h0, (~_slots_9_io_will_be_valid | (|next_8)) & ~issue_slots_9_in_uop_valid} + {1'h0, (~_slots_10_io_will_be_valid | (|next_9)) & ~issue_slots_10_in_uop_valid} + {1'h0, (~_slots_11_io_will_be_valid | (|next_10)) & ~issue_slots_11_in_uop_valid}}}}
    + {1'h0, {1'h0, {1'h0, {1'h0, (~_slots_12_io_will_be_valid | (|next_11)) & ~issue_slots_12_in_uop_valid} + {1'h0, (~_slots_13_io_will_be_valid | (|next_12)) & ~issue_slots_13_in_uop_valid} + {1'h0, (~_slots_14_io_will_be_valid | (|next_13)) & ~issue_slots_14_in_uop_valid}} + {1'h0, {1'h0, (~_slots_15_io_will_be_valid | (|next_14)) & ~issue_slots_15_in_uop_valid} + {1'h0, (~_slots_16_io_will_be_valid | (|next_15)) & ~issue_slots_16_in_uop_valid} + {1'h0, (~_slots_17_io_will_be_valid | (|next_16)) & ~issue_slots_17_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_18_io_will_be_valid | (|next_17)) & ~issue_slots_18_in_uop_valid} + {1'h0, (~_slots_19_io_will_be_valid | (|next_18)) & ~issue_slots_19_in_uop_valid} + {1'h0, (~_slots_20_io_will_be_valid | (|next_19)) & ~issue_slots_20_in_uop_valid}} + {1'h0, {1'h0, (~_slots_21_io_will_be_valid | (|next_20)) & ~issue_slots_21_in_uop_valid} + {1'h0, (~_slots_22_io_will_be_valid | (|next_21)) & ~issue_slots_22_in_uop_valid} + {1'h0, (~_slots_23_io_will_be_valid | (|next_22)) & ~issue_slots_23_in_uop_valid}}}};
  always @(posedge clock) begin
    io_dis_uops_0_ready_REG <= |num_available;
    io_dis_uops_1_ready_REG <= |(num_available[4:1]);
    io_dis_uops_2_ready_REG <= num_available > 5'h2;
    io_dis_uops_3_ready_REG <= |(num_available[4:2]);
  end // always @(posedge)
  IssueSlot_32 slots_0 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_0_io_valid),
    .io_will_be_valid               (_slots_0_io_will_be_valid),
    .io_request                     (_slots_0_io_request),
    .io_grant                       (issue_slots_0_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (1'h0),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_0_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_21 ? _slots_4_io_out_uop_uopc : _GEN_20 ? _slots_3_io_out_uop_uopc : _GEN_19 ? _slots_2_io_out_uop_uopc : _slots_1_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_21 ? _slots_4_io_out_uop_inst : _GEN_20 ? _slots_3_io_out_uop_inst : _GEN_19 ? _slots_2_io_out_uop_inst : _slots_1_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_21 ? _slots_4_io_out_uop_debug_inst : _GEN_20 ? _slots_3_io_out_uop_debug_inst : _GEN_19 ? _slots_2_io_out_uop_debug_inst : _slots_1_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_21 ? _slots_4_io_out_uop_is_rvc : _GEN_20 ? _slots_3_io_out_uop_is_rvc : _GEN_19 ? _slots_2_io_out_uop_is_rvc : _slots_1_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_21 ? _slots_4_io_out_uop_debug_pc : _GEN_20 ? _slots_3_io_out_uop_debug_pc : _GEN_19 ? _slots_2_io_out_uop_debug_pc : _slots_1_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_21 ? _slots_4_io_out_uop_iq_type : _GEN_20 ? _slots_3_io_out_uop_iq_type : _GEN_19 ? _slots_2_io_out_uop_iq_type : _slots_1_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_21 ? _slots_4_io_out_uop_fu_code : _GEN_20 ? _slots_3_io_out_uop_fu_code : _GEN_19 ? _slots_2_io_out_uop_fu_code : _slots_1_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_21 ? _slots_4_io_out_uop_iw_state : _GEN_20 ? _slots_3_io_out_uop_iw_state : _GEN_19 ? _slots_2_io_out_uop_iw_state : _slots_1_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_21 ? _slots_4_io_out_uop_iw_p1_poisoned : _GEN_20 ? _slots_3_io_out_uop_iw_p1_poisoned : _GEN_19 ? _slots_2_io_out_uop_iw_p1_poisoned : _slots_1_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_21 ? _slots_4_io_out_uop_iw_p2_poisoned : _GEN_20 ? _slots_3_io_out_uop_iw_p2_poisoned : _GEN_19 ? _slots_2_io_out_uop_iw_p2_poisoned : _slots_1_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_21 ? _slots_4_io_out_uop_is_br : _GEN_20 ? _slots_3_io_out_uop_is_br : _GEN_19 ? _slots_2_io_out_uop_is_br : _slots_1_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_21 ? _slots_4_io_out_uop_is_jalr : _GEN_20 ? _slots_3_io_out_uop_is_jalr : _GEN_19 ? _slots_2_io_out_uop_is_jalr : _slots_1_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_21 ? _slots_4_io_out_uop_is_jal : _GEN_20 ? _slots_3_io_out_uop_is_jal : _GEN_19 ? _slots_2_io_out_uop_is_jal : _slots_1_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_21 ? _slots_4_io_out_uop_is_sfb : _GEN_20 ? _slots_3_io_out_uop_is_sfb : _GEN_19 ? _slots_2_io_out_uop_is_sfb : _slots_1_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_21 ? _slots_4_io_out_uop_br_mask : _GEN_20 ? _slots_3_io_out_uop_br_mask : _GEN_19 ? _slots_2_io_out_uop_br_mask : _slots_1_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_21 ? _slots_4_io_out_uop_br_tag : _GEN_20 ? _slots_3_io_out_uop_br_tag : _GEN_19 ? _slots_2_io_out_uop_br_tag : _slots_1_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_21 ? _slots_4_io_out_uop_ftq_idx : _GEN_20 ? _slots_3_io_out_uop_ftq_idx : _GEN_19 ? _slots_2_io_out_uop_ftq_idx : _slots_1_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_21 ? _slots_4_io_out_uop_edge_inst : _GEN_20 ? _slots_3_io_out_uop_edge_inst : _GEN_19 ? _slots_2_io_out_uop_edge_inst : _slots_1_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_21 ? _slots_4_io_out_uop_pc_lob : _GEN_20 ? _slots_3_io_out_uop_pc_lob : _GEN_19 ? _slots_2_io_out_uop_pc_lob : _slots_1_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_21 ? _slots_4_io_out_uop_taken : _GEN_20 ? _slots_3_io_out_uop_taken : _GEN_19 ? _slots_2_io_out_uop_taken : _slots_1_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_21 ? _slots_4_io_out_uop_imm_packed : _GEN_20 ? _slots_3_io_out_uop_imm_packed : _GEN_19 ? _slots_2_io_out_uop_imm_packed : _slots_1_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_21 ? _slots_4_io_out_uop_csr_addr : _GEN_20 ? _slots_3_io_out_uop_csr_addr : _GEN_19 ? _slots_2_io_out_uop_csr_addr : _slots_1_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_21 ? _slots_4_io_out_uop_rob_idx : _GEN_20 ? _slots_3_io_out_uop_rob_idx : _GEN_19 ? _slots_2_io_out_uop_rob_idx : _slots_1_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_21 ? _slots_4_io_out_uop_ldq_idx : _GEN_20 ? _slots_3_io_out_uop_ldq_idx : _GEN_19 ? _slots_2_io_out_uop_ldq_idx : _slots_1_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_21 ? _slots_4_io_out_uop_stq_idx : _GEN_20 ? _slots_3_io_out_uop_stq_idx : _GEN_19 ? _slots_2_io_out_uop_stq_idx : _slots_1_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_21 ? _slots_4_io_out_uop_rxq_idx : _GEN_20 ? _slots_3_io_out_uop_rxq_idx : _GEN_19 ? _slots_2_io_out_uop_rxq_idx : _slots_1_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_21 ? _slots_4_io_out_uop_pdst : _GEN_20 ? _slots_3_io_out_uop_pdst : _GEN_19 ? _slots_2_io_out_uop_pdst : _slots_1_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_21 ? _slots_4_io_out_uop_prs1 : _GEN_20 ? _slots_3_io_out_uop_prs1 : _GEN_19 ? _slots_2_io_out_uop_prs1 : _slots_1_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_21 ? _slots_4_io_out_uop_prs2 : _GEN_20 ? _slots_3_io_out_uop_prs2 : _GEN_19 ? _slots_2_io_out_uop_prs2 : _slots_1_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_21 ? _slots_4_io_out_uop_prs3 : _GEN_20 ? _slots_3_io_out_uop_prs3 : _GEN_19 ? _slots_2_io_out_uop_prs3 : _slots_1_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_21 ? _slots_4_io_out_uop_ppred : _GEN_20 ? _slots_3_io_out_uop_ppred : _GEN_19 ? _slots_2_io_out_uop_ppred : _slots_1_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_21 ? _slots_4_io_out_uop_prs1_busy : _GEN_20 ? _slots_3_io_out_uop_prs1_busy : _GEN_19 ? _slots_2_io_out_uop_prs1_busy : _slots_1_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_21 ? _slots_4_io_out_uop_prs2_busy : _GEN_20 ? _slots_3_io_out_uop_prs2_busy : _GEN_19 ? _slots_2_io_out_uop_prs2_busy : _slots_1_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_21 ? _slots_4_io_out_uop_prs3_busy : _GEN_20 ? _slots_3_io_out_uop_prs3_busy : _GEN_19 ? _slots_2_io_out_uop_prs3_busy : _slots_1_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_21 ? _slots_4_io_out_uop_ppred_busy : _GEN_20 ? _slots_3_io_out_uop_ppred_busy : _GEN_19 ? _slots_2_io_out_uop_ppred_busy : _slots_1_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_21 ? _slots_4_io_out_uop_stale_pdst : _GEN_20 ? _slots_3_io_out_uop_stale_pdst : _GEN_19 ? _slots_2_io_out_uop_stale_pdst : _slots_1_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_21 ? _slots_4_io_out_uop_exception : _GEN_20 ? _slots_3_io_out_uop_exception : _GEN_19 ? _slots_2_io_out_uop_exception : _slots_1_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_21 ? _slots_4_io_out_uop_exc_cause : _GEN_20 ? _slots_3_io_out_uop_exc_cause : _GEN_19 ? _slots_2_io_out_uop_exc_cause : _slots_1_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_21 ? _slots_4_io_out_uop_bypassable : _GEN_20 ? _slots_3_io_out_uop_bypassable : _GEN_19 ? _slots_2_io_out_uop_bypassable : _slots_1_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_21 ? _slots_4_io_out_uop_mem_cmd : _GEN_20 ? _slots_3_io_out_uop_mem_cmd : _GEN_19 ? _slots_2_io_out_uop_mem_cmd : _slots_1_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_21 ? _slots_4_io_out_uop_mem_size : _GEN_20 ? _slots_3_io_out_uop_mem_size : _GEN_19 ? _slots_2_io_out_uop_mem_size : _slots_1_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_21 ? _slots_4_io_out_uop_mem_signed : _GEN_20 ? _slots_3_io_out_uop_mem_signed : _GEN_19 ? _slots_2_io_out_uop_mem_signed : _slots_1_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_21 ? _slots_4_io_out_uop_is_fence : _GEN_20 ? _slots_3_io_out_uop_is_fence : _GEN_19 ? _slots_2_io_out_uop_is_fence : _slots_1_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_21 ? _slots_4_io_out_uop_is_fencei : _GEN_20 ? _slots_3_io_out_uop_is_fencei : _GEN_19 ? _slots_2_io_out_uop_is_fencei : _slots_1_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_21 ? _slots_4_io_out_uop_is_amo : _GEN_20 ? _slots_3_io_out_uop_is_amo : _GEN_19 ? _slots_2_io_out_uop_is_amo : _slots_1_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_21 ? _slots_4_io_out_uop_uses_ldq : _GEN_20 ? _slots_3_io_out_uop_uses_ldq : _GEN_19 ? _slots_2_io_out_uop_uses_ldq : _slots_1_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_21 ? _slots_4_io_out_uop_uses_stq : _GEN_20 ? _slots_3_io_out_uop_uses_stq : _GEN_19 ? _slots_2_io_out_uop_uses_stq : _slots_1_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_21 ? _slots_4_io_out_uop_is_sys_pc2epc : _GEN_20 ? _slots_3_io_out_uop_is_sys_pc2epc : _GEN_19 ? _slots_2_io_out_uop_is_sys_pc2epc : _slots_1_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_21 ? _slots_4_io_out_uop_is_unique : _GEN_20 ? _slots_3_io_out_uop_is_unique : _GEN_19 ? _slots_2_io_out_uop_is_unique : _slots_1_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_21 ? _slots_4_io_out_uop_flush_on_commit : _GEN_20 ? _slots_3_io_out_uop_flush_on_commit : _GEN_19 ? _slots_2_io_out_uop_flush_on_commit : _slots_1_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_21 ? _slots_4_io_out_uop_ldst_is_rs1 : _GEN_20 ? _slots_3_io_out_uop_ldst_is_rs1 : _GEN_19 ? _slots_2_io_out_uop_ldst_is_rs1 : _slots_1_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_21 ? _slots_4_io_out_uop_ldst : _GEN_20 ? _slots_3_io_out_uop_ldst : _GEN_19 ? _slots_2_io_out_uop_ldst : _slots_1_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_21 ? _slots_4_io_out_uop_lrs1 : _GEN_20 ? _slots_3_io_out_uop_lrs1 : _GEN_19 ? _slots_2_io_out_uop_lrs1 : _slots_1_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_21 ? _slots_4_io_out_uop_lrs2 : _GEN_20 ? _slots_3_io_out_uop_lrs2 : _GEN_19 ? _slots_2_io_out_uop_lrs2 : _slots_1_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_21 ? _slots_4_io_out_uop_lrs3 : _GEN_20 ? _slots_3_io_out_uop_lrs3 : _GEN_19 ? _slots_2_io_out_uop_lrs3 : _slots_1_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_21 ? _slots_4_io_out_uop_ldst_val : _GEN_20 ? _slots_3_io_out_uop_ldst_val : _GEN_19 ? _slots_2_io_out_uop_ldst_val : _slots_1_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_21 ? _slots_4_io_out_uop_dst_rtype : _GEN_20 ? _slots_3_io_out_uop_dst_rtype : _GEN_19 ? _slots_2_io_out_uop_dst_rtype : _slots_1_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_21 ? _slots_4_io_out_uop_lrs1_rtype : _GEN_20 ? _slots_3_io_out_uop_lrs1_rtype : _GEN_19 ? _slots_2_io_out_uop_lrs1_rtype : _slots_1_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_21 ? _slots_4_io_out_uop_lrs2_rtype : _GEN_20 ? _slots_3_io_out_uop_lrs2_rtype : _GEN_19 ? _slots_2_io_out_uop_lrs2_rtype : _slots_1_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_21 ? _slots_4_io_out_uop_frs3_en : _GEN_20 ? _slots_3_io_out_uop_frs3_en : _GEN_19 ? _slots_2_io_out_uop_frs3_en : _slots_1_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_21 ? _slots_4_io_out_uop_fp_val : _GEN_20 ? _slots_3_io_out_uop_fp_val : _GEN_19 ? _slots_2_io_out_uop_fp_val : _slots_1_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_21 ? _slots_4_io_out_uop_fp_single : _GEN_20 ? _slots_3_io_out_uop_fp_single : _GEN_19 ? _slots_2_io_out_uop_fp_single : _slots_1_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_21 ? _slots_4_io_out_uop_xcpt_pf_if : _GEN_20 ? _slots_3_io_out_uop_xcpt_pf_if : _GEN_19 ? _slots_2_io_out_uop_xcpt_pf_if : _slots_1_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_21 ? _slots_4_io_out_uop_xcpt_ae_if : _GEN_20 ? _slots_3_io_out_uop_xcpt_ae_if : _GEN_19 ? _slots_2_io_out_uop_xcpt_ae_if : _slots_1_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_21 ? _slots_4_io_out_uop_xcpt_ma_if : _GEN_20 ? _slots_3_io_out_uop_xcpt_ma_if : _GEN_19 ? _slots_2_io_out_uop_xcpt_ma_if : _slots_1_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_21 ? _slots_4_io_out_uop_bp_debug_if : _GEN_20 ? _slots_3_io_out_uop_bp_debug_if : _GEN_19 ? _slots_2_io_out_uop_bp_debug_if : _slots_1_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_21 ? _slots_4_io_out_uop_bp_xcpt_if : _GEN_20 ? _slots_3_io_out_uop_bp_xcpt_if : _GEN_19 ? _slots_2_io_out_uop_bp_xcpt_if : _slots_1_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_21 ? _slots_4_io_out_uop_debug_fsrc : _GEN_20 ? _slots_3_io_out_uop_debug_fsrc : _GEN_19 ? _slots_2_io_out_uop_debug_fsrc : _slots_1_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_21 ? _slots_4_io_out_uop_debug_tsrc : _GEN_20 ? _slots_3_io_out_uop_debug_tsrc : _GEN_19 ? _slots_2_io_out_uop_debug_tsrc : _slots_1_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (/* unused */),
    .io_out_uop_inst                (/* unused */),
    .io_out_uop_debug_inst          (/* unused */),
    .io_out_uop_is_rvc              (/* unused */),
    .io_out_uop_debug_pc            (/* unused */),
    .io_out_uop_iq_type             (/* unused */),
    .io_out_uop_fu_code             (/* unused */),
    .io_out_uop_iw_state            (/* unused */),
    .io_out_uop_iw_p1_poisoned      (/* unused */),
    .io_out_uop_iw_p2_poisoned      (/* unused */),
    .io_out_uop_is_br               (/* unused */),
    .io_out_uop_is_jalr             (/* unused */),
    .io_out_uop_is_jal              (/* unused */),
    .io_out_uop_is_sfb              (/* unused */),
    .io_out_uop_br_mask             (/* unused */),
    .io_out_uop_br_tag              (/* unused */),
    .io_out_uop_ftq_idx             (/* unused */),
    .io_out_uop_edge_inst           (/* unused */),
    .io_out_uop_pc_lob              (/* unused */),
    .io_out_uop_taken               (/* unused */),
    .io_out_uop_imm_packed          (/* unused */),
    .io_out_uop_csr_addr            (/* unused */),
    .io_out_uop_rob_idx             (/* unused */),
    .io_out_uop_ldq_idx             (/* unused */),
    .io_out_uop_stq_idx             (/* unused */),
    .io_out_uop_rxq_idx             (/* unused */),
    .io_out_uop_pdst                (/* unused */),
    .io_out_uop_prs1                (/* unused */),
    .io_out_uop_prs2                (/* unused */),
    .io_out_uop_prs3                (/* unused */),
    .io_out_uop_ppred               (/* unused */),
    .io_out_uop_prs1_busy           (/* unused */),
    .io_out_uop_prs2_busy           (/* unused */),
    .io_out_uop_prs3_busy           (/* unused */),
    .io_out_uop_ppred_busy          (/* unused */),
    .io_out_uop_stale_pdst          (/* unused */),
    .io_out_uop_exception           (/* unused */),
    .io_out_uop_exc_cause           (/* unused */),
    .io_out_uop_bypassable          (/* unused */),
    .io_out_uop_mem_cmd             (/* unused */),
    .io_out_uop_mem_size            (/* unused */),
    .io_out_uop_mem_signed          (/* unused */),
    .io_out_uop_is_fence            (/* unused */),
    .io_out_uop_is_fencei           (/* unused */),
    .io_out_uop_is_amo              (/* unused */),
    .io_out_uop_uses_ldq            (/* unused */),
    .io_out_uop_uses_stq            (/* unused */),
    .io_out_uop_is_sys_pc2epc       (/* unused */),
    .io_out_uop_is_unique           (/* unused */),
    .io_out_uop_flush_on_commit     (/* unused */),
    .io_out_uop_ldst_is_rs1         (/* unused */),
    .io_out_uop_ldst                (/* unused */),
    .io_out_uop_lrs1                (/* unused */),
    .io_out_uop_lrs2                (/* unused */),
    .io_out_uop_lrs3                (/* unused */),
    .io_out_uop_ldst_val            (/* unused */),
    .io_out_uop_dst_rtype           (/* unused */),
    .io_out_uop_lrs1_rtype          (/* unused */),
    .io_out_uop_lrs2_rtype          (/* unused */),
    .io_out_uop_frs3_en             (/* unused */),
    .io_out_uop_fp_val              (/* unused */),
    .io_out_uop_fp_single           (/* unused */),
    .io_out_uop_xcpt_pf_if          (/* unused */),
    .io_out_uop_xcpt_ae_if          (/* unused */),
    .io_out_uop_xcpt_ma_if          (/* unused */),
    .io_out_uop_bp_debug_if         (/* unused */),
    .io_out_uop_bp_xcpt_if          (/* unused */),
    .io_out_uop_debug_fsrc          (/* unused */),
    .io_out_uop_debug_tsrc          (/* unused */),
    .io_uop_uopc                    (_slots_0_io_uop_uopc),
    .io_uop_inst                    (_slots_0_io_uop_inst),
    .io_uop_debug_inst              (_slots_0_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_0_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_0_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_0_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_0_io_uop_fu_code),
    .io_uop_iw_state                (_slots_0_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_0_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_0_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_0_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_0_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_0_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_0_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_0_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_0_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_0_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_0_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_0_io_uop_pc_lob),
    .io_uop_taken                   (_slots_0_io_uop_taken),
    .io_uop_imm_packed              (_slots_0_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_0_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_0_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_0_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_0_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_0_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_0_io_uop_pdst),
    .io_uop_prs1                    (_slots_0_io_uop_prs1),
    .io_uop_prs2                    (_slots_0_io_uop_prs2),
    .io_uop_prs3                    (_slots_0_io_uop_prs3),
    .io_uop_ppred                   (_slots_0_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_0_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_0_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_0_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_0_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_0_io_uop_stale_pdst),
    .io_uop_exception               (_slots_0_io_uop_exception),
    .io_uop_exc_cause               (_slots_0_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_0_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_0_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_0_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_0_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_0_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_0_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_0_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_0_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_0_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_0_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_0_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_0_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_0_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_0_io_uop_ldst),
    .io_uop_lrs1                    (_slots_0_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_0_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_0_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_0_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_0_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_0_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_0_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_0_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_0_io_uop_fp_val),
    .io_uop_fp_single               (_slots_0_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_0_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_0_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_0_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_0_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_0_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_0_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_0_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_1 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_1_io_valid),
    .io_will_be_valid               (_slots_1_io_will_be_valid),
    .io_request                     (_slots_1_io_request),
    .io_grant                       (issue_slots_1_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (~_slots_0_io_valid),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_1_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_24 ? _slots_5_io_out_uop_uopc : _GEN_23 ? _slots_4_io_out_uop_uopc : _GEN_22 ? _slots_3_io_out_uop_uopc : _slots_2_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_24 ? _slots_5_io_out_uop_inst : _GEN_23 ? _slots_4_io_out_uop_inst : _GEN_22 ? _slots_3_io_out_uop_inst : _slots_2_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_24 ? _slots_5_io_out_uop_debug_inst : _GEN_23 ? _slots_4_io_out_uop_debug_inst : _GEN_22 ? _slots_3_io_out_uop_debug_inst : _slots_2_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_24 ? _slots_5_io_out_uop_is_rvc : _GEN_23 ? _slots_4_io_out_uop_is_rvc : _GEN_22 ? _slots_3_io_out_uop_is_rvc : _slots_2_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_24 ? _slots_5_io_out_uop_debug_pc : _GEN_23 ? _slots_4_io_out_uop_debug_pc : _GEN_22 ? _slots_3_io_out_uop_debug_pc : _slots_2_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_24 ? _slots_5_io_out_uop_iq_type : _GEN_23 ? _slots_4_io_out_uop_iq_type : _GEN_22 ? _slots_3_io_out_uop_iq_type : _slots_2_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_24 ? _slots_5_io_out_uop_fu_code : _GEN_23 ? _slots_4_io_out_uop_fu_code : _GEN_22 ? _slots_3_io_out_uop_fu_code : _slots_2_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_24 ? _slots_5_io_out_uop_iw_state : _GEN_23 ? _slots_4_io_out_uop_iw_state : _GEN_22 ? _slots_3_io_out_uop_iw_state : _slots_2_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_24 ? _slots_5_io_out_uop_iw_p1_poisoned : _GEN_23 ? _slots_4_io_out_uop_iw_p1_poisoned : _GEN_22 ? _slots_3_io_out_uop_iw_p1_poisoned : _slots_2_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_24 ? _slots_5_io_out_uop_iw_p2_poisoned : _GEN_23 ? _slots_4_io_out_uop_iw_p2_poisoned : _GEN_22 ? _slots_3_io_out_uop_iw_p2_poisoned : _slots_2_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_24 ? _slots_5_io_out_uop_is_br : _GEN_23 ? _slots_4_io_out_uop_is_br : _GEN_22 ? _slots_3_io_out_uop_is_br : _slots_2_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_24 ? _slots_5_io_out_uop_is_jalr : _GEN_23 ? _slots_4_io_out_uop_is_jalr : _GEN_22 ? _slots_3_io_out_uop_is_jalr : _slots_2_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_24 ? _slots_5_io_out_uop_is_jal : _GEN_23 ? _slots_4_io_out_uop_is_jal : _GEN_22 ? _slots_3_io_out_uop_is_jal : _slots_2_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_24 ? _slots_5_io_out_uop_is_sfb : _GEN_23 ? _slots_4_io_out_uop_is_sfb : _GEN_22 ? _slots_3_io_out_uop_is_sfb : _slots_2_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_24 ? _slots_5_io_out_uop_br_mask : _GEN_23 ? _slots_4_io_out_uop_br_mask : _GEN_22 ? _slots_3_io_out_uop_br_mask : _slots_2_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_24 ? _slots_5_io_out_uop_br_tag : _GEN_23 ? _slots_4_io_out_uop_br_tag : _GEN_22 ? _slots_3_io_out_uop_br_tag : _slots_2_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_24 ? _slots_5_io_out_uop_ftq_idx : _GEN_23 ? _slots_4_io_out_uop_ftq_idx : _GEN_22 ? _slots_3_io_out_uop_ftq_idx : _slots_2_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_24 ? _slots_5_io_out_uop_edge_inst : _GEN_23 ? _slots_4_io_out_uop_edge_inst : _GEN_22 ? _slots_3_io_out_uop_edge_inst : _slots_2_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_24 ? _slots_5_io_out_uop_pc_lob : _GEN_23 ? _slots_4_io_out_uop_pc_lob : _GEN_22 ? _slots_3_io_out_uop_pc_lob : _slots_2_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_24 ? _slots_5_io_out_uop_taken : _GEN_23 ? _slots_4_io_out_uop_taken : _GEN_22 ? _slots_3_io_out_uop_taken : _slots_2_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_24 ? _slots_5_io_out_uop_imm_packed : _GEN_23 ? _slots_4_io_out_uop_imm_packed : _GEN_22 ? _slots_3_io_out_uop_imm_packed : _slots_2_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_24 ? _slots_5_io_out_uop_csr_addr : _GEN_23 ? _slots_4_io_out_uop_csr_addr : _GEN_22 ? _slots_3_io_out_uop_csr_addr : _slots_2_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_24 ? _slots_5_io_out_uop_rob_idx : _GEN_23 ? _slots_4_io_out_uop_rob_idx : _GEN_22 ? _slots_3_io_out_uop_rob_idx : _slots_2_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_24 ? _slots_5_io_out_uop_ldq_idx : _GEN_23 ? _slots_4_io_out_uop_ldq_idx : _GEN_22 ? _slots_3_io_out_uop_ldq_idx : _slots_2_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_24 ? _slots_5_io_out_uop_stq_idx : _GEN_23 ? _slots_4_io_out_uop_stq_idx : _GEN_22 ? _slots_3_io_out_uop_stq_idx : _slots_2_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_24 ? _slots_5_io_out_uop_rxq_idx : _GEN_23 ? _slots_4_io_out_uop_rxq_idx : _GEN_22 ? _slots_3_io_out_uop_rxq_idx : _slots_2_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_24 ? _slots_5_io_out_uop_pdst : _GEN_23 ? _slots_4_io_out_uop_pdst : _GEN_22 ? _slots_3_io_out_uop_pdst : _slots_2_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_24 ? _slots_5_io_out_uop_prs1 : _GEN_23 ? _slots_4_io_out_uop_prs1 : _GEN_22 ? _slots_3_io_out_uop_prs1 : _slots_2_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_24 ? _slots_5_io_out_uop_prs2 : _GEN_23 ? _slots_4_io_out_uop_prs2 : _GEN_22 ? _slots_3_io_out_uop_prs2 : _slots_2_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_24 ? _slots_5_io_out_uop_prs3 : _GEN_23 ? _slots_4_io_out_uop_prs3 : _GEN_22 ? _slots_3_io_out_uop_prs3 : _slots_2_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_24 ? _slots_5_io_out_uop_ppred : _GEN_23 ? _slots_4_io_out_uop_ppred : _GEN_22 ? _slots_3_io_out_uop_ppred : _slots_2_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_24 ? _slots_5_io_out_uop_prs1_busy : _GEN_23 ? _slots_4_io_out_uop_prs1_busy : _GEN_22 ? _slots_3_io_out_uop_prs1_busy : _slots_2_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_24 ? _slots_5_io_out_uop_prs2_busy : _GEN_23 ? _slots_4_io_out_uop_prs2_busy : _GEN_22 ? _slots_3_io_out_uop_prs2_busy : _slots_2_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_24 ? _slots_5_io_out_uop_prs3_busy : _GEN_23 ? _slots_4_io_out_uop_prs3_busy : _GEN_22 ? _slots_3_io_out_uop_prs3_busy : _slots_2_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_24 ? _slots_5_io_out_uop_ppred_busy : _GEN_23 ? _slots_4_io_out_uop_ppred_busy : _GEN_22 ? _slots_3_io_out_uop_ppred_busy : _slots_2_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_24 ? _slots_5_io_out_uop_stale_pdst : _GEN_23 ? _slots_4_io_out_uop_stale_pdst : _GEN_22 ? _slots_3_io_out_uop_stale_pdst : _slots_2_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_24 ? _slots_5_io_out_uop_exception : _GEN_23 ? _slots_4_io_out_uop_exception : _GEN_22 ? _slots_3_io_out_uop_exception : _slots_2_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_24 ? _slots_5_io_out_uop_exc_cause : _GEN_23 ? _slots_4_io_out_uop_exc_cause : _GEN_22 ? _slots_3_io_out_uop_exc_cause : _slots_2_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_24 ? _slots_5_io_out_uop_bypassable : _GEN_23 ? _slots_4_io_out_uop_bypassable : _GEN_22 ? _slots_3_io_out_uop_bypassable : _slots_2_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_24 ? _slots_5_io_out_uop_mem_cmd : _GEN_23 ? _slots_4_io_out_uop_mem_cmd : _GEN_22 ? _slots_3_io_out_uop_mem_cmd : _slots_2_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_24 ? _slots_5_io_out_uop_mem_size : _GEN_23 ? _slots_4_io_out_uop_mem_size : _GEN_22 ? _slots_3_io_out_uop_mem_size : _slots_2_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_24 ? _slots_5_io_out_uop_mem_signed : _GEN_23 ? _slots_4_io_out_uop_mem_signed : _GEN_22 ? _slots_3_io_out_uop_mem_signed : _slots_2_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_24 ? _slots_5_io_out_uop_is_fence : _GEN_23 ? _slots_4_io_out_uop_is_fence : _GEN_22 ? _slots_3_io_out_uop_is_fence : _slots_2_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_24 ? _slots_5_io_out_uop_is_fencei : _GEN_23 ? _slots_4_io_out_uop_is_fencei : _GEN_22 ? _slots_3_io_out_uop_is_fencei : _slots_2_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_24 ? _slots_5_io_out_uop_is_amo : _GEN_23 ? _slots_4_io_out_uop_is_amo : _GEN_22 ? _slots_3_io_out_uop_is_amo : _slots_2_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_24 ? _slots_5_io_out_uop_uses_ldq : _GEN_23 ? _slots_4_io_out_uop_uses_ldq : _GEN_22 ? _slots_3_io_out_uop_uses_ldq : _slots_2_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_24 ? _slots_5_io_out_uop_uses_stq : _GEN_23 ? _slots_4_io_out_uop_uses_stq : _GEN_22 ? _slots_3_io_out_uop_uses_stq : _slots_2_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_24 ? _slots_5_io_out_uop_is_sys_pc2epc : _GEN_23 ? _slots_4_io_out_uop_is_sys_pc2epc : _GEN_22 ? _slots_3_io_out_uop_is_sys_pc2epc : _slots_2_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_24 ? _slots_5_io_out_uop_is_unique : _GEN_23 ? _slots_4_io_out_uop_is_unique : _GEN_22 ? _slots_3_io_out_uop_is_unique : _slots_2_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_24 ? _slots_5_io_out_uop_flush_on_commit : _GEN_23 ? _slots_4_io_out_uop_flush_on_commit : _GEN_22 ? _slots_3_io_out_uop_flush_on_commit : _slots_2_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_24 ? _slots_5_io_out_uop_ldst_is_rs1 : _GEN_23 ? _slots_4_io_out_uop_ldst_is_rs1 : _GEN_22 ? _slots_3_io_out_uop_ldst_is_rs1 : _slots_2_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_24 ? _slots_5_io_out_uop_ldst : _GEN_23 ? _slots_4_io_out_uop_ldst : _GEN_22 ? _slots_3_io_out_uop_ldst : _slots_2_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_24 ? _slots_5_io_out_uop_lrs1 : _GEN_23 ? _slots_4_io_out_uop_lrs1 : _GEN_22 ? _slots_3_io_out_uop_lrs1 : _slots_2_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_24 ? _slots_5_io_out_uop_lrs2 : _GEN_23 ? _slots_4_io_out_uop_lrs2 : _GEN_22 ? _slots_3_io_out_uop_lrs2 : _slots_2_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_24 ? _slots_5_io_out_uop_lrs3 : _GEN_23 ? _slots_4_io_out_uop_lrs3 : _GEN_22 ? _slots_3_io_out_uop_lrs3 : _slots_2_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_24 ? _slots_5_io_out_uop_ldst_val : _GEN_23 ? _slots_4_io_out_uop_ldst_val : _GEN_22 ? _slots_3_io_out_uop_ldst_val : _slots_2_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_24 ? _slots_5_io_out_uop_dst_rtype : _GEN_23 ? _slots_4_io_out_uop_dst_rtype : _GEN_22 ? _slots_3_io_out_uop_dst_rtype : _slots_2_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_24 ? _slots_5_io_out_uop_lrs1_rtype : _GEN_23 ? _slots_4_io_out_uop_lrs1_rtype : _GEN_22 ? _slots_3_io_out_uop_lrs1_rtype : _slots_2_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_24 ? _slots_5_io_out_uop_lrs2_rtype : _GEN_23 ? _slots_4_io_out_uop_lrs2_rtype : _GEN_22 ? _slots_3_io_out_uop_lrs2_rtype : _slots_2_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_24 ? _slots_5_io_out_uop_frs3_en : _GEN_23 ? _slots_4_io_out_uop_frs3_en : _GEN_22 ? _slots_3_io_out_uop_frs3_en : _slots_2_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_24 ? _slots_5_io_out_uop_fp_val : _GEN_23 ? _slots_4_io_out_uop_fp_val : _GEN_22 ? _slots_3_io_out_uop_fp_val : _slots_2_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_24 ? _slots_5_io_out_uop_fp_single : _GEN_23 ? _slots_4_io_out_uop_fp_single : _GEN_22 ? _slots_3_io_out_uop_fp_single : _slots_2_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_24 ? _slots_5_io_out_uop_xcpt_pf_if : _GEN_23 ? _slots_4_io_out_uop_xcpt_pf_if : _GEN_22 ? _slots_3_io_out_uop_xcpt_pf_if : _slots_2_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_24 ? _slots_5_io_out_uop_xcpt_ae_if : _GEN_23 ? _slots_4_io_out_uop_xcpt_ae_if : _GEN_22 ? _slots_3_io_out_uop_xcpt_ae_if : _slots_2_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_24 ? _slots_5_io_out_uop_xcpt_ma_if : _GEN_23 ? _slots_4_io_out_uop_xcpt_ma_if : _GEN_22 ? _slots_3_io_out_uop_xcpt_ma_if : _slots_2_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_24 ? _slots_5_io_out_uop_bp_debug_if : _GEN_23 ? _slots_4_io_out_uop_bp_debug_if : _GEN_22 ? _slots_3_io_out_uop_bp_debug_if : _slots_2_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_24 ? _slots_5_io_out_uop_bp_xcpt_if : _GEN_23 ? _slots_4_io_out_uop_bp_xcpt_if : _GEN_22 ? _slots_3_io_out_uop_bp_xcpt_if : _slots_2_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_24 ? _slots_5_io_out_uop_debug_fsrc : _GEN_23 ? _slots_4_io_out_uop_debug_fsrc : _GEN_22 ? _slots_3_io_out_uop_debug_fsrc : _slots_2_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_24 ? _slots_5_io_out_uop_debug_tsrc : _GEN_23 ? _slots_4_io_out_uop_debug_tsrc : _GEN_22 ? _slots_3_io_out_uop_debug_tsrc : _slots_2_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_1_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_1_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_1_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_1_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_1_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_1_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_1_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_1_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_1_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_1_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_1_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_1_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_1_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_1_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_1_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_1_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_1_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_1_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_1_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_1_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_1_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_1_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_1_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_1_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_1_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_1_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_1_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_1_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_1_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_1_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_1_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_1_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_1_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_1_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_1_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_1_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_1_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_1_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_1_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_1_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_1_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_1_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_1_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_1_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_1_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_1_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_1_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_1_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_1_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_1_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_1_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_1_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_1_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_1_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_1_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_1_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_1_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_1_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_1_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_1_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_1_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_1_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_1_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_1_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_1_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_1_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_1_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_1_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_1_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_1_io_uop_uopc),
    .io_uop_inst                    (_slots_1_io_uop_inst),
    .io_uop_debug_inst              (_slots_1_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_1_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_1_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_1_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_1_io_uop_fu_code),
    .io_uop_iw_state                (_slots_1_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_1_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_1_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_1_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_1_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_1_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_1_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_1_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_1_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_1_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_1_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_1_io_uop_pc_lob),
    .io_uop_taken                   (_slots_1_io_uop_taken),
    .io_uop_imm_packed              (_slots_1_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_1_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_1_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_1_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_1_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_1_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_1_io_uop_pdst),
    .io_uop_prs1                    (_slots_1_io_uop_prs1),
    .io_uop_prs2                    (_slots_1_io_uop_prs2),
    .io_uop_prs3                    (_slots_1_io_uop_prs3),
    .io_uop_ppred                   (_slots_1_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_1_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_1_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_1_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_1_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_1_io_uop_stale_pdst),
    .io_uop_exception               (_slots_1_io_uop_exception),
    .io_uop_exc_cause               (_slots_1_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_1_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_1_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_1_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_1_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_1_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_1_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_1_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_1_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_1_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_1_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_1_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_1_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_1_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_1_io_uop_ldst),
    .io_uop_lrs1                    (_slots_1_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_1_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_1_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_1_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_1_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_1_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_1_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_1_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_1_io_uop_fp_val),
    .io_uop_fp_single               (_slots_1_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_1_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_1_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_1_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_1_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_1_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_1_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_1_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_2 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_2_io_valid),
    .io_will_be_valid               (_slots_2_io_will_be_valid),
    .io_request                     (_slots_2_io_request),
    .io_grant                       (issue_slots_2_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_next_1_1to0),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_2_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_27 ? _slots_6_io_out_uop_uopc : _GEN_26 ? _slots_5_io_out_uop_uopc : _GEN_25 ? _slots_4_io_out_uop_uopc : _slots_3_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_27 ? _slots_6_io_out_uop_inst : _GEN_26 ? _slots_5_io_out_uop_inst : _GEN_25 ? _slots_4_io_out_uop_inst : _slots_3_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_27 ? _slots_6_io_out_uop_debug_inst : _GEN_26 ? _slots_5_io_out_uop_debug_inst : _GEN_25 ? _slots_4_io_out_uop_debug_inst : _slots_3_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_27 ? _slots_6_io_out_uop_is_rvc : _GEN_26 ? _slots_5_io_out_uop_is_rvc : _GEN_25 ? _slots_4_io_out_uop_is_rvc : _slots_3_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_27 ? _slots_6_io_out_uop_debug_pc : _GEN_26 ? _slots_5_io_out_uop_debug_pc : _GEN_25 ? _slots_4_io_out_uop_debug_pc : _slots_3_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_27 ? _slots_6_io_out_uop_iq_type : _GEN_26 ? _slots_5_io_out_uop_iq_type : _GEN_25 ? _slots_4_io_out_uop_iq_type : _slots_3_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_27 ? _slots_6_io_out_uop_fu_code : _GEN_26 ? _slots_5_io_out_uop_fu_code : _GEN_25 ? _slots_4_io_out_uop_fu_code : _slots_3_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_27 ? _slots_6_io_out_uop_iw_state : _GEN_26 ? _slots_5_io_out_uop_iw_state : _GEN_25 ? _slots_4_io_out_uop_iw_state : _slots_3_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_27 ? _slots_6_io_out_uop_iw_p1_poisoned : _GEN_26 ? _slots_5_io_out_uop_iw_p1_poisoned : _GEN_25 ? _slots_4_io_out_uop_iw_p1_poisoned : _slots_3_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_27 ? _slots_6_io_out_uop_iw_p2_poisoned : _GEN_26 ? _slots_5_io_out_uop_iw_p2_poisoned : _GEN_25 ? _slots_4_io_out_uop_iw_p2_poisoned : _slots_3_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_27 ? _slots_6_io_out_uop_is_br : _GEN_26 ? _slots_5_io_out_uop_is_br : _GEN_25 ? _slots_4_io_out_uop_is_br : _slots_3_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_27 ? _slots_6_io_out_uop_is_jalr : _GEN_26 ? _slots_5_io_out_uop_is_jalr : _GEN_25 ? _slots_4_io_out_uop_is_jalr : _slots_3_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_27 ? _slots_6_io_out_uop_is_jal : _GEN_26 ? _slots_5_io_out_uop_is_jal : _GEN_25 ? _slots_4_io_out_uop_is_jal : _slots_3_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_27 ? _slots_6_io_out_uop_is_sfb : _GEN_26 ? _slots_5_io_out_uop_is_sfb : _GEN_25 ? _slots_4_io_out_uop_is_sfb : _slots_3_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_27 ? _slots_6_io_out_uop_br_mask : _GEN_26 ? _slots_5_io_out_uop_br_mask : _GEN_25 ? _slots_4_io_out_uop_br_mask : _slots_3_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_27 ? _slots_6_io_out_uop_br_tag : _GEN_26 ? _slots_5_io_out_uop_br_tag : _GEN_25 ? _slots_4_io_out_uop_br_tag : _slots_3_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_27 ? _slots_6_io_out_uop_ftq_idx : _GEN_26 ? _slots_5_io_out_uop_ftq_idx : _GEN_25 ? _slots_4_io_out_uop_ftq_idx : _slots_3_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_27 ? _slots_6_io_out_uop_edge_inst : _GEN_26 ? _slots_5_io_out_uop_edge_inst : _GEN_25 ? _slots_4_io_out_uop_edge_inst : _slots_3_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_27 ? _slots_6_io_out_uop_pc_lob : _GEN_26 ? _slots_5_io_out_uop_pc_lob : _GEN_25 ? _slots_4_io_out_uop_pc_lob : _slots_3_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_27 ? _slots_6_io_out_uop_taken : _GEN_26 ? _slots_5_io_out_uop_taken : _GEN_25 ? _slots_4_io_out_uop_taken : _slots_3_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_27 ? _slots_6_io_out_uop_imm_packed : _GEN_26 ? _slots_5_io_out_uop_imm_packed : _GEN_25 ? _slots_4_io_out_uop_imm_packed : _slots_3_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_27 ? _slots_6_io_out_uop_csr_addr : _GEN_26 ? _slots_5_io_out_uop_csr_addr : _GEN_25 ? _slots_4_io_out_uop_csr_addr : _slots_3_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_27 ? _slots_6_io_out_uop_rob_idx : _GEN_26 ? _slots_5_io_out_uop_rob_idx : _GEN_25 ? _slots_4_io_out_uop_rob_idx : _slots_3_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_27 ? _slots_6_io_out_uop_ldq_idx : _GEN_26 ? _slots_5_io_out_uop_ldq_idx : _GEN_25 ? _slots_4_io_out_uop_ldq_idx : _slots_3_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_27 ? _slots_6_io_out_uop_stq_idx : _GEN_26 ? _slots_5_io_out_uop_stq_idx : _GEN_25 ? _slots_4_io_out_uop_stq_idx : _slots_3_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_27 ? _slots_6_io_out_uop_rxq_idx : _GEN_26 ? _slots_5_io_out_uop_rxq_idx : _GEN_25 ? _slots_4_io_out_uop_rxq_idx : _slots_3_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_27 ? _slots_6_io_out_uop_pdst : _GEN_26 ? _slots_5_io_out_uop_pdst : _GEN_25 ? _slots_4_io_out_uop_pdst : _slots_3_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_27 ? _slots_6_io_out_uop_prs1 : _GEN_26 ? _slots_5_io_out_uop_prs1 : _GEN_25 ? _slots_4_io_out_uop_prs1 : _slots_3_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_27 ? _slots_6_io_out_uop_prs2 : _GEN_26 ? _slots_5_io_out_uop_prs2 : _GEN_25 ? _slots_4_io_out_uop_prs2 : _slots_3_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_27 ? _slots_6_io_out_uop_prs3 : _GEN_26 ? _slots_5_io_out_uop_prs3 : _GEN_25 ? _slots_4_io_out_uop_prs3 : _slots_3_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_27 ? _slots_6_io_out_uop_ppred : _GEN_26 ? _slots_5_io_out_uop_ppred : _GEN_25 ? _slots_4_io_out_uop_ppred : _slots_3_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_27 ? _slots_6_io_out_uop_prs1_busy : _GEN_26 ? _slots_5_io_out_uop_prs1_busy : _GEN_25 ? _slots_4_io_out_uop_prs1_busy : _slots_3_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_27 ? _slots_6_io_out_uop_prs2_busy : _GEN_26 ? _slots_5_io_out_uop_prs2_busy : _GEN_25 ? _slots_4_io_out_uop_prs2_busy : _slots_3_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_27 ? _slots_6_io_out_uop_prs3_busy : _GEN_26 ? _slots_5_io_out_uop_prs3_busy : _GEN_25 ? _slots_4_io_out_uop_prs3_busy : _slots_3_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_27 ? _slots_6_io_out_uop_ppred_busy : _GEN_26 ? _slots_5_io_out_uop_ppred_busy : _GEN_25 ? _slots_4_io_out_uop_ppred_busy : _slots_3_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_27 ? _slots_6_io_out_uop_stale_pdst : _GEN_26 ? _slots_5_io_out_uop_stale_pdst : _GEN_25 ? _slots_4_io_out_uop_stale_pdst : _slots_3_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_27 ? _slots_6_io_out_uop_exception : _GEN_26 ? _slots_5_io_out_uop_exception : _GEN_25 ? _slots_4_io_out_uop_exception : _slots_3_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_27 ? _slots_6_io_out_uop_exc_cause : _GEN_26 ? _slots_5_io_out_uop_exc_cause : _GEN_25 ? _slots_4_io_out_uop_exc_cause : _slots_3_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_27 ? _slots_6_io_out_uop_bypassable : _GEN_26 ? _slots_5_io_out_uop_bypassable : _GEN_25 ? _slots_4_io_out_uop_bypassable : _slots_3_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_27 ? _slots_6_io_out_uop_mem_cmd : _GEN_26 ? _slots_5_io_out_uop_mem_cmd : _GEN_25 ? _slots_4_io_out_uop_mem_cmd : _slots_3_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_27 ? _slots_6_io_out_uop_mem_size : _GEN_26 ? _slots_5_io_out_uop_mem_size : _GEN_25 ? _slots_4_io_out_uop_mem_size : _slots_3_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_27 ? _slots_6_io_out_uop_mem_signed : _GEN_26 ? _slots_5_io_out_uop_mem_signed : _GEN_25 ? _slots_4_io_out_uop_mem_signed : _slots_3_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_27 ? _slots_6_io_out_uop_is_fence : _GEN_26 ? _slots_5_io_out_uop_is_fence : _GEN_25 ? _slots_4_io_out_uop_is_fence : _slots_3_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_27 ? _slots_6_io_out_uop_is_fencei : _GEN_26 ? _slots_5_io_out_uop_is_fencei : _GEN_25 ? _slots_4_io_out_uop_is_fencei : _slots_3_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_27 ? _slots_6_io_out_uop_is_amo : _GEN_26 ? _slots_5_io_out_uop_is_amo : _GEN_25 ? _slots_4_io_out_uop_is_amo : _slots_3_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_27 ? _slots_6_io_out_uop_uses_ldq : _GEN_26 ? _slots_5_io_out_uop_uses_ldq : _GEN_25 ? _slots_4_io_out_uop_uses_ldq : _slots_3_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_27 ? _slots_6_io_out_uop_uses_stq : _GEN_26 ? _slots_5_io_out_uop_uses_stq : _GEN_25 ? _slots_4_io_out_uop_uses_stq : _slots_3_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_27 ? _slots_6_io_out_uop_is_sys_pc2epc : _GEN_26 ? _slots_5_io_out_uop_is_sys_pc2epc : _GEN_25 ? _slots_4_io_out_uop_is_sys_pc2epc : _slots_3_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_27 ? _slots_6_io_out_uop_is_unique : _GEN_26 ? _slots_5_io_out_uop_is_unique : _GEN_25 ? _slots_4_io_out_uop_is_unique : _slots_3_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_27 ? _slots_6_io_out_uop_flush_on_commit : _GEN_26 ? _slots_5_io_out_uop_flush_on_commit : _GEN_25 ? _slots_4_io_out_uop_flush_on_commit : _slots_3_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_27 ? _slots_6_io_out_uop_ldst_is_rs1 : _GEN_26 ? _slots_5_io_out_uop_ldst_is_rs1 : _GEN_25 ? _slots_4_io_out_uop_ldst_is_rs1 : _slots_3_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_27 ? _slots_6_io_out_uop_ldst : _GEN_26 ? _slots_5_io_out_uop_ldst : _GEN_25 ? _slots_4_io_out_uop_ldst : _slots_3_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_27 ? _slots_6_io_out_uop_lrs1 : _GEN_26 ? _slots_5_io_out_uop_lrs1 : _GEN_25 ? _slots_4_io_out_uop_lrs1 : _slots_3_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_27 ? _slots_6_io_out_uop_lrs2 : _GEN_26 ? _slots_5_io_out_uop_lrs2 : _GEN_25 ? _slots_4_io_out_uop_lrs2 : _slots_3_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_27 ? _slots_6_io_out_uop_lrs3 : _GEN_26 ? _slots_5_io_out_uop_lrs3 : _GEN_25 ? _slots_4_io_out_uop_lrs3 : _slots_3_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_27 ? _slots_6_io_out_uop_ldst_val : _GEN_26 ? _slots_5_io_out_uop_ldst_val : _GEN_25 ? _slots_4_io_out_uop_ldst_val : _slots_3_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_27 ? _slots_6_io_out_uop_dst_rtype : _GEN_26 ? _slots_5_io_out_uop_dst_rtype : _GEN_25 ? _slots_4_io_out_uop_dst_rtype : _slots_3_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_27 ? _slots_6_io_out_uop_lrs1_rtype : _GEN_26 ? _slots_5_io_out_uop_lrs1_rtype : _GEN_25 ? _slots_4_io_out_uop_lrs1_rtype : _slots_3_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_27 ? _slots_6_io_out_uop_lrs2_rtype : _GEN_26 ? _slots_5_io_out_uop_lrs2_rtype : _GEN_25 ? _slots_4_io_out_uop_lrs2_rtype : _slots_3_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_27 ? _slots_6_io_out_uop_frs3_en : _GEN_26 ? _slots_5_io_out_uop_frs3_en : _GEN_25 ? _slots_4_io_out_uop_frs3_en : _slots_3_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_27 ? _slots_6_io_out_uop_fp_val : _GEN_26 ? _slots_5_io_out_uop_fp_val : _GEN_25 ? _slots_4_io_out_uop_fp_val : _slots_3_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_27 ? _slots_6_io_out_uop_fp_single : _GEN_26 ? _slots_5_io_out_uop_fp_single : _GEN_25 ? _slots_4_io_out_uop_fp_single : _slots_3_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_27 ? _slots_6_io_out_uop_xcpt_pf_if : _GEN_26 ? _slots_5_io_out_uop_xcpt_pf_if : _GEN_25 ? _slots_4_io_out_uop_xcpt_pf_if : _slots_3_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_27 ? _slots_6_io_out_uop_xcpt_ae_if : _GEN_26 ? _slots_5_io_out_uop_xcpt_ae_if : _GEN_25 ? _slots_4_io_out_uop_xcpt_ae_if : _slots_3_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_27 ? _slots_6_io_out_uop_xcpt_ma_if : _GEN_26 ? _slots_5_io_out_uop_xcpt_ma_if : _GEN_25 ? _slots_4_io_out_uop_xcpt_ma_if : _slots_3_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_27 ? _slots_6_io_out_uop_bp_debug_if : _GEN_26 ? _slots_5_io_out_uop_bp_debug_if : _GEN_25 ? _slots_4_io_out_uop_bp_debug_if : _slots_3_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_27 ? _slots_6_io_out_uop_bp_xcpt_if : _GEN_26 ? _slots_5_io_out_uop_bp_xcpt_if : _GEN_25 ? _slots_4_io_out_uop_bp_xcpt_if : _slots_3_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_27 ? _slots_6_io_out_uop_debug_fsrc : _GEN_26 ? _slots_5_io_out_uop_debug_fsrc : _GEN_25 ? _slots_4_io_out_uop_debug_fsrc : _slots_3_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_27 ? _slots_6_io_out_uop_debug_tsrc : _GEN_26 ? _slots_5_io_out_uop_debug_tsrc : _GEN_25 ? _slots_4_io_out_uop_debug_tsrc : _slots_3_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_2_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_2_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_2_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_2_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_2_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_2_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_2_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_2_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_2_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_2_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_2_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_2_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_2_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_2_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_2_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_2_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_2_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_2_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_2_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_2_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_2_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_2_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_2_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_2_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_2_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_2_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_2_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_2_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_2_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_2_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_2_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_2_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_2_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_2_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_2_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_2_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_2_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_2_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_2_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_2_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_2_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_2_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_2_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_2_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_2_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_2_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_2_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_2_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_2_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_2_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_2_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_2_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_2_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_2_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_2_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_2_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_2_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_2_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_2_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_2_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_2_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_2_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_2_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_2_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_2_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_2_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_2_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_2_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_2_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_2_io_uop_uopc),
    .io_uop_inst                    (_slots_2_io_uop_inst),
    .io_uop_debug_inst              (_slots_2_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_2_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_2_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_2_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_2_io_uop_fu_code),
    .io_uop_iw_state                (_slots_2_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_2_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_2_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_2_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_2_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_2_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_2_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_2_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_2_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_2_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_2_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_2_io_uop_pc_lob),
    .io_uop_taken                   (_slots_2_io_uop_taken),
    .io_uop_imm_packed              (_slots_2_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_2_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_2_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_2_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_2_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_2_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_2_io_uop_pdst),
    .io_uop_prs1                    (_slots_2_io_uop_prs1),
    .io_uop_prs2                    (_slots_2_io_uop_prs2),
    .io_uop_prs3                    (_slots_2_io_uop_prs3),
    .io_uop_ppred                   (_slots_2_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_2_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_2_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_2_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_2_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_2_io_uop_stale_pdst),
    .io_uop_exception               (_slots_2_io_uop_exception),
    .io_uop_exc_cause               (_slots_2_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_2_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_2_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_2_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_2_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_2_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_2_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_2_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_2_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_2_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_2_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_2_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_2_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_2_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_2_io_uop_ldst),
    .io_uop_lrs1                    (_slots_2_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_2_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_2_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_2_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_2_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_2_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_2_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_2_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_2_io_uop_fp_val),
    .io_uop_fp_single               (_slots_2_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_2_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_2_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_2_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_2_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_2_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_2_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_2_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_3 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_3_io_valid),
    .io_will_be_valid               (_slots_3_io_will_be_valid),
    .io_request                     (_slots_3_io_request),
    .io_grant                       (issue_slots_3_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_2),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_3_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_30 ? _slots_7_io_out_uop_uopc : _GEN_29 ? _slots_6_io_out_uop_uopc : _GEN_28 ? _slots_5_io_out_uop_uopc : _slots_4_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_30 ? _slots_7_io_out_uop_inst : _GEN_29 ? _slots_6_io_out_uop_inst : _GEN_28 ? _slots_5_io_out_uop_inst : _slots_4_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_30 ? _slots_7_io_out_uop_debug_inst : _GEN_29 ? _slots_6_io_out_uop_debug_inst : _GEN_28 ? _slots_5_io_out_uop_debug_inst : _slots_4_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_30 ? _slots_7_io_out_uop_is_rvc : _GEN_29 ? _slots_6_io_out_uop_is_rvc : _GEN_28 ? _slots_5_io_out_uop_is_rvc : _slots_4_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_30 ? _slots_7_io_out_uop_debug_pc : _GEN_29 ? _slots_6_io_out_uop_debug_pc : _GEN_28 ? _slots_5_io_out_uop_debug_pc : _slots_4_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_30 ? _slots_7_io_out_uop_iq_type : _GEN_29 ? _slots_6_io_out_uop_iq_type : _GEN_28 ? _slots_5_io_out_uop_iq_type : _slots_4_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_30 ? _slots_7_io_out_uop_fu_code : _GEN_29 ? _slots_6_io_out_uop_fu_code : _GEN_28 ? _slots_5_io_out_uop_fu_code : _slots_4_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_30 ? _slots_7_io_out_uop_iw_state : _GEN_29 ? _slots_6_io_out_uop_iw_state : _GEN_28 ? _slots_5_io_out_uop_iw_state : _slots_4_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_30 ? _slots_7_io_out_uop_iw_p1_poisoned : _GEN_29 ? _slots_6_io_out_uop_iw_p1_poisoned : _GEN_28 ? _slots_5_io_out_uop_iw_p1_poisoned : _slots_4_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_30 ? _slots_7_io_out_uop_iw_p2_poisoned : _GEN_29 ? _slots_6_io_out_uop_iw_p2_poisoned : _GEN_28 ? _slots_5_io_out_uop_iw_p2_poisoned : _slots_4_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_30 ? _slots_7_io_out_uop_is_br : _GEN_29 ? _slots_6_io_out_uop_is_br : _GEN_28 ? _slots_5_io_out_uop_is_br : _slots_4_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_30 ? _slots_7_io_out_uop_is_jalr : _GEN_29 ? _slots_6_io_out_uop_is_jalr : _GEN_28 ? _slots_5_io_out_uop_is_jalr : _slots_4_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_30 ? _slots_7_io_out_uop_is_jal : _GEN_29 ? _slots_6_io_out_uop_is_jal : _GEN_28 ? _slots_5_io_out_uop_is_jal : _slots_4_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_30 ? _slots_7_io_out_uop_is_sfb : _GEN_29 ? _slots_6_io_out_uop_is_sfb : _GEN_28 ? _slots_5_io_out_uop_is_sfb : _slots_4_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_30 ? _slots_7_io_out_uop_br_mask : _GEN_29 ? _slots_6_io_out_uop_br_mask : _GEN_28 ? _slots_5_io_out_uop_br_mask : _slots_4_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_30 ? _slots_7_io_out_uop_br_tag : _GEN_29 ? _slots_6_io_out_uop_br_tag : _GEN_28 ? _slots_5_io_out_uop_br_tag : _slots_4_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_30 ? _slots_7_io_out_uop_ftq_idx : _GEN_29 ? _slots_6_io_out_uop_ftq_idx : _GEN_28 ? _slots_5_io_out_uop_ftq_idx : _slots_4_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_30 ? _slots_7_io_out_uop_edge_inst : _GEN_29 ? _slots_6_io_out_uop_edge_inst : _GEN_28 ? _slots_5_io_out_uop_edge_inst : _slots_4_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_30 ? _slots_7_io_out_uop_pc_lob : _GEN_29 ? _slots_6_io_out_uop_pc_lob : _GEN_28 ? _slots_5_io_out_uop_pc_lob : _slots_4_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_30 ? _slots_7_io_out_uop_taken : _GEN_29 ? _slots_6_io_out_uop_taken : _GEN_28 ? _slots_5_io_out_uop_taken : _slots_4_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_30 ? _slots_7_io_out_uop_imm_packed : _GEN_29 ? _slots_6_io_out_uop_imm_packed : _GEN_28 ? _slots_5_io_out_uop_imm_packed : _slots_4_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_30 ? _slots_7_io_out_uop_csr_addr : _GEN_29 ? _slots_6_io_out_uop_csr_addr : _GEN_28 ? _slots_5_io_out_uop_csr_addr : _slots_4_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_30 ? _slots_7_io_out_uop_rob_idx : _GEN_29 ? _slots_6_io_out_uop_rob_idx : _GEN_28 ? _slots_5_io_out_uop_rob_idx : _slots_4_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_30 ? _slots_7_io_out_uop_ldq_idx : _GEN_29 ? _slots_6_io_out_uop_ldq_idx : _GEN_28 ? _slots_5_io_out_uop_ldq_idx : _slots_4_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_30 ? _slots_7_io_out_uop_stq_idx : _GEN_29 ? _slots_6_io_out_uop_stq_idx : _GEN_28 ? _slots_5_io_out_uop_stq_idx : _slots_4_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_30 ? _slots_7_io_out_uop_rxq_idx : _GEN_29 ? _slots_6_io_out_uop_rxq_idx : _GEN_28 ? _slots_5_io_out_uop_rxq_idx : _slots_4_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_30 ? _slots_7_io_out_uop_pdst : _GEN_29 ? _slots_6_io_out_uop_pdst : _GEN_28 ? _slots_5_io_out_uop_pdst : _slots_4_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_30 ? _slots_7_io_out_uop_prs1 : _GEN_29 ? _slots_6_io_out_uop_prs1 : _GEN_28 ? _slots_5_io_out_uop_prs1 : _slots_4_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_30 ? _slots_7_io_out_uop_prs2 : _GEN_29 ? _slots_6_io_out_uop_prs2 : _GEN_28 ? _slots_5_io_out_uop_prs2 : _slots_4_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_30 ? _slots_7_io_out_uop_prs3 : _GEN_29 ? _slots_6_io_out_uop_prs3 : _GEN_28 ? _slots_5_io_out_uop_prs3 : _slots_4_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_30 ? _slots_7_io_out_uop_ppred : _GEN_29 ? _slots_6_io_out_uop_ppred : _GEN_28 ? _slots_5_io_out_uop_ppred : _slots_4_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_30 ? _slots_7_io_out_uop_prs1_busy : _GEN_29 ? _slots_6_io_out_uop_prs1_busy : _GEN_28 ? _slots_5_io_out_uop_prs1_busy : _slots_4_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_30 ? _slots_7_io_out_uop_prs2_busy : _GEN_29 ? _slots_6_io_out_uop_prs2_busy : _GEN_28 ? _slots_5_io_out_uop_prs2_busy : _slots_4_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_30 ? _slots_7_io_out_uop_prs3_busy : _GEN_29 ? _slots_6_io_out_uop_prs3_busy : _GEN_28 ? _slots_5_io_out_uop_prs3_busy : _slots_4_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_30 ? _slots_7_io_out_uop_ppred_busy : _GEN_29 ? _slots_6_io_out_uop_ppred_busy : _GEN_28 ? _slots_5_io_out_uop_ppred_busy : _slots_4_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_30 ? _slots_7_io_out_uop_stale_pdst : _GEN_29 ? _slots_6_io_out_uop_stale_pdst : _GEN_28 ? _slots_5_io_out_uop_stale_pdst : _slots_4_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_30 ? _slots_7_io_out_uop_exception : _GEN_29 ? _slots_6_io_out_uop_exception : _GEN_28 ? _slots_5_io_out_uop_exception : _slots_4_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_30 ? _slots_7_io_out_uop_exc_cause : _GEN_29 ? _slots_6_io_out_uop_exc_cause : _GEN_28 ? _slots_5_io_out_uop_exc_cause : _slots_4_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_30 ? _slots_7_io_out_uop_bypassable : _GEN_29 ? _slots_6_io_out_uop_bypassable : _GEN_28 ? _slots_5_io_out_uop_bypassable : _slots_4_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_30 ? _slots_7_io_out_uop_mem_cmd : _GEN_29 ? _slots_6_io_out_uop_mem_cmd : _GEN_28 ? _slots_5_io_out_uop_mem_cmd : _slots_4_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_30 ? _slots_7_io_out_uop_mem_size : _GEN_29 ? _slots_6_io_out_uop_mem_size : _GEN_28 ? _slots_5_io_out_uop_mem_size : _slots_4_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_30 ? _slots_7_io_out_uop_mem_signed : _GEN_29 ? _slots_6_io_out_uop_mem_signed : _GEN_28 ? _slots_5_io_out_uop_mem_signed : _slots_4_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_30 ? _slots_7_io_out_uop_is_fence : _GEN_29 ? _slots_6_io_out_uop_is_fence : _GEN_28 ? _slots_5_io_out_uop_is_fence : _slots_4_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_30 ? _slots_7_io_out_uop_is_fencei : _GEN_29 ? _slots_6_io_out_uop_is_fencei : _GEN_28 ? _slots_5_io_out_uop_is_fencei : _slots_4_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_30 ? _slots_7_io_out_uop_is_amo : _GEN_29 ? _slots_6_io_out_uop_is_amo : _GEN_28 ? _slots_5_io_out_uop_is_amo : _slots_4_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_30 ? _slots_7_io_out_uop_uses_ldq : _GEN_29 ? _slots_6_io_out_uop_uses_ldq : _GEN_28 ? _slots_5_io_out_uop_uses_ldq : _slots_4_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_30 ? _slots_7_io_out_uop_uses_stq : _GEN_29 ? _slots_6_io_out_uop_uses_stq : _GEN_28 ? _slots_5_io_out_uop_uses_stq : _slots_4_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_30 ? _slots_7_io_out_uop_is_sys_pc2epc : _GEN_29 ? _slots_6_io_out_uop_is_sys_pc2epc : _GEN_28 ? _slots_5_io_out_uop_is_sys_pc2epc : _slots_4_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_30 ? _slots_7_io_out_uop_is_unique : _GEN_29 ? _slots_6_io_out_uop_is_unique : _GEN_28 ? _slots_5_io_out_uop_is_unique : _slots_4_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_30 ? _slots_7_io_out_uop_flush_on_commit : _GEN_29 ? _slots_6_io_out_uop_flush_on_commit : _GEN_28 ? _slots_5_io_out_uop_flush_on_commit : _slots_4_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_30 ? _slots_7_io_out_uop_ldst_is_rs1 : _GEN_29 ? _slots_6_io_out_uop_ldst_is_rs1 : _GEN_28 ? _slots_5_io_out_uop_ldst_is_rs1 : _slots_4_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_30 ? _slots_7_io_out_uop_ldst : _GEN_29 ? _slots_6_io_out_uop_ldst : _GEN_28 ? _slots_5_io_out_uop_ldst : _slots_4_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_30 ? _slots_7_io_out_uop_lrs1 : _GEN_29 ? _slots_6_io_out_uop_lrs1 : _GEN_28 ? _slots_5_io_out_uop_lrs1 : _slots_4_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_30 ? _slots_7_io_out_uop_lrs2 : _GEN_29 ? _slots_6_io_out_uop_lrs2 : _GEN_28 ? _slots_5_io_out_uop_lrs2 : _slots_4_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_30 ? _slots_7_io_out_uop_lrs3 : _GEN_29 ? _slots_6_io_out_uop_lrs3 : _GEN_28 ? _slots_5_io_out_uop_lrs3 : _slots_4_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_30 ? _slots_7_io_out_uop_ldst_val : _GEN_29 ? _slots_6_io_out_uop_ldst_val : _GEN_28 ? _slots_5_io_out_uop_ldst_val : _slots_4_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_30 ? _slots_7_io_out_uop_dst_rtype : _GEN_29 ? _slots_6_io_out_uop_dst_rtype : _GEN_28 ? _slots_5_io_out_uop_dst_rtype : _slots_4_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_30 ? _slots_7_io_out_uop_lrs1_rtype : _GEN_29 ? _slots_6_io_out_uop_lrs1_rtype : _GEN_28 ? _slots_5_io_out_uop_lrs1_rtype : _slots_4_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_30 ? _slots_7_io_out_uop_lrs2_rtype : _GEN_29 ? _slots_6_io_out_uop_lrs2_rtype : _GEN_28 ? _slots_5_io_out_uop_lrs2_rtype : _slots_4_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_30 ? _slots_7_io_out_uop_frs3_en : _GEN_29 ? _slots_6_io_out_uop_frs3_en : _GEN_28 ? _slots_5_io_out_uop_frs3_en : _slots_4_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_30 ? _slots_7_io_out_uop_fp_val : _GEN_29 ? _slots_6_io_out_uop_fp_val : _GEN_28 ? _slots_5_io_out_uop_fp_val : _slots_4_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_30 ? _slots_7_io_out_uop_fp_single : _GEN_29 ? _slots_6_io_out_uop_fp_single : _GEN_28 ? _slots_5_io_out_uop_fp_single : _slots_4_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_30 ? _slots_7_io_out_uop_xcpt_pf_if : _GEN_29 ? _slots_6_io_out_uop_xcpt_pf_if : _GEN_28 ? _slots_5_io_out_uop_xcpt_pf_if : _slots_4_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_30 ? _slots_7_io_out_uop_xcpt_ae_if : _GEN_29 ? _slots_6_io_out_uop_xcpt_ae_if : _GEN_28 ? _slots_5_io_out_uop_xcpt_ae_if : _slots_4_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_30 ? _slots_7_io_out_uop_xcpt_ma_if : _GEN_29 ? _slots_6_io_out_uop_xcpt_ma_if : _GEN_28 ? _slots_5_io_out_uop_xcpt_ma_if : _slots_4_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_30 ? _slots_7_io_out_uop_bp_debug_if : _GEN_29 ? _slots_6_io_out_uop_bp_debug_if : _GEN_28 ? _slots_5_io_out_uop_bp_debug_if : _slots_4_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_30 ? _slots_7_io_out_uop_bp_xcpt_if : _GEN_29 ? _slots_6_io_out_uop_bp_xcpt_if : _GEN_28 ? _slots_5_io_out_uop_bp_xcpt_if : _slots_4_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_30 ? _slots_7_io_out_uop_debug_fsrc : _GEN_29 ? _slots_6_io_out_uop_debug_fsrc : _GEN_28 ? _slots_5_io_out_uop_debug_fsrc : _slots_4_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_30 ? _slots_7_io_out_uop_debug_tsrc : _GEN_29 ? _slots_6_io_out_uop_debug_tsrc : _GEN_28 ? _slots_5_io_out_uop_debug_tsrc : _slots_4_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_3_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_3_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_3_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_3_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_3_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_3_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_3_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_3_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_3_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_3_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_3_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_3_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_3_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_3_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_3_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_3_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_3_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_3_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_3_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_3_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_3_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_3_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_3_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_3_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_3_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_3_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_3_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_3_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_3_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_3_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_3_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_3_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_3_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_3_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_3_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_3_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_3_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_3_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_3_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_3_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_3_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_3_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_3_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_3_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_3_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_3_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_3_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_3_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_3_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_3_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_3_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_3_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_3_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_3_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_3_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_3_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_3_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_3_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_3_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_3_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_3_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_3_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_3_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_3_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_3_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_3_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_3_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_3_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_3_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_3_io_uop_uopc),
    .io_uop_inst                    (_slots_3_io_uop_inst),
    .io_uop_debug_inst              (_slots_3_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_3_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_3_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_3_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_3_io_uop_fu_code),
    .io_uop_iw_state                (_slots_3_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_3_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_3_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_3_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_3_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_3_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_3_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_3_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_3_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_3_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_3_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_3_io_uop_pc_lob),
    .io_uop_taken                   (_slots_3_io_uop_taken),
    .io_uop_imm_packed              (_slots_3_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_3_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_3_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_3_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_3_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_3_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_3_io_uop_pdst),
    .io_uop_prs1                    (_slots_3_io_uop_prs1),
    .io_uop_prs2                    (_slots_3_io_uop_prs2),
    .io_uop_prs3                    (_slots_3_io_uop_prs3),
    .io_uop_ppred                   (_slots_3_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_3_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_3_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_3_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_3_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_3_io_uop_stale_pdst),
    .io_uop_exception               (_slots_3_io_uop_exception),
    .io_uop_exc_cause               (_slots_3_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_3_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_3_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_3_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_3_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_3_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_3_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_3_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_3_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_3_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_3_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_3_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_3_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_3_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_3_io_uop_ldst),
    .io_uop_lrs1                    (_slots_3_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_3_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_3_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_3_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_3_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_3_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_3_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_3_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_3_io_uop_fp_val),
    .io_uop_fp_single               (_slots_3_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_3_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_3_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_3_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_3_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_3_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_3_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_3_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_4 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_4_io_valid),
    .io_will_be_valid               (_slots_4_io_will_be_valid),
    .io_request                     (_slots_4_io_request),
    .io_grant                       (issue_slots_4_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_3),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_4_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_33 ? _slots_8_io_out_uop_uopc : _GEN_32 ? _slots_7_io_out_uop_uopc : _GEN_31 ? _slots_6_io_out_uop_uopc : _slots_5_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_33 ? _slots_8_io_out_uop_inst : _GEN_32 ? _slots_7_io_out_uop_inst : _GEN_31 ? _slots_6_io_out_uop_inst : _slots_5_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_33 ? _slots_8_io_out_uop_debug_inst : _GEN_32 ? _slots_7_io_out_uop_debug_inst : _GEN_31 ? _slots_6_io_out_uop_debug_inst : _slots_5_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_33 ? _slots_8_io_out_uop_is_rvc : _GEN_32 ? _slots_7_io_out_uop_is_rvc : _GEN_31 ? _slots_6_io_out_uop_is_rvc : _slots_5_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_33 ? _slots_8_io_out_uop_debug_pc : _GEN_32 ? _slots_7_io_out_uop_debug_pc : _GEN_31 ? _slots_6_io_out_uop_debug_pc : _slots_5_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_33 ? _slots_8_io_out_uop_iq_type : _GEN_32 ? _slots_7_io_out_uop_iq_type : _GEN_31 ? _slots_6_io_out_uop_iq_type : _slots_5_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_33 ? _slots_8_io_out_uop_fu_code : _GEN_32 ? _slots_7_io_out_uop_fu_code : _GEN_31 ? _slots_6_io_out_uop_fu_code : _slots_5_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_33 ? _slots_8_io_out_uop_iw_state : _GEN_32 ? _slots_7_io_out_uop_iw_state : _GEN_31 ? _slots_6_io_out_uop_iw_state : _slots_5_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_33 ? _slots_8_io_out_uop_iw_p1_poisoned : _GEN_32 ? _slots_7_io_out_uop_iw_p1_poisoned : _GEN_31 ? _slots_6_io_out_uop_iw_p1_poisoned : _slots_5_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_33 ? _slots_8_io_out_uop_iw_p2_poisoned : _GEN_32 ? _slots_7_io_out_uop_iw_p2_poisoned : _GEN_31 ? _slots_6_io_out_uop_iw_p2_poisoned : _slots_5_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_33 ? _slots_8_io_out_uop_is_br : _GEN_32 ? _slots_7_io_out_uop_is_br : _GEN_31 ? _slots_6_io_out_uop_is_br : _slots_5_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_33 ? _slots_8_io_out_uop_is_jalr : _GEN_32 ? _slots_7_io_out_uop_is_jalr : _GEN_31 ? _slots_6_io_out_uop_is_jalr : _slots_5_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_33 ? _slots_8_io_out_uop_is_jal : _GEN_32 ? _slots_7_io_out_uop_is_jal : _GEN_31 ? _slots_6_io_out_uop_is_jal : _slots_5_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_33 ? _slots_8_io_out_uop_is_sfb : _GEN_32 ? _slots_7_io_out_uop_is_sfb : _GEN_31 ? _slots_6_io_out_uop_is_sfb : _slots_5_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_33 ? _slots_8_io_out_uop_br_mask : _GEN_32 ? _slots_7_io_out_uop_br_mask : _GEN_31 ? _slots_6_io_out_uop_br_mask : _slots_5_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_33 ? _slots_8_io_out_uop_br_tag : _GEN_32 ? _slots_7_io_out_uop_br_tag : _GEN_31 ? _slots_6_io_out_uop_br_tag : _slots_5_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_33 ? _slots_8_io_out_uop_ftq_idx : _GEN_32 ? _slots_7_io_out_uop_ftq_idx : _GEN_31 ? _slots_6_io_out_uop_ftq_idx : _slots_5_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_33 ? _slots_8_io_out_uop_edge_inst : _GEN_32 ? _slots_7_io_out_uop_edge_inst : _GEN_31 ? _slots_6_io_out_uop_edge_inst : _slots_5_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_33 ? _slots_8_io_out_uop_pc_lob : _GEN_32 ? _slots_7_io_out_uop_pc_lob : _GEN_31 ? _slots_6_io_out_uop_pc_lob : _slots_5_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_33 ? _slots_8_io_out_uop_taken : _GEN_32 ? _slots_7_io_out_uop_taken : _GEN_31 ? _slots_6_io_out_uop_taken : _slots_5_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_33 ? _slots_8_io_out_uop_imm_packed : _GEN_32 ? _slots_7_io_out_uop_imm_packed : _GEN_31 ? _slots_6_io_out_uop_imm_packed : _slots_5_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_33 ? _slots_8_io_out_uop_csr_addr : _GEN_32 ? _slots_7_io_out_uop_csr_addr : _GEN_31 ? _slots_6_io_out_uop_csr_addr : _slots_5_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_33 ? _slots_8_io_out_uop_rob_idx : _GEN_32 ? _slots_7_io_out_uop_rob_idx : _GEN_31 ? _slots_6_io_out_uop_rob_idx : _slots_5_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_33 ? _slots_8_io_out_uop_ldq_idx : _GEN_32 ? _slots_7_io_out_uop_ldq_idx : _GEN_31 ? _slots_6_io_out_uop_ldq_idx : _slots_5_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_33 ? _slots_8_io_out_uop_stq_idx : _GEN_32 ? _slots_7_io_out_uop_stq_idx : _GEN_31 ? _slots_6_io_out_uop_stq_idx : _slots_5_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_33 ? _slots_8_io_out_uop_rxq_idx : _GEN_32 ? _slots_7_io_out_uop_rxq_idx : _GEN_31 ? _slots_6_io_out_uop_rxq_idx : _slots_5_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_33 ? _slots_8_io_out_uop_pdst : _GEN_32 ? _slots_7_io_out_uop_pdst : _GEN_31 ? _slots_6_io_out_uop_pdst : _slots_5_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_33 ? _slots_8_io_out_uop_prs1 : _GEN_32 ? _slots_7_io_out_uop_prs1 : _GEN_31 ? _slots_6_io_out_uop_prs1 : _slots_5_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_33 ? _slots_8_io_out_uop_prs2 : _GEN_32 ? _slots_7_io_out_uop_prs2 : _GEN_31 ? _slots_6_io_out_uop_prs2 : _slots_5_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_33 ? _slots_8_io_out_uop_prs3 : _GEN_32 ? _slots_7_io_out_uop_prs3 : _GEN_31 ? _slots_6_io_out_uop_prs3 : _slots_5_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_33 ? _slots_8_io_out_uop_ppred : _GEN_32 ? _slots_7_io_out_uop_ppred : _GEN_31 ? _slots_6_io_out_uop_ppred : _slots_5_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_33 ? _slots_8_io_out_uop_prs1_busy : _GEN_32 ? _slots_7_io_out_uop_prs1_busy : _GEN_31 ? _slots_6_io_out_uop_prs1_busy : _slots_5_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_33 ? _slots_8_io_out_uop_prs2_busy : _GEN_32 ? _slots_7_io_out_uop_prs2_busy : _GEN_31 ? _slots_6_io_out_uop_prs2_busy : _slots_5_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_33 ? _slots_8_io_out_uop_prs3_busy : _GEN_32 ? _slots_7_io_out_uop_prs3_busy : _GEN_31 ? _slots_6_io_out_uop_prs3_busy : _slots_5_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_33 ? _slots_8_io_out_uop_ppred_busy : _GEN_32 ? _slots_7_io_out_uop_ppred_busy : _GEN_31 ? _slots_6_io_out_uop_ppred_busy : _slots_5_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_33 ? _slots_8_io_out_uop_stale_pdst : _GEN_32 ? _slots_7_io_out_uop_stale_pdst : _GEN_31 ? _slots_6_io_out_uop_stale_pdst : _slots_5_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_33 ? _slots_8_io_out_uop_exception : _GEN_32 ? _slots_7_io_out_uop_exception : _GEN_31 ? _slots_6_io_out_uop_exception : _slots_5_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_33 ? _slots_8_io_out_uop_exc_cause : _GEN_32 ? _slots_7_io_out_uop_exc_cause : _GEN_31 ? _slots_6_io_out_uop_exc_cause : _slots_5_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_33 ? _slots_8_io_out_uop_bypassable : _GEN_32 ? _slots_7_io_out_uop_bypassable : _GEN_31 ? _slots_6_io_out_uop_bypassable : _slots_5_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_33 ? _slots_8_io_out_uop_mem_cmd : _GEN_32 ? _slots_7_io_out_uop_mem_cmd : _GEN_31 ? _slots_6_io_out_uop_mem_cmd : _slots_5_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_33 ? _slots_8_io_out_uop_mem_size : _GEN_32 ? _slots_7_io_out_uop_mem_size : _GEN_31 ? _slots_6_io_out_uop_mem_size : _slots_5_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_33 ? _slots_8_io_out_uop_mem_signed : _GEN_32 ? _slots_7_io_out_uop_mem_signed : _GEN_31 ? _slots_6_io_out_uop_mem_signed : _slots_5_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_33 ? _slots_8_io_out_uop_is_fence : _GEN_32 ? _slots_7_io_out_uop_is_fence : _GEN_31 ? _slots_6_io_out_uop_is_fence : _slots_5_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_33 ? _slots_8_io_out_uop_is_fencei : _GEN_32 ? _slots_7_io_out_uop_is_fencei : _GEN_31 ? _slots_6_io_out_uop_is_fencei : _slots_5_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_33 ? _slots_8_io_out_uop_is_amo : _GEN_32 ? _slots_7_io_out_uop_is_amo : _GEN_31 ? _slots_6_io_out_uop_is_amo : _slots_5_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_33 ? _slots_8_io_out_uop_uses_ldq : _GEN_32 ? _slots_7_io_out_uop_uses_ldq : _GEN_31 ? _slots_6_io_out_uop_uses_ldq : _slots_5_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_33 ? _slots_8_io_out_uop_uses_stq : _GEN_32 ? _slots_7_io_out_uop_uses_stq : _GEN_31 ? _slots_6_io_out_uop_uses_stq : _slots_5_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_33 ? _slots_8_io_out_uop_is_sys_pc2epc : _GEN_32 ? _slots_7_io_out_uop_is_sys_pc2epc : _GEN_31 ? _slots_6_io_out_uop_is_sys_pc2epc : _slots_5_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_33 ? _slots_8_io_out_uop_is_unique : _GEN_32 ? _slots_7_io_out_uop_is_unique : _GEN_31 ? _slots_6_io_out_uop_is_unique : _slots_5_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_33 ? _slots_8_io_out_uop_flush_on_commit : _GEN_32 ? _slots_7_io_out_uop_flush_on_commit : _GEN_31 ? _slots_6_io_out_uop_flush_on_commit : _slots_5_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_33 ? _slots_8_io_out_uop_ldst_is_rs1 : _GEN_32 ? _slots_7_io_out_uop_ldst_is_rs1 : _GEN_31 ? _slots_6_io_out_uop_ldst_is_rs1 : _slots_5_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_33 ? _slots_8_io_out_uop_ldst : _GEN_32 ? _slots_7_io_out_uop_ldst : _GEN_31 ? _slots_6_io_out_uop_ldst : _slots_5_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_33 ? _slots_8_io_out_uop_lrs1 : _GEN_32 ? _slots_7_io_out_uop_lrs1 : _GEN_31 ? _slots_6_io_out_uop_lrs1 : _slots_5_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_33 ? _slots_8_io_out_uop_lrs2 : _GEN_32 ? _slots_7_io_out_uop_lrs2 : _GEN_31 ? _slots_6_io_out_uop_lrs2 : _slots_5_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_33 ? _slots_8_io_out_uop_lrs3 : _GEN_32 ? _slots_7_io_out_uop_lrs3 : _GEN_31 ? _slots_6_io_out_uop_lrs3 : _slots_5_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_33 ? _slots_8_io_out_uop_ldst_val : _GEN_32 ? _slots_7_io_out_uop_ldst_val : _GEN_31 ? _slots_6_io_out_uop_ldst_val : _slots_5_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_33 ? _slots_8_io_out_uop_dst_rtype : _GEN_32 ? _slots_7_io_out_uop_dst_rtype : _GEN_31 ? _slots_6_io_out_uop_dst_rtype : _slots_5_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_33 ? _slots_8_io_out_uop_lrs1_rtype : _GEN_32 ? _slots_7_io_out_uop_lrs1_rtype : _GEN_31 ? _slots_6_io_out_uop_lrs1_rtype : _slots_5_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_33 ? _slots_8_io_out_uop_lrs2_rtype : _GEN_32 ? _slots_7_io_out_uop_lrs2_rtype : _GEN_31 ? _slots_6_io_out_uop_lrs2_rtype : _slots_5_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_33 ? _slots_8_io_out_uop_frs3_en : _GEN_32 ? _slots_7_io_out_uop_frs3_en : _GEN_31 ? _slots_6_io_out_uop_frs3_en : _slots_5_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_33 ? _slots_8_io_out_uop_fp_val : _GEN_32 ? _slots_7_io_out_uop_fp_val : _GEN_31 ? _slots_6_io_out_uop_fp_val : _slots_5_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_33 ? _slots_8_io_out_uop_fp_single : _GEN_32 ? _slots_7_io_out_uop_fp_single : _GEN_31 ? _slots_6_io_out_uop_fp_single : _slots_5_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_33 ? _slots_8_io_out_uop_xcpt_pf_if : _GEN_32 ? _slots_7_io_out_uop_xcpt_pf_if : _GEN_31 ? _slots_6_io_out_uop_xcpt_pf_if : _slots_5_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_33 ? _slots_8_io_out_uop_xcpt_ae_if : _GEN_32 ? _slots_7_io_out_uop_xcpt_ae_if : _GEN_31 ? _slots_6_io_out_uop_xcpt_ae_if : _slots_5_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_33 ? _slots_8_io_out_uop_xcpt_ma_if : _GEN_32 ? _slots_7_io_out_uop_xcpt_ma_if : _GEN_31 ? _slots_6_io_out_uop_xcpt_ma_if : _slots_5_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_33 ? _slots_8_io_out_uop_bp_debug_if : _GEN_32 ? _slots_7_io_out_uop_bp_debug_if : _GEN_31 ? _slots_6_io_out_uop_bp_debug_if : _slots_5_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_33 ? _slots_8_io_out_uop_bp_xcpt_if : _GEN_32 ? _slots_7_io_out_uop_bp_xcpt_if : _GEN_31 ? _slots_6_io_out_uop_bp_xcpt_if : _slots_5_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_33 ? _slots_8_io_out_uop_debug_fsrc : _GEN_32 ? _slots_7_io_out_uop_debug_fsrc : _GEN_31 ? _slots_6_io_out_uop_debug_fsrc : _slots_5_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_33 ? _slots_8_io_out_uop_debug_tsrc : _GEN_32 ? _slots_7_io_out_uop_debug_tsrc : _GEN_31 ? _slots_6_io_out_uop_debug_tsrc : _slots_5_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_4_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_4_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_4_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_4_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_4_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_4_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_4_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_4_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_4_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_4_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_4_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_4_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_4_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_4_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_4_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_4_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_4_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_4_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_4_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_4_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_4_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_4_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_4_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_4_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_4_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_4_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_4_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_4_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_4_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_4_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_4_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_4_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_4_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_4_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_4_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_4_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_4_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_4_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_4_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_4_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_4_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_4_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_4_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_4_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_4_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_4_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_4_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_4_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_4_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_4_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_4_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_4_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_4_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_4_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_4_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_4_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_4_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_4_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_4_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_4_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_4_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_4_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_4_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_4_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_4_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_4_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_4_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_4_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_4_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_4_io_uop_uopc),
    .io_uop_inst                    (_slots_4_io_uop_inst),
    .io_uop_debug_inst              (_slots_4_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_4_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_4_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_4_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_4_io_uop_fu_code),
    .io_uop_iw_state                (_slots_4_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_4_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_4_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_4_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_4_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_4_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_4_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_4_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_4_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_4_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_4_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_4_io_uop_pc_lob),
    .io_uop_taken                   (_slots_4_io_uop_taken),
    .io_uop_imm_packed              (_slots_4_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_4_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_4_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_4_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_4_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_4_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_4_io_uop_pdst),
    .io_uop_prs1                    (_slots_4_io_uop_prs1),
    .io_uop_prs2                    (_slots_4_io_uop_prs2),
    .io_uop_prs3                    (_slots_4_io_uop_prs3),
    .io_uop_ppred                   (_slots_4_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_4_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_4_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_4_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_4_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_4_io_uop_stale_pdst),
    .io_uop_exception               (_slots_4_io_uop_exception),
    .io_uop_exc_cause               (_slots_4_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_4_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_4_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_4_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_4_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_4_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_4_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_4_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_4_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_4_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_4_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_4_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_4_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_4_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_4_io_uop_ldst),
    .io_uop_lrs1                    (_slots_4_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_4_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_4_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_4_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_4_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_4_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_4_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_4_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_4_io_uop_fp_val),
    .io_uop_fp_single               (_slots_4_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_4_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_4_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_4_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_4_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_4_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_4_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_4_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_5 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_5_io_valid),
    .io_will_be_valid               (_slots_5_io_will_be_valid),
    .io_request                     (_slots_5_io_request),
    .io_grant                       (issue_slots_5_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_4),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_5_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_36 ? _slots_9_io_out_uop_uopc : _GEN_35 ? _slots_8_io_out_uop_uopc : _GEN_34 ? _slots_7_io_out_uop_uopc : _slots_6_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_36 ? _slots_9_io_out_uop_inst : _GEN_35 ? _slots_8_io_out_uop_inst : _GEN_34 ? _slots_7_io_out_uop_inst : _slots_6_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_36 ? _slots_9_io_out_uop_debug_inst : _GEN_35 ? _slots_8_io_out_uop_debug_inst : _GEN_34 ? _slots_7_io_out_uop_debug_inst : _slots_6_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_36 ? _slots_9_io_out_uop_is_rvc : _GEN_35 ? _slots_8_io_out_uop_is_rvc : _GEN_34 ? _slots_7_io_out_uop_is_rvc : _slots_6_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_36 ? _slots_9_io_out_uop_debug_pc : _GEN_35 ? _slots_8_io_out_uop_debug_pc : _GEN_34 ? _slots_7_io_out_uop_debug_pc : _slots_6_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_36 ? _slots_9_io_out_uop_iq_type : _GEN_35 ? _slots_8_io_out_uop_iq_type : _GEN_34 ? _slots_7_io_out_uop_iq_type : _slots_6_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_36 ? _slots_9_io_out_uop_fu_code : _GEN_35 ? _slots_8_io_out_uop_fu_code : _GEN_34 ? _slots_7_io_out_uop_fu_code : _slots_6_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_36 ? _slots_9_io_out_uop_iw_state : _GEN_35 ? _slots_8_io_out_uop_iw_state : _GEN_34 ? _slots_7_io_out_uop_iw_state : _slots_6_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_36 ? _slots_9_io_out_uop_iw_p1_poisoned : _GEN_35 ? _slots_8_io_out_uop_iw_p1_poisoned : _GEN_34 ? _slots_7_io_out_uop_iw_p1_poisoned : _slots_6_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_36 ? _slots_9_io_out_uop_iw_p2_poisoned : _GEN_35 ? _slots_8_io_out_uop_iw_p2_poisoned : _GEN_34 ? _slots_7_io_out_uop_iw_p2_poisoned : _slots_6_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_36 ? _slots_9_io_out_uop_is_br : _GEN_35 ? _slots_8_io_out_uop_is_br : _GEN_34 ? _slots_7_io_out_uop_is_br : _slots_6_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_36 ? _slots_9_io_out_uop_is_jalr : _GEN_35 ? _slots_8_io_out_uop_is_jalr : _GEN_34 ? _slots_7_io_out_uop_is_jalr : _slots_6_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_36 ? _slots_9_io_out_uop_is_jal : _GEN_35 ? _slots_8_io_out_uop_is_jal : _GEN_34 ? _slots_7_io_out_uop_is_jal : _slots_6_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_36 ? _slots_9_io_out_uop_is_sfb : _GEN_35 ? _slots_8_io_out_uop_is_sfb : _GEN_34 ? _slots_7_io_out_uop_is_sfb : _slots_6_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_36 ? _slots_9_io_out_uop_br_mask : _GEN_35 ? _slots_8_io_out_uop_br_mask : _GEN_34 ? _slots_7_io_out_uop_br_mask : _slots_6_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_36 ? _slots_9_io_out_uop_br_tag : _GEN_35 ? _slots_8_io_out_uop_br_tag : _GEN_34 ? _slots_7_io_out_uop_br_tag : _slots_6_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_36 ? _slots_9_io_out_uop_ftq_idx : _GEN_35 ? _slots_8_io_out_uop_ftq_idx : _GEN_34 ? _slots_7_io_out_uop_ftq_idx : _slots_6_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_36 ? _slots_9_io_out_uop_edge_inst : _GEN_35 ? _slots_8_io_out_uop_edge_inst : _GEN_34 ? _slots_7_io_out_uop_edge_inst : _slots_6_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_36 ? _slots_9_io_out_uop_pc_lob : _GEN_35 ? _slots_8_io_out_uop_pc_lob : _GEN_34 ? _slots_7_io_out_uop_pc_lob : _slots_6_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_36 ? _slots_9_io_out_uop_taken : _GEN_35 ? _slots_8_io_out_uop_taken : _GEN_34 ? _slots_7_io_out_uop_taken : _slots_6_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_36 ? _slots_9_io_out_uop_imm_packed : _GEN_35 ? _slots_8_io_out_uop_imm_packed : _GEN_34 ? _slots_7_io_out_uop_imm_packed : _slots_6_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_36 ? _slots_9_io_out_uop_csr_addr : _GEN_35 ? _slots_8_io_out_uop_csr_addr : _GEN_34 ? _slots_7_io_out_uop_csr_addr : _slots_6_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_36 ? _slots_9_io_out_uop_rob_idx : _GEN_35 ? _slots_8_io_out_uop_rob_idx : _GEN_34 ? _slots_7_io_out_uop_rob_idx : _slots_6_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_36 ? _slots_9_io_out_uop_ldq_idx : _GEN_35 ? _slots_8_io_out_uop_ldq_idx : _GEN_34 ? _slots_7_io_out_uop_ldq_idx : _slots_6_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_36 ? _slots_9_io_out_uop_stq_idx : _GEN_35 ? _slots_8_io_out_uop_stq_idx : _GEN_34 ? _slots_7_io_out_uop_stq_idx : _slots_6_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_36 ? _slots_9_io_out_uop_rxq_idx : _GEN_35 ? _slots_8_io_out_uop_rxq_idx : _GEN_34 ? _slots_7_io_out_uop_rxq_idx : _slots_6_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_36 ? _slots_9_io_out_uop_pdst : _GEN_35 ? _slots_8_io_out_uop_pdst : _GEN_34 ? _slots_7_io_out_uop_pdst : _slots_6_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_36 ? _slots_9_io_out_uop_prs1 : _GEN_35 ? _slots_8_io_out_uop_prs1 : _GEN_34 ? _slots_7_io_out_uop_prs1 : _slots_6_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_36 ? _slots_9_io_out_uop_prs2 : _GEN_35 ? _slots_8_io_out_uop_prs2 : _GEN_34 ? _slots_7_io_out_uop_prs2 : _slots_6_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_36 ? _slots_9_io_out_uop_prs3 : _GEN_35 ? _slots_8_io_out_uop_prs3 : _GEN_34 ? _slots_7_io_out_uop_prs3 : _slots_6_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_36 ? _slots_9_io_out_uop_ppred : _GEN_35 ? _slots_8_io_out_uop_ppred : _GEN_34 ? _slots_7_io_out_uop_ppred : _slots_6_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_36 ? _slots_9_io_out_uop_prs1_busy : _GEN_35 ? _slots_8_io_out_uop_prs1_busy : _GEN_34 ? _slots_7_io_out_uop_prs1_busy : _slots_6_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_36 ? _slots_9_io_out_uop_prs2_busy : _GEN_35 ? _slots_8_io_out_uop_prs2_busy : _GEN_34 ? _slots_7_io_out_uop_prs2_busy : _slots_6_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_36 ? _slots_9_io_out_uop_prs3_busy : _GEN_35 ? _slots_8_io_out_uop_prs3_busy : _GEN_34 ? _slots_7_io_out_uop_prs3_busy : _slots_6_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_36 ? _slots_9_io_out_uop_ppred_busy : _GEN_35 ? _slots_8_io_out_uop_ppred_busy : _GEN_34 ? _slots_7_io_out_uop_ppred_busy : _slots_6_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_36 ? _slots_9_io_out_uop_stale_pdst : _GEN_35 ? _slots_8_io_out_uop_stale_pdst : _GEN_34 ? _slots_7_io_out_uop_stale_pdst : _slots_6_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_36 ? _slots_9_io_out_uop_exception : _GEN_35 ? _slots_8_io_out_uop_exception : _GEN_34 ? _slots_7_io_out_uop_exception : _slots_6_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_36 ? _slots_9_io_out_uop_exc_cause : _GEN_35 ? _slots_8_io_out_uop_exc_cause : _GEN_34 ? _slots_7_io_out_uop_exc_cause : _slots_6_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_36 ? _slots_9_io_out_uop_bypassable : _GEN_35 ? _slots_8_io_out_uop_bypassable : _GEN_34 ? _slots_7_io_out_uop_bypassable : _slots_6_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_36 ? _slots_9_io_out_uop_mem_cmd : _GEN_35 ? _slots_8_io_out_uop_mem_cmd : _GEN_34 ? _slots_7_io_out_uop_mem_cmd : _slots_6_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_36 ? _slots_9_io_out_uop_mem_size : _GEN_35 ? _slots_8_io_out_uop_mem_size : _GEN_34 ? _slots_7_io_out_uop_mem_size : _slots_6_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_36 ? _slots_9_io_out_uop_mem_signed : _GEN_35 ? _slots_8_io_out_uop_mem_signed : _GEN_34 ? _slots_7_io_out_uop_mem_signed : _slots_6_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_36 ? _slots_9_io_out_uop_is_fence : _GEN_35 ? _slots_8_io_out_uop_is_fence : _GEN_34 ? _slots_7_io_out_uop_is_fence : _slots_6_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_36 ? _slots_9_io_out_uop_is_fencei : _GEN_35 ? _slots_8_io_out_uop_is_fencei : _GEN_34 ? _slots_7_io_out_uop_is_fencei : _slots_6_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_36 ? _slots_9_io_out_uop_is_amo : _GEN_35 ? _slots_8_io_out_uop_is_amo : _GEN_34 ? _slots_7_io_out_uop_is_amo : _slots_6_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_36 ? _slots_9_io_out_uop_uses_ldq : _GEN_35 ? _slots_8_io_out_uop_uses_ldq : _GEN_34 ? _slots_7_io_out_uop_uses_ldq : _slots_6_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_36 ? _slots_9_io_out_uop_uses_stq : _GEN_35 ? _slots_8_io_out_uop_uses_stq : _GEN_34 ? _slots_7_io_out_uop_uses_stq : _slots_6_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_36 ? _slots_9_io_out_uop_is_sys_pc2epc : _GEN_35 ? _slots_8_io_out_uop_is_sys_pc2epc : _GEN_34 ? _slots_7_io_out_uop_is_sys_pc2epc : _slots_6_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_36 ? _slots_9_io_out_uop_is_unique : _GEN_35 ? _slots_8_io_out_uop_is_unique : _GEN_34 ? _slots_7_io_out_uop_is_unique : _slots_6_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_36 ? _slots_9_io_out_uop_flush_on_commit : _GEN_35 ? _slots_8_io_out_uop_flush_on_commit : _GEN_34 ? _slots_7_io_out_uop_flush_on_commit : _slots_6_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_36 ? _slots_9_io_out_uop_ldst_is_rs1 : _GEN_35 ? _slots_8_io_out_uop_ldst_is_rs1 : _GEN_34 ? _slots_7_io_out_uop_ldst_is_rs1 : _slots_6_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_36 ? _slots_9_io_out_uop_ldst : _GEN_35 ? _slots_8_io_out_uop_ldst : _GEN_34 ? _slots_7_io_out_uop_ldst : _slots_6_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_36 ? _slots_9_io_out_uop_lrs1 : _GEN_35 ? _slots_8_io_out_uop_lrs1 : _GEN_34 ? _slots_7_io_out_uop_lrs1 : _slots_6_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_36 ? _slots_9_io_out_uop_lrs2 : _GEN_35 ? _slots_8_io_out_uop_lrs2 : _GEN_34 ? _slots_7_io_out_uop_lrs2 : _slots_6_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_36 ? _slots_9_io_out_uop_lrs3 : _GEN_35 ? _slots_8_io_out_uop_lrs3 : _GEN_34 ? _slots_7_io_out_uop_lrs3 : _slots_6_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_36 ? _slots_9_io_out_uop_ldst_val : _GEN_35 ? _slots_8_io_out_uop_ldst_val : _GEN_34 ? _slots_7_io_out_uop_ldst_val : _slots_6_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_36 ? _slots_9_io_out_uop_dst_rtype : _GEN_35 ? _slots_8_io_out_uop_dst_rtype : _GEN_34 ? _slots_7_io_out_uop_dst_rtype : _slots_6_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_36 ? _slots_9_io_out_uop_lrs1_rtype : _GEN_35 ? _slots_8_io_out_uop_lrs1_rtype : _GEN_34 ? _slots_7_io_out_uop_lrs1_rtype : _slots_6_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_36 ? _slots_9_io_out_uop_lrs2_rtype : _GEN_35 ? _slots_8_io_out_uop_lrs2_rtype : _GEN_34 ? _slots_7_io_out_uop_lrs2_rtype : _slots_6_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_36 ? _slots_9_io_out_uop_frs3_en : _GEN_35 ? _slots_8_io_out_uop_frs3_en : _GEN_34 ? _slots_7_io_out_uop_frs3_en : _slots_6_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_36 ? _slots_9_io_out_uop_fp_val : _GEN_35 ? _slots_8_io_out_uop_fp_val : _GEN_34 ? _slots_7_io_out_uop_fp_val : _slots_6_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_36 ? _slots_9_io_out_uop_fp_single : _GEN_35 ? _slots_8_io_out_uop_fp_single : _GEN_34 ? _slots_7_io_out_uop_fp_single : _slots_6_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_36 ? _slots_9_io_out_uop_xcpt_pf_if : _GEN_35 ? _slots_8_io_out_uop_xcpt_pf_if : _GEN_34 ? _slots_7_io_out_uop_xcpt_pf_if : _slots_6_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_36 ? _slots_9_io_out_uop_xcpt_ae_if : _GEN_35 ? _slots_8_io_out_uop_xcpt_ae_if : _GEN_34 ? _slots_7_io_out_uop_xcpt_ae_if : _slots_6_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_36 ? _slots_9_io_out_uop_xcpt_ma_if : _GEN_35 ? _slots_8_io_out_uop_xcpt_ma_if : _GEN_34 ? _slots_7_io_out_uop_xcpt_ma_if : _slots_6_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_36 ? _slots_9_io_out_uop_bp_debug_if : _GEN_35 ? _slots_8_io_out_uop_bp_debug_if : _GEN_34 ? _slots_7_io_out_uop_bp_debug_if : _slots_6_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_36 ? _slots_9_io_out_uop_bp_xcpt_if : _GEN_35 ? _slots_8_io_out_uop_bp_xcpt_if : _GEN_34 ? _slots_7_io_out_uop_bp_xcpt_if : _slots_6_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_36 ? _slots_9_io_out_uop_debug_fsrc : _GEN_35 ? _slots_8_io_out_uop_debug_fsrc : _GEN_34 ? _slots_7_io_out_uop_debug_fsrc : _slots_6_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_36 ? _slots_9_io_out_uop_debug_tsrc : _GEN_35 ? _slots_8_io_out_uop_debug_tsrc : _GEN_34 ? _slots_7_io_out_uop_debug_tsrc : _slots_6_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_5_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_5_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_5_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_5_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_5_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_5_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_5_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_5_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_5_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_5_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_5_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_5_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_5_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_5_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_5_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_5_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_5_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_5_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_5_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_5_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_5_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_5_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_5_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_5_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_5_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_5_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_5_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_5_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_5_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_5_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_5_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_5_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_5_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_5_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_5_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_5_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_5_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_5_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_5_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_5_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_5_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_5_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_5_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_5_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_5_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_5_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_5_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_5_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_5_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_5_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_5_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_5_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_5_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_5_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_5_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_5_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_5_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_5_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_5_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_5_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_5_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_5_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_5_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_5_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_5_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_5_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_5_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_5_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_5_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_5_io_uop_uopc),
    .io_uop_inst                    (_slots_5_io_uop_inst),
    .io_uop_debug_inst              (_slots_5_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_5_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_5_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_5_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_5_io_uop_fu_code),
    .io_uop_iw_state                (_slots_5_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_5_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_5_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_5_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_5_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_5_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_5_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_5_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_5_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_5_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_5_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_5_io_uop_pc_lob),
    .io_uop_taken                   (_slots_5_io_uop_taken),
    .io_uop_imm_packed              (_slots_5_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_5_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_5_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_5_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_5_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_5_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_5_io_uop_pdst),
    .io_uop_prs1                    (_slots_5_io_uop_prs1),
    .io_uop_prs2                    (_slots_5_io_uop_prs2),
    .io_uop_prs3                    (_slots_5_io_uop_prs3),
    .io_uop_ppred                   (_slots_5_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_5_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_5_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_5_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_5_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_5_io_uop_stale_pdst),
    .io_uop_exception               (_slots_5_io_uop_exception),
    .io_uop_exc_cause               (_slots_5_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_5_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_5_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_5_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_5_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_5_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_5_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_5_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_5_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_5_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_5_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_5_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_5_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_5_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_5_io_uop_ldst),
    .io_uop_lrs1                    (_slots_5_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_5_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_5_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_5_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_5_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_5_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_5_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_5_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_5_io_uop_fp_val),
    .io_uop_fp_single               (_slots_5_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_5_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_5_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_5_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_5_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_5_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_5_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_5_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_6 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_6_io_valid),
    .io_will_be_valid               (_slots_6_io_will_be_valid),
    .io_request                     (_slots_6_io_request),
    .io_grant                       (issue_slots_6_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_5),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_6_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_39 ? _slots_10_io_out_uop_uopc : _GEN_38 ? _slots_9_io_out_uop_uopc : _GEN_37 ? _slots_8_io_out_uop_uopc : _slots_7_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_39 ? _slots_10_io_out_uop_inst : _GEN_38 ? _slots_9_io_out_uop_inst : _GEN_37 ? _slots_8_io_out_uop_inst : _slots_7_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_39 ? _slots_10_io_out_uop_debug_inst : _GEN_38 ? _slots_9_io_out_uop_debug_inst : _GEN_37 ? _slots_8_io_out_uop_debug_inst : _slots_7_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_39 ? _slots_10_io_out_uop_is_rvc : _GEN_38 ? _slots_9_io_out_uop_is_rvc : _GEN_37 ? _slots_8_io_out_uop_is_rvc : _slots_7_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_39 ? _slots_10_io_out_uop_debug_pc : _GEN_38 ? _slots_9_io_out_uop_debug_pc : _GEN_37 ? _slots_8_io_out_uop_debug_pc : _slots_7_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_39 ? _slots_10_io_out_uop_iq_type : _GEN_38 ? _slots_9_io_out_uop_iq_type : _GEN_37 ? _slots_8_io_out_uop_iq_type : _slots_7_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_39 ? _slots_10_io_out_uop_fu_code : _GEN_38 ? _slots_9_io_out_uop_fu_code : _GEN_37 ? _slots_8_io_out_uop_fu_code : _slots_7_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_39 ? _slots_10_io_out_uop_iw_state : _GEN_38 ? _slots_9_io_out_uop_iw_state : _GEN_37 ? _slots_8_io_out_uop_iw_state : _slots_7_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_39 ? _slots_10_io_out_uop_iw_p1_poisoned : _GEN_38 ? _slots_9_io_out_uop_iw_p1_poisoned : _GEN_37 ? _slots_8_io_out_uop_iw_p1_poisoned : _slots_7_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_39 ? _slots_10_io_out_uop_iw_p2_poisoned : _GEN_38 ? _slots_9_io_out_uop_iw_p2_poisoned : _GEN_37 ? _slots_8_io_out_uop_iw_p2_poisoned : _slots_7_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_39 ? _slots_10_io_out_uop_is_br : _GEN_38 ? _slots_9_io_out_uop_is_br : _GEN_37 ? _slots_8_io_out_uop_is_br : _slots_7_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_39 ? _slots_10_io_out_uop_is_jalr : _GEN_38 ? _slots_9_io_out_uop_is_jalr : _GEN_37 ? _slots_8_io_out_uop_is_jalr : _slots_7_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_39 ? _slots_10_io_out_uop_is_jal : _GEN_38 ? _slots_9_io_out_uop_is_jal : _GEN_37 ? _slots_8_io_out_uop_is_jal : _slots_7_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_39 ? _slots_10_io_out_uop_is_sfb : _GEN_38 ? _slots_9_io_out_uop_is_sfb : _GEN_37 ? _slots_8_io_out_uop_is_sfb : _slots_7_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_39 ? _slots_10_io_out_uop_br_mask : _GEN_38 ? _slots_9_io_out_uop_br_mask : _GEN_37 ? _slots_8_io_out_uop_br_mask : _slots_7_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_39 ? _slots_10_io_out_uop_br_tag : _GEN_38 ? _slots_9_io_out_uop_br_tag : _GEN_37 ? _slots_8_io_out_uop_br_tag : _slots_7_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_39 ? _slots_10_io_out_uop_ftq_idx : _GEN_38 ? _slots_9_io_out_uop_ftq_idx : _GEN_37 ? _slots_8_io_out_uop_ftq_idx : _slots_7_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_39 ? _slots_10_io_out_uop_edge_inst : _GEN_38 ? _slots_9_io_out_uop_edge_inst : _GEN_37 ? _slots_8_io_out_uop_edge_inst : _slots_7_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_39 ? _slots_10_io_out_uop_pc_lob : _GEN_38 ? _slots_9_io_out_uop_pc_lob : _GEN_37 ? _slots_8_io_out_uop_pc_lob : _slots_7_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_39 ? _slots_10_io_out_uop_taken : _GEN_38 ? _slots_9_io_out_uop_taken : _GEN_37 ? _slots_8_io_out_uop_taken : _slots_7_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_39 ? _slots_10_io_out_uop_imm_packed : _GEN_38 ? _slots_9_io_out_uop_imm_packed : _GEN_37 ? _slots_8_io_out_uop_imm_packed : _slots_7_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_39 ? _slots_10_io_out_uop_csr_addr : _GEN_38 ? _slots_9_io_out_uop_csr_addr : _GEN_37 ? _slots_8_io_out_uop_csr_addr : _slots_7_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_39 ? _slots_10_io_out_uop_rob_idx : _GEN_38 ? _slots_9_io_out_uop_rob_idx : _GEN_37 ? _slots_8_io_out_uop_rob_idx : _slots_7_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_39 ? _slots_10_io_out_uop_ldq_idx : _GEN_38 ? _slots_9_io_out_uop_ldq_idx : _GEN_37 ? _slots_8_io_out_uop_ldq_idx : _slots_7_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_39 ? _slots_10_io_out_uop_stq_idx : _GEN_38 ? _slots_9_io_out_uop_stq_idx : _GEN_37 ? _slots_8_io_out_uop_stq_idx : _slots_7_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_39 ? _slots_10_io_out_uop_rxq_idx : _GEN_38 ? _slots_9_io_out_uop_rxq_idx : _GEN_37 ? _slots_8_io_out_uop_rxq_idx : _slots_7_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_39 ? _slots_10_io_out_uop_pdst : _GEN_38 ? _slots_9_io_out_uop_pdst : _GEN_37 ? _slots_8_io_out_uop_pdst : _slots_7_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_39 ? _slots_10_io_out_uop_prs1 : _GEN_38 ? _slots_9_io_out_uop_prs1 : _GEN_37 ? _slots_8_io_out_uop_prs1 : _slots_7_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_39 ? _slots_10_io_out_uop_prs2 : _GEN_38 ? _slots_9_io_out_uop_prs2 : _GEN_37 ? _slots_8_io_out_uop_prs2 : _slots_7_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_39 ? _slots_10_io_out_uop_prs3 : _GEN_38 ? _slots_9_io_out_uop_prs3 : _GEN_37 ? _slots_8_io_out_uop_prs3 : _slots_7_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_39 ? _slots_10_io_out_uop_ppred : _GEN_38 ? _slots_9_io_out_uop_ppred : _GEN_37 ? _slots_8_io_out_uop_ppred : _slots_7_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_39 ? _slots_10_io_out_uop_prs1_busy : _GEN_38 ? _slots_9_io_out_uop_prs1_busy : _GEN_37 ? _slots_8_io_out_uop_prs1_busy : _slots_7_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_39 ? _slots_10_io_out_uop_prs2_busy : _GEN_38 ? _slots_9_io_out_uop_prs2_busy : _GEN_37 ? _slots_8_io_out_uop_prs2_busy : _slots_7_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_39 ? _slots_10_io_out_uop_prs3_busy : _GEN_38 ? _slots_9_io_out_uop_prs3_busy : _GEN_37 ? _slots_8_io_out_uop_prs3_busy : _slots_7_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_39 ? _slots_10_io_out_uop_ppred_busy : _GEN_38 ? _slots_9_io_out_uop_ppred_busy : _GEN_37 ? _slots_8_io_out_uop_ppred_busy : _slots_7_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_39 ? _slots_10_io_out_uop_stale_pdst : _GEN_38 ? _slots_9_io_out_uop_stale_pdst : _GEN_37 ? _slots_8_io_out_uop_stale_pdst : _slots_7_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_39 ? _slots_10_io_out_uop_exception : _GEN_38 ? _slots_9_io_out_uop_exception : _GEN_37 ? _slots_8_io_out_uop_exception : _slots_7_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_39 ? _slots_10_io_out_uop_exc_cause : _GEN_38 ? _slots_9_io_out_uop_exc_cause : _GEN_37 ? _slots_8_io_out_uop_exc_cause : _slots_7_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_39 ? _slots_10_io_out_uop_bypassable : _GEN_38 ? _slots_9_io_out_uop_bypassable : _GEN_37 ? _slots_8_io_out_uop_bypassable : _slots_7_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_39 ? _slots_10_io_out_uop_mem_cmd : _GEN_38 ? _slots_9_io_out_uop_mem_cmd : _GEN_37 ? _slots_8_io_out_uop_mem_cmd : _slots_7_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_39 ? _slots_10_io_out_uop_mem_size : _GEN_38 ? _slots_9_io_out_uop_mem_size : _GEN_37 ? _slots_8_io_out_uop_mem_size : _slots_7_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_39 ? _slots_10_io_out_uop_mem_signed : _GEN_38 ? _slots_9_io_out_uop_mem_signed : _GEN_37 ? _slots_8_io_out_uop_mem_signed : _slots_7_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_39 ? _slots_10_io_out_uop_is_fence : _GEN_38 ? _slots_9_io_out_uop_is_fence : _GEN_37 ? _slots_8_io_out_uop_is_fence : _slots_7_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_39 ? _slots_10_io_out_uop_is_fencei : _GEN_38 ? _slots_9_io_out_uop_is_fencei : _GEN_37 ? _slots_8_io_out_uop_is_fencei : _slots_7_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_39 ? _slots_10_io_out_uop_is_amo : _GEN_38 ? _slots_9_io_out_uop_is_amo : _GEN_37 ? _slots_8_io_out_uop_is_amo : _slots_7_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_39 ? _slots_10_io_out_uop_uses_ldq : _GEN_38 ? _slots_9_io_out_uop_uses_ldq : _GEN_37 ? _slots_8_io_out_uop_uses_ldq : _slots_7_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_39 ? _slots_10_io_out_uop_uses_stq : _GEN_38 ? _slots_9_io_out_uop_uses_stq : _GEN_37 ? _slots_8_io_out_uop_uses_stq : _slots_7_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_39 ? _slots_10_io_out_uop_is_sys_pc2epc : _GEN_38 ? _slots_9_io_out_uop_is_sys_pc2epc : _GEN_37 ? _slots_8_io_out_uop_is_sys_pc2epc : _slots_7_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_39 ? _slots_10_io_out_uop_is_unique : _GEN_38 ? _slots_9_io_out_uop_is_unique : _GEN_37 ? _slots_8_io_out_uop_is_unique : _slots_7_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_39 ? _slots_10_io_out_uop_flush_on_commit : _GEN_38 ? _slots_9_io_out_uop_flush_on_commit : _GEN_37 ? _slots_8_io_out_uop_flush_on_commit : _slots_7_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_39 ? _slots_10_io_out_uop_ldst_is_rs1 : _GEN_38 ? _slots_9_io_out_uop_ldst_is_rs1 : _GEN_37 ? _slots_8_io_out_uop_ldst_is_rs1 : _slots_7_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_39 ? _slots_10_io_out_uop_ldst : _GEN_38 ? _slots_9_io_out_uop_ldst : _GEN_37 ? _slots_8_io_out_uop_ldst : _slots_7_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_39 ? _slots_10_io_out_uop_lrs1 : _GEN_38 ? _slots_9_io_out_uop_lrs1 : _GEN_37 ? _slots_8_io_out_uop_lrs1 : _slots_7_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_39 ? _slots_10_io_out_uop_lrs2 : _GEN_38 ? _slots_9_io_out_uop_lrs2 : _GEN_37 ? _slots_8_io_out_uop_lrs2 : _slots_7_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_39 ? _slots_10_io_out_uop_lrs3 : _GEN_38 ? _slots_9_io_out_uop_lrs3 : _GEN_37 ? _slots_8_io_out_uop_lrs3 : _slots_7_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_39 ? _slots_10_io_out_uop_ldst_val : _GEN_38 ? _slots_9_io_out_uop_ldst_val : _GEN_37 ? _slots_8_io_out_uop_ldst_val : _slots_7_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_39 ? _slots_10_io_out_uop_dst_rtype : _GEN_38 ? _slots_9_io_out_uop_dst_rtype : _GEN_37 ? _slots_8_io_out_uop_dst_rtype : _slots_7_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_39 ? _slots_10_io_out_uop_lrs1_rtype : _GEN_38 ? _slots_9_io_out_uop_lrs1_rtype : _GEN_37 ? _slots_8_io_out_uop_lrs1_rtype : _slots_7_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_39 ? _slots_10_io_out_uop_lrs2_rtype : _GEN_38 ? _slots_9_io_out_uop_lrs2_rtype : _GEN_37 ? _slots_8_io_out_uop_lrs2_rtype : _slots_7_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_39 ? _slots_10_io_out_uop_frs3_en : _GEN_38 ? _slots_9_io_out_uop_frs3_en : _GEN_37 ? _slots_8_io_out_uop_frs3_en : _slots_7_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_39 ? _slots_10_io_out_uop_fp_val : _GEN_38 ? _slots_9_io_out_uop_fp_val : _GEN_37 ? _slots_8_io_out_uop_fp_val : _slots_7_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_39 ? _slots_10_io_out_uop_fp_single : _GEN_38 ? _slots_9_io_out_uop_fp_single : _GEN_37 ? _slots_8_io_out_uop_fp_single : _slots_7_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_39 ? _slots_10_io_out_uop_xcpt_pf_if : _GEN_38 ? _slots_9_io_out_uop_xcpt_pf_if : _GEN_37 ? _slots_8_io_out_uop_xcpt_pf_if : _slots_7_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_39 ? _slots_10_io_out_uop_xcpt_ae_if : _GEN_38 ? _slots_9_io_out_uop_xcpt_ae_if : _GEN_37 ? _slots_8_io_out_uop_xcpt_ae_if : _slots_7_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_39 ? _slots_10_io_out_uop_xcpt_ma_if : _GEN_38 ? _slots_9_io_out_uop_xcpt_ma_if : _GEN_37 ? _slots_8_io_out_uop_xcpt_ma_if : _slots_7_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_39 ? _slots_10_io_out_uop_bp_debug_if : _GEN_38 ? _slots_9_io_out_uop_bp_debug_if : _GEN_37 ? _slots_8_io_out_uop_bp_debug_if : _slots_7_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_39 ? _slots_10_io_out_uop_bp_xcpt_if : _GEN_38 ? _slots_9_io_out_uop_bp_xcpt_if : _GEN_37 ? _slots_8_io_out_uop_bp_xcpt_if : _slots_7_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_39 ? _slots_10_io_out_uop_debug_fsrc : _GEN_38 ? _slots_9_io_out_uop_debug_fsrc : _GEN_37 ? _slots_8_io_out_uop_debug_fsrc : _slots_7_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_39 ? _slots_10_io_out_uop_debug_tsrc : _GEN_38 ? _slots_9_io_out_uop_debug_tsrc : _GEN_37 ? _slots_8_io_out_uop_debug_tsrc : _slots_7_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_6_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_6_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_6_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_6_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_6_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_6_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_6_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_6_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_6_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_6_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_6_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_6_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_6_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_6_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_6_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_6_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_6_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_6_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_6_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_6_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_6_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_6_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_6_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_6_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_6_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_6_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_6_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_6_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_6_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_6_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_6_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_6_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_6_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_6_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_6_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_6_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_6_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_6_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_6_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_6_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_6_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_6_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_6_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_6_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_6_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_6_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_6_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_6_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_6_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_6_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_6_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_6_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_6_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_6_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_6_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_6_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_6_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_6_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_6_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_6_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_6_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_6_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_6_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_6_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_6_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_6_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_6_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_6_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_6_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_6_io_uop_uopc),
    .io_uop_inst                    (_slots_6_io_uop_inst),
    .io_uop_debug_inst              (_slots_6_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_6_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_6_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_6_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_6_io_uop_fu_code),
    .io_uop_iw_state                (_slots_6_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_6_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_6_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_6_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_6_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_6_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_6_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_6_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_6_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_6_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_6_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_6_io_uop_pc_lob),
    .io_uop_taken                   (_slots_6_io_uop_taken),
    .io_uop_imm_packed              (_slots_6_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_6_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_6_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_6_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_6_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_6_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_6_io_uop_pdst),
    .io_uop_prs1                    (_slots_6_io_uop_prs1),
    .io_uop_prs2                    (_slots_6_io_uop_prs2),
    .io_uop_prs3                    (_slots_6_io_uop_prs3),
    .io_uop_ppred                   (_slots_6_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_6_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_6_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_6_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_6_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_6_io_uop_stale_pdst),
    .io_uop_exception               (_slots_6_io_uop_exception),
    .io_uop_exc_cause               (_slots_6_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_6_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_6_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_6_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_6_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_6_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_6_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_6_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_6_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_6_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_6_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_6_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_6_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_6_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_6_io_uop_ldst),
    .io_uop_lrs1                    (_slots_6_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_6_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_6_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_6_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_6_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_6_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_6_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_6_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_6_io_uop_fp_val),
    .io_uop_fp_single               (_slots_6_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_6_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_6_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_6_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_6_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_6_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_6_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_6_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_7 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_7_io_valid),
    .io_will_be_valid               (_slots_7_io_will_be_valid),
    .io_request                     (_slots_7_io_request),
    .io_grant                       (issue_slots_7_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_6),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_7_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_42 ? _slots_11_io_out_uop_uopc : _GEN_41 ? _slots_10_io_out_uop_uopc : _GEN_40 ? _slots_9_io_out_uop_uopc : _slots_8_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_42 ? _slots_11_io_out_uop_inst : _GEN_41 ? _slots_10_io_out_uop_inst : _GEN_40 ? _slots_9_io_out_uop_inst : _slots_8_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_42 ? _slots_11_io_out_uop_debug_inst : _GEN_41 ? _slots_10_io_out_uop_debug_inst : _GEN_40 ? _slots_9_io_out_uop_debug_inst : _slots_8_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_42 ? _slots_11_io_out_uop_is_rvc : _GEN_41 ? _slots_10_io_out_uop_is_rvc : _GEN_40 ? _slots_9_io_out_uop_is_rvc : _slots_8_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_42 ? _slots_11_io_out_uop_debug_pc : _GEN_41 ? _slots_10_io_out_uop_debug_pc : _GEN_40 ? _slots_9_io_out_uop_debug_pc : _slots_8_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_42 ? _slots_11_io_out_uop_iq_type : _GEN_41 ? _slots_10_io_out_uop_iq_type : _GEN_40 ? _slots_9_io_out_uop_iq_type : _slots_8_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_42 ? _slots_11_io_out_uop_fu_code : _GEN_41 ? _slots_10_io_out_uop_fu_code : _GEN_40 ? _slots_9_io_out_uop_fu_code : _slots_8_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_42 ? _slots_11_io_out_uop_iw_state : _GEN_41 ? _slots_10_io_out_uop_iw_state : _GEN_40 ? _slots_9_io_out_uop_iw_state : _slots_8_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_42 ? _slots_11_io_out_uop_iw_p1_poisoned : _GEN_41 ? _slots_10_io_out_uop_iw_p1_poisoned : _GEN_40 ? _slots_9_io_out_uop_iw_p1_poisoned : _slots_8_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_42 ? _slots_11_io_out_uop_iw_p2_poisoned : _GEN_41 ? _slots_10_io_out_uop_iw_p2_poisoned : _GEN_40 ? _slots_9_io_out_uop_iw_p2_poisoned : _slots_8_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_42 ? _slots_11_io_out_uop_is_br : _GEN_41 ? _slots_10_io_out_uop_is_br : _GEN_40 ? _slots_9_io_out_uop_is_br : _slots_8_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_42 ? _slots_11_io_out_uop_is_jalr : _GEN_41 ? _slots_10_io_out_uop_is_jalr : _GEN_40 ? _slots_9_io_out_uop_is_jalr : _slots_8_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_42 ? _slots_11_io_out_uop_is_jal : _GEN_41 ? _slots_10_io_out_uop_is_jal : _GEN_40 ? _slots_9_io_out_uop_is_jal : _slots_8_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_42 ? _slots_11_io_out_uop_is_sfb : _GEN_41 ? _slots_10_io_out_uop_is_sfb : _GEN_40 ? _slots_9_io_out_uop_is_sfb : _slots_8_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_42 ? _slots_11_io_out_uop_br_mask : _GEN_41 ? _slots_10_io_out_uop_br_mask : _GEN_40 ? _slots_9_io_out_uop_br_mask : _slots_8_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_42 ? _slots_11_io_out_uop_br_tag : _GEN_41 ? _slots_10_io_out_uop_br_tag : _GEN_40 ? _slots_9_io_out_uop_br_tag : _slots_8_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_42 ? _slots_11_io_out_uop_ftq_idx : _GEN_41 ? _slots_10_io_out_uop_ftq_idx : _GEN_40 ? _slots_9_io_out_uop_ftq_idx : _slots_8_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_42 ? _slots_11_io_out_uop_edge_inst : _GEN_41 ? _slots_10_io_out_uop_edge_inst : _GEN_40 ? _slots_9_io_out_uop_edge_inst : _slots_8_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_42 ? _slots_11_io_out_uop_pc_lob : _GEN_41 ? _slots_10_io_out_uop_pc_lob : _GEN_40 ? _slots_9_io_out_uop_pc_lob : _slots_8_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_42 ? _slots_11_io_out_uop_taken : _GEN_41 ? _slots_10_io_out_uop_taken : _GEN_40 ? _slots_9_io_out_uop_taken : _slots_8_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_42 ? _slots_11_io_out_uop_imm_packed : _GEN_41 ? _slots_10_io_out_uop_imm_packed : _GEN_40 ? _slots_9_io_out_uop_imm_packed : _slots_8_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_42 ? _slots_11_io_out_uop_csr_addr : _GEN_41 ? _slots_10_io_out_uop_csr_addr : _GEN_40 ? _slots_9_io_out_uop_csr_addr : _slots_8_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_42 ? _slots_11_io_out_uop_rob_idx : _GEN_41 ? _slots_10_io_out_uop_rob_idx : _GEN_40 ? _slots_9_io_out_uop_rob_idx : _slots_8_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_42 ? _slots_11_io_out_uop_ldq_idx : _GEN_41 ? _slots_10_io_out_uop_ldq_idx : _GEN_40 ? _slots_9_io_out_uop_ldq_idx : _slots_8_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_42 ? _slots_11_io_out_uop_stq_idx : _GEN_41 ? _slots_10_io_out_uop_stq_idx : _GEN_40 ? _slots_9_io_out_uop_stq_idx : _slots_8_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_42 ? _slots_11_io_out_uop_rxq_idx : _GEN_41 ? _slots_10_io_out_uop_rxq_idx : _GEN_40 ? _slots_9_io_out_uop_rxq_idx : _slots_8_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_42 ? _slots_11_io_out_uop_pdst : _GEN_41 ? _slots_10_io_out_uop_pdst : _GEN_40 ? _slots_9_io_out_uop_pdst : _slots_8_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_42 ? _slots_11_io_out_uop_prs1 : _GEN_41 ? _slots_10_io_out_uop_prs1 : _GEN_40 ? _slots_9_io_out_uop_prs1 : _slots_8_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_42 ? _slots_11_io_out_uop_prs2 : _GEN_41 ? _slots_10_io_out_uop_prs2 : _GEN_40 ? _slots_9_io_out_uop_prs2 : _slots_8_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_42 ? _slots_11_io_out_uop_prs3 : _GEN_41 ? _slots_10_io_out_uop_prs3 : _GEN_40 ? _slots_9_io_out_uop_prs3 : _slots_8_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_42 ? _slots_11_io_out_uop_ppred : _GEN_41 ? _slots_10_io_out_uop_ppred : _GEN_40 ? _slots_9_io_out_uop_ppred : _slots_8_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_42 ? _slots_11_io_out_uop_prs1_busy : _GEN_41 ? _slots_10_io_out_uop_prs1_busy : _GEN_40 ? _slots_9_io_out_uop_prs1_busy : _slots_8_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_42 ? _slots_11_io_out_uop_prs2_busy : _GEN_41 ? _slots_10_io_out_uop_prs2_busy : _GEN_40 ? _slots_9_io_out_uop_prs2_busy : _slots_8_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_42 ? _slots_11_io_out_uop_prs3_busy : _GEN_41 ? _slots_10_io_out_uop_prs3_busy : _GEN_40 ? _slots_9_io_out_uop_prs3_busy : _slots_8_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_42 ? _slots_11_io_out_uop_ppred_busy : _GEN_41 ? _slots_10_io_out_uop_ppred_busy : _GEN_40 ? _slots_9_io_out_uop_ppred_busy : _slots_8_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_42 ? _slots_11_io_out_uop_stale_pdst : _GEN_41 ? _slots_10_io_out_uop_stale_pdst : _GEN_40 ? _slots_9_io_out_uop_stale_pdst : _slots_8_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_42 ? _slots_11_io_out_uop_exception : _GEN_41 ? _slots_10_io_out_uop_exception : _GEN_40 ? _slots_9_io_out_uop_exception : _slots_8_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_42 ? _slots_11_io_out_uop_exc_cause : _GEN_41 ? _slots_10_io_out_uop_exc_cause : _GEN_40 ? _slots_9_io_out_uop_exc_cause : _slots_8_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_42 ? _slots_11_io_out_uop_bypassable : _GEN_41 ? _slots_10_io_out_uop_bypassable : _GEN_40 ? _slots_9_io_out_uop_bypassable : _slots_8_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_42 ? _slots_11_io_out_uop_mem_cmd : _GEN_41 ? _slots_10_io_out_uop_mem_cmd : _GEN_40 ? _slots_9_io_out_uop_mem_cmd : _slots_8_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_42 ? _slots_11_io_out_uop_mem_size : _GEN_41 ? _slots_10_io_out_uop_mem_size : _GEN_40 ? _slots_9_io_out_uop_mem_size : _slots_8_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_42 ? _slots_11_io_out_uop_mem_signed : _GEN_41 ? _slots_10_io_out_uop_mem_signed : _GEN_40 ? _slots_9_io_out_uop_mem_signed : _slots_8_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_42 ? _slots_11_io_out_uop_is_fence : _GEN_41 ? _slots_10_io_out_uop_is_fence : _GEN_40 ? _slots_9_io_out_uop_is_fence : _slots_8_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_42 ? _slots_11_io_out_uop_is_fencei : _GEN_41 ? _slots_10_io_out_uop_is_fencei : _GEN_40 ? _slots_9_io_out_uop_is_fencei : _slots_8_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_42 ? _slots_11_io_out_uop_is_amo : _GEN_41 ? _slots_10_io_out_uop_is_amo : _GEN_40 ? _slots_9_io_out_uop_is_amo : _slots_8_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_42 ? _slots_11_io_out_uop_uses_ldq : _GEN_41 ? _slots_10_io_out_uop_uses_ldq : _GEN_40 ? _slots_9_io_out_uop_uses_ldq : _slots_8_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_42 ? _slots_11_io_out_uop_uses_stq : _GEN_41 ? _slots_10_io_out_uop_uses_stq : _GEN_40 ? _slots_9_io_out_uop_uses_stq : _slots_8_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_42 ? _slots_11_io_out_uop_is_sys_pc2epc : _GEN_41 ? _slots_10_io_out_uop_is_sys_pc2epc : _GEN_40 ? _slots_9_io_out_uop_is_sys_pc2epc : _slots_8_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_42 ? _slots_11_io_out_uop_is_unique : _GEN_41 ? _slots_10_io_out_uop_is_unique : _GEN_40 ? _slots_9_io_out_uop_is_unique : _slots_8_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_42 ? _slots_11_io_out_uop_flush_on_commit : _GEN_41 ? _slots_10_io_out_uop_flush_on_commit : _GEN_40 ? _slots_9_io_out_uop_flush_on_commit : _slots_8_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_42 ? _slots_11_io_out_uop_ldst_is_rs1 : _GEN_41 ? _slots_10_io_out_uop_ldst_is_rs1 : _GEN_40 ? _slots_9_io_out_uop_ldst_is_rs1 : _slots_8_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_42 ? _slots_11_io_out_uop_ldst : _GEN_41 ? _slots_10_io_out_uop_ldst : _GEN_40 ? _slots_9_io_out_uop_ldst : _slots_8_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_42 ? _slots_11_io_out_uop_lrs1 : _GEN_41 ? _slots_10_io_out_uop_lrs1 : _GEN_40 ? _slots_9_io_out_uop_lrs1 : _slots_8_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_42 ? _slots_11_io_out_uop_lrs2 : _GEN_41 ? _slots_10_io_out_uop_lrs2 : _GEN_40 ? _slots_9_io_out_uop_lrs2 : _slots_8_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_42 ? _slots_11_io_out_uop_lrs3 : _GEN_41 ? _slots_10_io_out_uop_lrs3 : _GEN_40 ? _slots_9_io_out_uop_lrs3 : _slots_8_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_42 ? _slots_11_io_out_uop_ldst_val : _GEN_41 ? _slots_10_io_out_uop_ldst_val : _GEN_40 ? _slots_9_io_out_uop_ldst_val : _slots_8_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_42 ? _slots_11_io_out_uop_dst_rtype : _GEN_41 ? _slots_10_io_out_uop_dst_rtype : _GEN_40 ? _slots_9_io_out_uop_dst_rtype : _slots_8_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_42 ? _slots_11_io_out_uop_lrs1_rtype : _GEN_41 ? _slots_10_io_out_uop_lrs1_rtype : _GEN_40 ? _slots_9_io_out_uop_lrs1_rtype : _slots_8_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_42 ? _slots_11_io_out_uop_lrs2_rtype : _GEN_41 ? _slots_10_io_out_uop_lrs2_rtype : _GEN_40 ? _slots_9_io_out_uop_lrs2_rtype : _slots_8_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_42 ? _slots_11_io_out_uop_frs3_en : _GEN_41 ? _slots_10_io_out_uop_frs3_en : _GEN_40 ? _slots_9_io_out_uop_frs3_en : _slots_8_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_42 ? _slots_11_io_out_uop_fp_val : _GEN_41 ? _slots_10_io_out_uop_fp_val : _GEN_40 ? _slots_9_io_out_uop_fp_val : _slots_8_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_42 ? _slots_11_io_out_uop_fp_single : _GEN_41 ? _slots_10_io_out_uop_fp_single : _GEN_40 ? _slots_9_io_out_uop_fp_single : _slots_8_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_42 ? _slots_11_io_out_uop_xcpt_pf_if : _GEN_41 ? _slots_10_io_out_uop_xcpt_pf_if : _GEN_40 ? _slots_9_io_out_uop_xcpt_pf_if : _slots_8_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_42 ? _slots_11_io_out_uop_xcpt_ae_if : _GEN_41 ? _slots_10_io_out_uop_xcpt_ae_if : _GEN_40 ? _slots_9_io_out_uop_xcpt_ae_if : _slots_8_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_42 ? _slots_11_io_out_uop_xcpt_ma_if : _GEN_41 ? _slots_10_io_out_uop_xcpt_ma_if : _GEN_40 ? _slots_9_io_out_uop_xcpt_ma_if : _slots_8_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_42 ? _slots_11_io_out_uop_bp_debug_if : _GEN_41 ? _slots_10_io_out_uop_bp_debug_if : _GEN_40 ? _slots_9_io_out_uop_bp_debug_if : _slots_8_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_42 ? _slots_11_io_out_uop_bp_xcpt_if : _GEN_41 ? _slots_10_io_out_uop_bp_xcpt_if : _GEN_40 ? _slots_9_io_out_uop_bp_xcpt_if : _slots_8_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_42 ? _slots_11_io_out_uop_debug_fsrc : _GEN_41 ? _slots_10_io_out_uop_debug_fsrc : _GEN_40 ? _slots_9_io_out_uop_debug_fsrc : _slots_8_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_42 ? _slots_11_io_out_uop_debug_tsrc : _GEN_41 ? _slots_10_io_out_uop_debug_tsrc : _GEN_40 ? _slots_9_io_out_uop_debug_tsrc : _slots_8_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_7_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_7_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_7_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_7_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_7_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_7_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_7_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_7_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_7_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_7_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_7_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_7_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_7_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_7_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_7_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_7_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_7_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_7_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_7_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_7_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_7_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_7_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_7_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_7_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_7_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_7_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_7_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_7_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_7_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_7_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_7_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_7_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_7_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_7_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_7_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_7_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_7_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_7_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_7_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_7_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_7_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_7_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_7_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_7_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_7_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_7_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_7_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_7_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_7_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_7_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_7_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_7_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_7_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_7_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_7_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_7_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_7_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_7_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_7_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_7_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_7_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_7_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_7_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_7_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_7_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_7_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_7_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_7_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_7_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_7_io_uop_uopc),
    .io_uop_inst                    (_slots_7_io_uop_inst),
    .io_uop_debug_inst              (_slots_7_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_7_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_7_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_7_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_7_io_uop_fu_code),
    .io_uop_iw_state                (_slots_7_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_7_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_7_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_7_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_7_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_7_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_7_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_7_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_7_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_7_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_7_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_7_io_uop_pc_lob),
    .io_uop_taken                   (_slots_7_io_uop_taken),
    .io_uop_imm_packed              (_slots_7_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_7_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_7_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_7_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_7_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_7_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_7_io_uop_pdst),
    .io_uop_prs1                    (_slots_7_io_uop_prs1),
    .io_uop_prs2                    (_slots_7_io_uop_prs2),
    .io_uop_prs3                    (_slots_7_io_uop_prs3),
    .io_uop_ppred                   (_slots_7_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_7_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_7_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_7_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_7_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_7_io_uop_stale_pdst),
    .io_uop_exception               (_slots_7_io_uop_exception),
    .io_uop_exc_cause               (_slots_7_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_7_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_7_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_7_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_7_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_7_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_7_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_7_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_7_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_7_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_7_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_7_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_7_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_7_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_7_io_uop_ldst),
    .io_uop_lrs1                    (_slots_7_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_7_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_7_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_7_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_7_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_7_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_7_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_7_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_7_io_uop_fp_val),
    .io_uop_fp_single               (_slots_7_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_7_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_7_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_7_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_7_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_7_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_7_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_7_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_8 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_8_io_valid),
    .io_will_be_valid               (_slots_8_io_will_be_valid),
    .io_request                     (_slots_8_io_request),
    .io_grant                       (issue_slots_8_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_7),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_8_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_45 ? _slots_12_io_out_uop_uopc : _GEN_44 ? _slots_11_io_out_uop_uopc : _GEN_43 ? _slots_10_io_out_uop_uopc : _slots_9_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_45 ? _slots_12_io_out_uop_inst : _GEN_44 ? _slots_11_io_out_uop_inst : _GEN_43 ? _slots_10_io_out_uop_inst : _slots_9_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_45 ? _slots_12_io_out_uop_debug_inst : _GEN_44 ? _slots_11_io_out_uop_debug_inst : _GEN_43 ? _slots_10_io_out_uop_debug_inst : _slots_9_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_45 ? _slots_12_io_out_uop_is_rvc : _GEN_44 ? _slots_11_io_out_uop_is_rvc : _GEN_43 ? _slots_10_io_out_uop_is_rvc : _slots_9_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_45 ? _slots_12_io_out_uop_debug_pc : _GEN_44 ? _slots_11_io_out_uop_debug_pc : _GEN_43 ? _slots_10_io_out_uop_debug_pc : _slots_9_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_45 ? _slots_12_io_out_uop_iq_type : _GEN_44 ? _slots_11_io_out_uop_iq_type : _GEN_43 ? _slots_10_io_out_uop_iq_type : _slots_9_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_45 ? _slots_12_io_out_uop_fu_code : _GEN_44 ? _slots_11_io_out_uop_fu_code : _GEN_43 ? _slots_10_io_out_uop_fu_code : _slots_9_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_45 ? _slots_12_io_out_uop_iw_state : _GEN_44 ? _slots_11_io_out_uop_iw_state : _GEN_43 ? _slots_10_io_out_uop_iw_state : _slots_9_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_45 ? _slots_12_io_out_uop_iw_p1_poisoned : _GEN_44 ? _slots_11_io_out_uop_iw_p1_poisoned : _GEN_43 ? _slots_10_io_out_uop_iw_p1_poisoned : _slots_9_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_45 ? _slots_12_io_out_uop_iw_p2_poisoned : _GEN_44 ? _slots_11_io_out_uop_iw_p2_poisoned : _GEN_43 ? _slots_10_io_out_uop_iw_p2_poisoned : _slots_9_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_45 ? _slots_12_io_out_uop_is_br : _GEN_44 ? _slots_11_io_out_uop_is_br : _GEN_43 ? _slots_10_io_out_uop_is_br : _slots_9_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_45 ? _slots_12_io_out_uop_is_jalr : _GEN_44 ? _slots_11_io_out_uop_is_jalr : _GEN_43 ? _slots_10_io_out_uop_is_jalr : _slots_9_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_45 ? _slots_12_io_out_uop_is_jal : _GEN_44 ? _slots_11_io_out_uop_is_jal : _GEN_43 ? _slots_10_io_out_uop_is_jal : _slots_9_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_45 ? _slots_12_io_out_uop_is_sfb : _GEN_44 ? _slots_11_io_out_uop_is_sfb : _GEN_43 ? _slots_10_io_out_uop_is_sfb : _slots_9_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_45 ? _slots_12_io_out_uop_br_mask : _GEN_44 ? _slots_11_io_out_uop_br_mask : _GEN_43 ? _slots_10_io_out_uop_br_mask : _slots_9_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_45 ? _slots_12_io_out_uop_br_tag : _GEN_44 ? _slots_11_io_out_uop_br_tag : _GEN_43 ? _slots_10_io_out_uop_br_tag : _slots_9_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_45 ? _slots_12_io_out_uop_ftq_idx : _GEN_44 ? _slots_11_io_out_uop_ftq_idx : _GEN_43 ? _slots_10_io_out_uop_ftq_idx : _slots_9_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_45 ? _slots_12_io_out_uop_edge_inst : _GEN_44 ? _slots_11_io_out_uop_edge_inst : _GEN_43 ? _slots_10_io_out_uop_edge_inst : _slots_9_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_45 ? _slots_12_io_out_uop_pc_lob : _GEN_44 ? _slots_11_io_out_uop_pc_lob : _GEN_43 ? _slots_10_io_out_uop_pc_lob : _slots_9_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_45 ? _slots_12_io_out_uop_taken : _GEN_44 ? _slots_11_io_out_uop_taken : _GEN_43 ? _slots_10_io_out_uop_taken : _slots_9_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_45 ? _slots_12_io_out_uop_imm_packed : _GEN_44 ? _slots_11_io_out_uop_imm_packed : _GEN_43 ? _slots_10_io_out_uop_imm_packed : _slots_9_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_45 ? _slots_12_io_out_uop_csr_addr : _GEN_44 ? _slots_11_io_out_uop_csr_addr : _GEN_43 ? _slots_10_io_out_uop_csr_addr : _slots_9_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_45 ? _slots_12_io_out_uop_rob_idx : _GEN_44 ? _slots_11_io_out_uop_rob_idx : _GEN_43 ? _slots_10_io_out_uop_rob_idx : _slots_9_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_45 ? _slots_12_io_out_uop_ldq_idx : _GEN_44 ? _slots_11_io_out_uop_ldq_idx : _GEN_43 ? _slots_10_io_out_uop_ldq_idx : _slots_9_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_45 ? _slots_12_io_out_uop_stq_idx : _GEN_44 ? _slots_11_io_out_uop_stq_idx : _GEN_43 ? _slots_10_io_out_uop_stq_idx : _slots_9_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_45 ? _slots_12_io_out_uop_rxq_idx : _GEN_44 ? _slots_11_io_out_uop_rxq_idx : _GEN_43 ? _slots_10_io_out_uop_rxq_idx : _slots_9_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_45 ? _slots_12_io_out_uop_pdst : _GEN_44 ? _slots_11_io_out_uop_pdst : _GEN_43 ? _slots_10_io_out_uop_pdst : _slots_9_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_45 ? _slots_12_io_out_uop_prs1 : _GEN_44 ? _slots_11_io_out_uop_prs1 : _GEN_43 ? _slots_10_io_out_uop_prs1 : _slots_9_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_45 ? _slots_12_io_out_uop_prs2 : _GEN_44 ? _slots_11_io_out_uop_prs2 : _GEN_43 ? _slots_10_io_out_uop_prs2 : _slots_9_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_45 ? _slots_12_io_out_uop_prs3 : _GEN_44 ? _slots_11_io_out_uop_prs3 : _GEN_43 ? _slots_10_io_out_uop_prs3 : _slots_9_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_45 ? _slots_12_io_out_uop_ppred : _GEN_44 ? _slots_11_io_out_uop_ppred : _GEN_43 ? _slots_10_io_out_uop_ppred : _slots_9_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_45 ? _slots_12_io_out_uop_prs1_busy : _GEN_44 ? _slots_11_io_out_uop_prs1_busy : _GEN_43 ? _slots_10_io_out_uop_prs1_busy : _slots_9_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_45 ? _slots_12_io_out_uop_prs2_busy : _GEN_44 ? _slots_11_io_out_uop_prs2_busy : _GEN_43 ? _slots_10_io_out_uop_prs2_busy : _slots_9_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_45 ? _slots_12_io_out_uop_prs3_busy : _GEN_44 ? _slots_11_io_out_uop_prs3_busy : _GEN_43 ? _slots_10_io_out_uop_prs3_busy : _slots_9_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_45 ? _slots_12_io_out_uop_ppred_busy : _GEN_44 ? _slots_11_io_out_uop_ppred_busy : _GEN_43 ? _slots_10_io_out_uop_ppred_busy : _slots_9_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_45 ? _slots_12_io_out_uop_stale_pdst : _GEN_44 ? _slots_11_io_out_uop_stale_pdst : _GEN_43 ? _slots_10_io_out_uop_stale_pdst : _slots_9_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_45 ? _slots_12_io_out_uop_exception : _GEN_44 ? _slots_11_io_out_uop_exception : _GEN_43 ? _slots_10_io_out_uop_exception : _slots_9_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_45 ? _slots_12_io_out_uop_exc_cause : _GEN_44 ? _slots_11_io_out_uop_exc_cause : _GEN_43 ? _slots_10_io_out_uop_exc_cause : _slots_9_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_45 ? _slots_12_io_out_uop_bypassable : _GEN_44 ? _slots_11_io_out_uop_bypassable : _GEN_43 ? _slots_10_io_out_uop_bypassable : _slots_9_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_45 ? _slots_12_io_out_uop_mem_cmd : _GEN_44 ? _slots_11_io_out_uop_mem_cmd : _GEN_43 ? _slots_10_io_out_uop_mem_cmd : _slots_9_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_45 ? _slots_12_io_out_uop_mem_size : _GEN_44 ? _slots_11_io_out_uop_mem_size : _GEN_43 ? _slots_10_io_out_uop_mem_size : _slots_9_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_45 ? _slots_12_io_out_uop_mem_signed : _GEN_44 ? _slots_11_io_out_uop_mem_signed : _GEN_43 ? _slots_10_io_out_uop_mem_signed : _slots_9_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_45 ? _slots_12_io_out_uop_is_fence : _GEN_44 ? _slots_11_io_out_uop_is_fence : _GEN_43 ? _slots_10_io_out_uop_is_fence : _slots_9_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_45 ? _slots_12_io_out_uop_is_fencei : _GEN_44 ? _slots_11_io_out_uop_is_fencei : _GEN_43 ? _slots_10_io_out_uop_is_fencei : _slots_9_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_45 ? _slots_12_io_out_uop_is_amo : _GEN_44 ? _slots_11_io_out_uop_is_amo : _GEN_43 ? _slots_10_io_out_uop_is_amo : _slots_9_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_45 ? _slots_12_io_out_uop_uses_ldq : _GEN_44 ? _slots_11_io_out_uop_uses_ldq : _GEN_43 ? _slots_10_io_out_uop_uses_ldq : _slots_9_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_45 ? _slots_12_io_out_uop_uses_stq : _GEN_44 ? _slots_11_io_out_uop_uses_stq : _GEN_43 ? _slots_10_io_out_uop_uses_stq : _slots_9_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_45 ? _slots_12_io_out_uop_is_sys_pc2epc : _GEN_44 ? _slots_11_io_out_uop_is_sys_pc2epc : _GEN_43 ? _slots_10_io_out_uop_is_sys_pc2epc : _slots_9_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_45 ? _slots_12_io_out_uop_is_unique : _GEN_44 ? _slots_11_io_out_uop_is_unique : _GEN_43 ? _slots_10_io_out_uop_is_unique : _slots_9_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_45 ? _slots_12_io_out_uop_flush_on_commit : _GEN_44 ? _slots_11_io_out_uop_flush_on_commit : _GEN_43 ? _slots_10_io_out_uop_flush_on_commit : _slots_9_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_45 ? _slots_12_io_out_uop_ldst_is_rs1 : _GEN_44 ? _slots_11_io_out_uop_ldst_is_rs1 : _GEN_43 ? _slots_10_io_out_uop_ldst_is_rs1 : _slots_9_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_45 ? _slots_12_io_out_uop_ldst : _GEN_44 ? _slots_11_io_out_uop_ldst : _GEN_43 ? _slots_10_io_out_uop_ldst : _slots_9_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_45 ? _slots_12_io_out_uop_lrs1 : _GEN_44 ? _slots_11_io_out_uop_lrs1 : _GEN_43 ? _slots_10_io_out_uop_lrs1 : _slots_9_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_45 ? _slots_12_io_out_uop_lrs2 : _GEN_44 ? _slots_11_io_out_uop_lrs2 : _GEN_43 ? _slots_10_io_out_uop_lrs2 : _slots_9_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_45 ? _slots_12_io_out_uop_lrs3 : _GEN_44 ? _slots_11_io_out_uop_lrs3 : _GEN_43 ? _slots_10_io_out_uop_lrs3 : _slots_9_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_45 ? _slots_12_io_out_uop_ldst_val : _GEN_44 ? _slots_11_io_out_uop_ldst_val : _GEN_43 ? _slots_10_io_out_uop_ldst_val : _slots_9_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_45 ? _slots_12_io_out_uop_dst_rtype : _GEN_44 ? _slots_11_io_out_uop_dst_rtype : _GEN_43 ? _slots_10_io_out_uop_dst_rtype : _slots_9_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_45 ? _slots_12_io_out_uop_lrs1_rtype : _GEN_44 ? _slots_11_io_out_uop_lrs1_rtype : _GEN_43 ? _slots_10_io_out_uop_lrs1_rtype : _slots_9_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_45 ? _slots_12_io_out_uop_lrs2_rtype : _GEN_44 ? _slots_11_io_out_uop_lrs2_rtype : _GEN_43 ? _slots_10_io_out_uop_lrs2_rtype : _slots_9_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_45 ? _slots_12_io_out_uop_frs3_en : _GEN_44 ? _slots_11_io_out_uop_frs3_en : _GEN_43 ? _slots_10_io_out_uop_frs3_en : _slots_9_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_45 ? _slots_12_io_out_uop_fp_val : _GEN_44 ? _slots_11_io_out_uop_fp_val : _GEN_43 ? _slots_10_io_out_uop_fp_val : _slots_9_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_45 ? _slots_12_io_out_uop_fp_single : _GEN_44 ? _slots_11_io_out_uop_fp_single : _GEN_43 ? _slots_10_io_out_uop_fp_single : _slots_9_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_45 ? _slots_12_io_out_uop_xcpt_pf_if : _GEN_44 ? _slots_11_io_out_uop_xcpt_pf_if : _GEN_43 ? _slots_10_io_out_uop_xcpt_pf_if : _slots_9_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_45 ? _slots_12_io_out_uop_xcpt_ae_if : _GEN_44 ? _slots_11_io_out_uop_xcpt_ae_if : _GEN_43 ? _slots_10_io_out_uop_xcpt_ae_if : _slots_9_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_45 ? _slots_12_io_out_uop_xcpt_ma_if : _GEN_44 ? _slots_11_io_out_uop_xcpt_ma_if : _GEN_43 ? _slots_10_io_out_uop_xcpt_ma_if : _slots_9_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_45 ? _slots_12_io_out_uop_bp_debug_if : _GEN_44 ? _slots_11_io_out_uop_bp_debug_if : _GEN_43 ? _slots_10_io_out_uop_bp_debug_if : _slots_9_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_45 ? _slots_12_io_out_uop_bp_xcpt_if : _GEN_44 ? _slots_11_io_out_uop_bp_xcpt_if : _GEN_43 ? _slots_10_io_out_uop_bp_xcpt_if : _slots_9_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_45 ? _slots_12_io_out_uop_debug_fsrc : _GEN_44 ? _slots_11_io_out_uop_debug_fsrc : _GEN_43 ? _slots_10_io_out_uop_debug_fsrc : _slots_9_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_45 ? _slots_12_io_out_uop_debug_tsrc : _GEN_44 ? _slots_11_io_out_uop_debug_tsrc : _GEN_43 ? _slots_10_io_out_uop_debug_tsrc : _slots_9_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_8_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_8_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_8_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_8_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_8_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_8_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_8_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_8_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_8_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_8_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_8_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_8_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_8_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_8_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_8_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_8_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_8_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_8_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_8_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_8_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_8_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_8_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_8_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_8_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_8_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_8_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_8_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_8_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_8_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_8_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_8_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_8_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_8_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_8_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_8_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_8_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_8_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_8_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_8_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_8_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_8_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_8_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_8_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_8_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_8_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_8_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_8_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_8_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_8_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_8_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_8_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_8_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_8_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_8_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_8_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_8_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_8_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_8_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_8_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_8_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_8_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_8_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_8_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_8_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_8_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_8_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_8_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_8_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_8_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_8_io_uop_uopc),
    .io_uop_inst                    (_slots_8_io_uop_inst),
    .io_uop_debug_inst              (_slots_8_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_8_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_8_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_8_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_8_io_uop_fu_code),
    .io_uop_iw_state                (_slots_8_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_8_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_8_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_8_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_8_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_8_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_8_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_8_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_8_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_8_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_8_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_8_io_uop_pc_lob),
    .io_uop_taken                   (_slots_8_io_uop_taken),
    .io_uop_imm_packed              (_slots_8_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_8_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_8_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_8_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_8_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_8_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_8_io_uop_pdst),
    .io_uop_prs1                    (_slots_8_io_uop_prs1),
    .io_uop_prs2                    (_slots_8_io_uop_prs2),
    .io_uop_prs3                    (_slots_8_io_uop_prs3),
    .io_uop_ppred                   (_slots_8_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_8_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_8_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_8_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_8_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_8_io_uop_stale_pdst),
    .io_uop_exception               (_slots_8_io_uop_exception),
    .io_uop_exc_cause               (_slots_8_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_8_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_8_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_8_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_8_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_8_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_8_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_8_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_8_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_8_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_8_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_8_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_8_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_8_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_8_io_uop_ldst),
    .io_uop_lrs1                    (_slots_8_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_8_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_8_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_8_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_8_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_8_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_8_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_8_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_8_io_uop_fp_val),
    .io_uop_fp_single               (_slots_8_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_8_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_8_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_8_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_8_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_8_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_8_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_8_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_9 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_9_io_valid),
    .io_will_be_valid               (_slots_9_io_will_be_valid),
    .io_request                     (_slots_9_io_request),
    .io_grant                       (issue_slots_9_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_8),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_9_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_48 ? _slots_13_io_out_uop_uopc : _GEN_47 ? _slots_12_io_out_uop_uopc : _GEN_46 ? _slots_11_io_out_uop_uopc : _slots_10_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_48 ? _slots_13_io_out_uop_inst : _GEN_47 ? _slots_12_io_out_uop_inst : _GEN_46 ? _slots_11_io_out_uop_inst : _slots_10_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_48 ? _slots_13_io_out_uop_debug_inst : _GEN_47 ? _slots_12_io_out_uop_debug_inst : _GEN_46 ? _slots_11_io_out_uop_debug_inst : _slots_10_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_48 ? _slots_13_io_out_uop_is_rvc : _GEN_47 ? _slots_12_io_out_uop_is_rvc : _GEN_46 ? _slots_11_io_out_uop_is_rvc : _slots_10_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_48 ? _slots_13_io_out_uop_debug_pc : _GEN_47 ? _slots_12_io_out_uop_debug_pc : _GEN_46 ? _slots_11_io_out_uop_debug_pc : _slots_10_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_48 ? _slots_13_io_out_uop_iq_type : _GEN_47 ? _slots_12_io_out_uop_iq_type : _GEN_46 ? _slots_11_io_out_uop_iq_type : _slots_10_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_48 ? _slots_13_io_out_uop_fu_code : _GEN_47 ? _slots_12_io_out_uop_fu_code : _GEN_46 ? _slots_11_io_out_uop_fu_code : _slots_10_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_48 ? _slots_13_io_out_uop_iw_state : _GEN_47 ? _slots_12_io_out_uop_iw_state : _GEN_46 ? _slots_11_io_out_uop_iw_state : _slots_10_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_48 ? _slots_13_io_out_uop_iw_p1_poisoned : _GEN_47 ? _slots_12_io_out_uop_iw_p1_poisoned : _GEN_46 ? _slots_11_io_out_uop_iw_p1_poisoned : _slots_10_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_48 ? _slots_13_io_out_uop_iw_p2_poisoned : _GEN_47 ? _slots_12_io_out_uop_iw_p2_poisoned : _GEN_46 ? _slots_11_io_out_uop_iw_p2_poisoned : _slots_10_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_48 ? _slots_13_io_out_uop_is_br : _GEN_47 ? _slots_12_io_out_uop_is_br : _GEN_46 ? _slots_11_io_out_uop_is_br : _slots_10_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_48 ? _slots_13_io_out_uop_is_jalr : _GEN_47 ? _slots_12_io_out_uop_is_jalr : _GEN_46 ? _slots_11_io_out_uop_is_jalr : _slots_10_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_48 ? _slots_13_io_out_uop_is_jal : _GEN_47 ? _slots_12_io_out_uop_is_jal : _GEN_46 ? _slots_11_io_out_uop_is_jal : _slots_10_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_48 ? _slots_13_io_out_uop_is_sfb : _GEN_47 ? _slots_12_io_out_uop_is_sfb : _GEN_46 ? _slots_11_io_out_uop_is_sfb : _slots_10_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_48 ? _slots_13_io_out_uop_br_mask : _GEN_47 ? _slots_12_io_out_uop_br_mask : _GEN_46 ? _slots_11_io_out_uop_br_mask : _slots_10_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_48 ? _slots_13_io_out_uop_br_tag : _GEN_47 ? _slots_12_io_out_uop_br_tag : _GEN_46 ? _slots_11_io_out_uop_br_tag : _slots_10_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_48 ? _slots_13_io_out_uop_ftq_idx : _GEN_47 ? _slots_12_io_out_uop_ftq_idx : _GEN_46 ? _slots_11_io_out_uop_ftq_idx : _slots_10_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_48 ? _slots_13_io_out_uop_edge_inst : _GEN_47 ? _slots_12_io_out_uop_edge_inst : _GEN_46 ? _slots_11_io_out_uop_edge_inst : _slots_10_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_48 ? _slots_13_io_out_uop_pc_lob : _GEN_47 ? _slots_12_io_out_uop_pc_lob : _GEN_46 ? _slots_11_io_out_uop_pc_lob : _slots_10_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_48 ? _slots_13_io_out_uop_taken : _GEN_47 ? _slots_12_io_out_uop_taken : _GEN_46 ? _slots_11_io_out_uop_taken : _slots_10_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_48 ? _slots_13_io_out_uop_imm_packed : _GEN_47 ? _slots_12_io_out_uop_imm_packed : _GEN_46 ? _slots_11_io_out_uop_imm_packed : _slots_10_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_48 ? _slots_13_io_out_uop_csr_addr : _GEN_47 ? _slots_12_io_out_uop_csr_addr : _GEN_46 ? _slots_11_io_out_uop_csr_addr : _slots_10_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_48 ? _slots_13_io_out_uop_rob_idx : _GEN_47 ? _slots_12_io_out_uop_rob_idx : _GEN_46 ? _slots_11_io_out_uop_rob_idx : _slots_10_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_48 ? _slots_13_io_out_uop_ldq_idx : _GEN_47 ? _slots_12_io_out_uop_ldq_idx : _GEN_46 ? _slots_11_io_out_uop_ldq_idx : _slots_10_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_48 ? _slots_13_io_out_uop_stq_idx : _GEN_47 ? _slots_12_io_out_uop_stq_idx : _GEN_46 ? _slots_11_io_out_uop_stq_idx : _slots_10_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_48 ? _slots_13_io_out_uop_rxq_idx : _GEN_47 ? _slots_12_io_out_uop_rxq_idx : _GEN_46 ? _slots_11_io_out_uop_rxq_idx : _slots_10_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_48 ? _slots_13_io_out_uop_pdst : _GEN_47 ? _slots_12_io_out_uop_pdst : _GEN_46 ? _slots_11_io_out_uop_pdst : _slots_10_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_48 ? _slots_13_io_out_uop_prs1 : _GEN_47 ? _slots_12_io_out_uop_prs1 : _GEN_46 ? _slots_11_io_out_uop_prs1 : _slots_10_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_48 ? _slots_13_io_out_uop_prs2 : _GEN_47 ? _slots_12_io_out_uop_prs2 : _GEN_46 ? _slots_11_io_out_uop_prs2 : _slots_10_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_48 ? _slots_13_io_out_uop_prs3 : _GEN_47 ? _slots_12_io_out_uop_prs3 : _GEN_46 ? _slots_11_io_out_uop_prs3 : _slots_10_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_48 ? _slots_13_io_out_uop_ppred : _GEN_47 ? _slots_12_io_out_uop_ppred : _GEN_46 ? _slots_11_io_out_uop_ppred : _slots_10_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_48 ? _slots_13_io_out_uop_prs1_busy : _GEN_47 ? _slots_12_io_out_uop_prs1_busy : _GEN_46 ? _slots_11_io_out_uop_prs1_busy : _slots_10_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_48 ? _slots_13_io_out_uop_prs2_busy : _GEN_47 ? _slots_12_io_out_uop_prs2_busy : _GEN_46 ? _slots_11_io_out_uop_prs2_busy : _slots_10_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_48 ? _slots_13_io_out_uop_prs3_busy : _GEN_47 ? _slots_12_io_out_uop_prs3_busy : _GEN_46 ? _slots_11_io_out_uop_prs3_busy : _slots_10_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_48 ? _slots_13_io_out_uop_ppred_busy : _GEN_47 ? _slots_12_io_out_uop_ppred_busy : _GEN_46 ? _slots_11_io_out_uop_ppred_busy : _slots_10_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_48 ? _slots_13_io_out_uop_stale_pdst : _GEN_47 ? _slots_12_io_out_uop_stale_pdst : _GEN_46 ? _slots_11_io_out_uop_stale_pdst : _slots_10_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_48 ? _slots_13_io_out_uop_exception : _GEN_47 ? _slots_12_io_out_uop_exception : _GEN_46 ? _slots_11_io_out_uop_exception : _slots_10_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_48 ? _slots_13_io_out_uop_exc_cause : _GEN_47 ? _slots_12_io_out_uop_exc_cause : _GEN_46 ? _slots_11_io_out_uop_exc_cause : _slots_10_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_48 ? _slots_13_io_out_uop_bypassable : _GEN_47 ? _slots_12_io_out_uop_bypassable : _GEN_46 ? _slots_11_io_out_uop_bypassable : _slots_10_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_48 ? _slots_13_io_out_uop_mem_cmd : _GEN_47 ? _slots_12_io_out_uop_mem_cmd : _GEN_46 ? _slots_11_io_out_uop_mem_cmd : _slots_10_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_48 ? _slots_13_io_out_uop_mem_size : _GEN_47 ? _slots_12_io_out_uop_mem_size : _GEN_46 ? _slots_11_io_out_uop_mem_size : _slots_10_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_48 ? _slots_13_io_out_uop_mem_signed : _GEN_47 ? _slots_12_io_out_uop_mem_signed : _GEN_46 ? _slots_11_io_out_uop_mem_signed : _slots_10_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_48 ? _slots_13_io_out_uop_is_fence : _GEN_47 ? _slots_12_io_out_uop_is_fence : _GEN_46 ? _slots_11_io_out_uop_is_fence : _slots_10_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_48 ? _slots_13_io_out_uop_is_fencei : _GEN_47 ? _slots_12_io_out_uop_is_fencei : _GEN_46 ? _slots_11_io_out_uop_is_fencei : _slots_10_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_48 ? _slots_13_io_out_uop_is_amo : _GEN_47 ? _slots_12_io_out_uop_is_amo : _GEN_46 ? _slots_11_io_out_uop_is_amo : _slots_10_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_48 ? _slots_13_io_out_uop_uses_ldq : _GEN_47 ? _slots_12_io_out_uop_uses_ldq : _GEN_46 ? _slots_11_io_out_uop_uses_ldq : _slots_10_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_48 ? _slots_13_io_out_uop_uses_stq : _GEN_47 ? _slots_12_io_out_uop_uses_stq : _GEN_46 ? _slots_11_io_out_uop_uses_stq : _slots_10_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_48 ? _slots_13_io_out_uop_is_sys_pc2epc : _GEN_47 ? _slots_12_io_out_uop_is_sys_pc2epc : _GEN_46 ? _slots_11_io_out_uop_is_sys_pc2epc : _slots_10_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_48 ? _slots_13_io_out_uop_is_unique : _GEN_47 ? _slots_12_io_out_uop_is_unique : _GEN_46 ? _slots_11_io_out_uop_is_unique : _slots_10_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_48 ? _slots_13_io_out_uop_flush_on_commit : _GEN_47 ? _slots_12_io_out_uop_flush_on_commit : _GEN_46 ? _slots_11_io_out_uop_flush_on_commit : _slots_10_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_48 ? _slots_13_io_out_uop_ldst_is_rs1 : _GEN_47 ? _slots_12_io_out_uop_ldst_is_rs1 : _GEN_46 ? _slots_11_io_out_uop_ldst_is_rs1 : _slots_10_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_48 ? _slots_13_io_out_uop_ldst : _GEN_47 ? _slots_12_io_out_uop_ldst : _GEN_46 ? _slots_11_io_out_uop_ldst : _slots_10_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_48 ? _slots_13_io_out_uop_lrs1 : _GEN_47 ? _slots_12_io_out_uop_lrs1 : _GEN_46 ? _slots_11_io_out_uop_lrs1 : _slots_10_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_48 ? _slots_13_io_out_uop_lrs2 : _GEN_47 ? _slots_12_io_out_uop_lrs2 : _GEN_46 ? _slots_11_io_out_uop_lrs2 : _slots_10_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_48 ? _slots_13_io_out_uop_lrs3 : _GEN_47 ? _slots_12_io_out_uop_lrs3 : _GEN_46 ? _slots_11_io_out_uop_lrs3 : _slots_10_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_48 ? _slots_13_io_out_uop_ldst_val : _GEN_47 ? _slots_12_io_out_uop_ldst_val : _GEN_46 ? _slots_11_io_out_uop_ldst_val : _slots_10_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_48 ? _slots_13_io_out_uop_dst_rtype : _GEN_47 ? _slots_12_io_out_uop_dst_rtype : _GEN_46 ? _slots_11_io_out_uop_dst_rtype : _slots_10_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_48 ? _slots_13_io_out_uop_lrs1_rtype : _GEN_47 ? _slots_12_io_out_uop_lrs1_rtype : _GEN_46 ? _slots_11_io_out_uop_lrs1_rtype : _slots_10_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_48 ? _slots_13_io_out_uop_lrs2_rtype : _GEN_47 ? _slots_12_io_out_uop_lrs2_rtype : _GEN_46 ? _slots_11_io_out_uop_lrs2_rtype : _slots_10_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_48 ? _slots_13_io_out_uop_frs3_en : _GEN_47 ? _slots_12_io_out_uop_frs3_en : _GEN_46 ? _slots_11_io_out_uop_frs3_en : _slots_10_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_48 ? _slots_13_io_out_uop_fp_val : _GEN_47 ? _slots_12_io_out_uop_fp_val : _GEN_46 ? _slots_11_io_out_uop_fp_val : _slots_10_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_48 ? _slots_13_io_out_uop_fp_single : _GEN_47 ? _slots_12_io_out_uop_fp_single : _GEN_46 ? _slots_11_io_out_uop_fp_single : _slots_10_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_48 ? _slots_13_io_out_uop_xcpt_pf_if : _GEN_47 ? _slots_12_io_out_uop_xcpt_pf_if : _GEN_46 ? _slots_11_io_out_uop_xcpt_pf_if : _slots_10_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_48 ? _slots_13_io_out_uop_xcpt_ae_if : _GEN_47 ? _slots_12_io_out_uop_xcpt_ae_if : _GEN_46 ? _slots_11_io_out_uop_xcpt_ae_if : _slots_10_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_48 ? _slots_13_io_out_uop_xcpt_ma_if : _GEN_47 ? _slots_12_io_out_uop_xcpt_ma_if : _GEN_46 ? _slots_11_io_out_uop_xcpt_ma_if : _slots_10_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_48 ? _slots_13_io_out_uop_bp_debug_if : _GEN_47 ? _slots_12_io_out_uop_bp_debug_if : _GEN_46 ? _slots_11_io_out_uop_bp_debug_if : _slots_10_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_48 ? _slots_13_io_out_uop_bp_xcpt_if : _GEN_47 ? _slots_12_io_out_uop_bp_xcpt_if : _GEN_46 ? _slots_11_io_out_uop_bp_xcpt_if : _slots_10_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_48 ? _slots_13_io_out_uop_debug_fsrc : _GEN_47 ? _slots_12_io_out_uop_debug_fsrc : _GEN_46 ? _slots_11_io_out_uop_debug_fsrc : _slots_10_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_48 ? _slots_13_io_out_uop_debug_tsrc : _GEN_47 ? _slots_12_io_out_uop_debug_tsrc : _GEN_46 ? _slots_11_io_out_uop_debug_tsrc : _slots_10_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_9_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_9_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_9_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_9_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_9_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_9_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_9_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_9_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_9_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_9_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_9_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_9_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_9_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_9_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_9_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_9_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_9_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_9_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_9_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_9_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_9_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_9_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_9_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_9_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_9_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_9_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_9_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_9_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_9_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_9_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_9_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_9_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_9_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_9_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_9_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_9_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_9_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_9_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_9_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_9_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_9_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_9_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_9_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_9_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_9_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_9_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_9_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_9_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_9_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_9_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_9_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_9_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_9_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_9_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_9_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_9_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_9_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_9_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_9_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_9_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_9_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_9_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_9_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_9_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_9_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_9_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_9_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_9_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_9_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_9_io_uop_uopc),
    .io_uop_inst                    (_slots_9_io_uop_inst),
    .io_uop_debug_inst              (_slots_9_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_9_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_9_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_9_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_9_io_uop_fu_code),
    .io_uop_iw_state                (_slots_9_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_9_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_9_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_9_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_9_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_9_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_9_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_9_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_9_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_9_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_9_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_9_io_uop_pc_lob),
    .io_uop_taken                   (_slots_9_io_uop_taken),
    .io_uop_imm_packed              (_slots_9_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_9_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_9_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_9_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_9_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_9_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_9_io_uop_pdst),
    .io_uop_prs1                    (_slots_9_io_uop_prs1),
    .io_uop_prs2                    (_slots_9_io_uop_prs2),
    .io_uop_prs3                    (_slots_9_io_uop_prs3),
    .io_uop_ppred                   (_slots_9_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_9_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_9_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_9_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_9_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_9_io_uop_stale_pdst),
    .io_uop_exception               (_slots_9_io_uop_exception),
    .io_uop_exc_cause               (_slots_9_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_9_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_9_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_9_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_9_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_9_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_9_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_9_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_9_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_9_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_9_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_9_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_9_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_9_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_9_io_uop_ldst),
    .io_uop_lrs1                    (_slots_9_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_9_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_9_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_9_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_9_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_9_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_9_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_9_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_9_io_uop_fp_val),
    .io_uop_fp_single               (_slots_9_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_9_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_9_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_9_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_9_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_9_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_9_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_9_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_10 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_10_io_valid),
    .io_will_be_valid               (_slots_10_io_will_be_valid),
    .io_request                     (_slots_10_io_request),
    .io_grant                       (issue_slots_10_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_9),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_10_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_51 ? _slots_14_io_out_uop_uopc : _GEN_50 ? _slots_13_io_out_uop_uopc : _GEN_49 ? _slots_12_io_out_uop_uopc : _slots_11_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_51 ? _slots_14_io_out_uop_inst : _GEN_50 ? _slots_13_io_out_uop_inst : _GEN_49 ? _slots_12_io_out_uop_inst : _slots_11_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_51 ? _slots_14_io_out_uop_debug_inst : _GEN_50 ? _slots_13_io_out_uop_debug_inst : _GEN_49 ? _slots_12_io_out_uop_debug_inst : _slots_11_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_51 ? _slots_14_io_out_uop_is_rvc : _GEN_50 ? _slots_13_io_out_uop_is_rvc : _GEN_49 ? _slots_12_io_out_uop_is_rvc : _slots_11_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_51 ? _slots_14_io_out_uop_debug_pc : _GEN_50 ? _slots_13_io_out_uop_debug_pc : _GEN_49 ? _slots_12_io_out_uop_debug_pc : _slots_11_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_51 ? _slots_14_io_out_uop_iq_type : _GEN_50 ? _slots_13_io_out_uop_iq_type : _GEN_49 ? _slots_12_io_out_uop_iq_type : _slots_11_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_51 ? _slots_14_io_out_uop_fu_code : _GEN_50 ? _slots_13_io_out_uop_fu_code : _GEN_49 ? _slots_12_io_out_uop_fu_code : _slots_11_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_51 ? _slots_14_io_out_uop_iw_state : _GEN_50 ? _slots_13_io_out_uop_iw_state : _GEN_49 ? _slots_12_io_out_uop_iw_state : _slots_11_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_51 ? _slots_14_io_out_uop_iw_p1_poisoned : _GEN_50 ? _slots_13_io_out_uop_iw_p1_poisoned : _GEN_49 ? _slots_12_io_out_uop_iw_p1_poisoned : _slots_11_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_51 ? _slots_14_io_out_uop_iw_p2_poisoned : _GEN_50 ? _slots_13_io_out_uop_iw_p2_poisoned : _GEN_49 ? _slots_12_io_out_uop_iw_p2_poisoned : _slots_11_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_51 ? _slots_14_io_out_uop_is_br : _GEN_50 ? _slots_13_io_out_uop_is_br : _GEN_49 ? _slots_12_io_out_uop_is_br : _slots_11_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_51 ? _slots_14_io_out_uop_is_jalr : _GEN_50 ? _slots_13_io_out_uop_is_jalr : _GEN_49 ? _slots_12_io_out_uop_is_jalr : _slots_11_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_51 ? _slots_14_io_out_uop_is_jal : _GEN_50 ? _slots_13_io_out_uop_is_jal : _GEN_49 ? _slots_12_io_out_uop_is_jal : _slots_11_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_51 ? _slots_14_io_out_uop_is_sfb : _GEN_50 ? _slots_13_io_out_uop_is_sfb : _GEN_49 ? _slots_12_io_out_uop_is_sfb : _slots_11_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_51 ? _slots_14_io_out_uop_br_mask : _GEN_50 ? _slots_13_io_out_uop_br_mask : _GEN_49 ? _slots_12_io_out_uop_br_mask : _slots_11_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_51 ? _slots_14_io_out_uop_br_tag : _GEN_50 ? _slots_13_io_out_uop_br_tag : _GEN_49 ? _slots_12_io_out_uop_br_tag : _slots_11_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_51 ? _slots_14_io_out_uop_ftq_idx : _GEN_50 ? _slots_13_io_out_uop_ftq_idx : _GEN_49 ? _slots_12_io_out_uop_ftq_idx : _slots_11_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_51 ? _slots_14_io_out_uop_edge_inst : _GEN_50 ? _slots_13_io_out_uop_edge_inst : _GEN_49 ? _slots_12_io_out_uop_edge_inst : _slots_11_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_51 ? _slots_14_io_out_uop_pc_lob : _GEN_50 ? _slots_13_io_out_uop_pc_lob : _GEN_49 ? _slots_12_io_out_uop_pc_lob : _slots_11_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_51 ? _slots_14_io_out_uop_taken : _GEN_50 ? _slots_13_io_out_uop_taken : _GEN_49 ? _slots_12_io_out_uop_taken : _slots_11_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_51 ? _slots_14_io_out_uop_imm_packed : _GEN_50 ? _slots_13_io_out_uop_imm_packed : _GEN_49 ? _slots_12_io_out_uop_imm_packed : _slots_11_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_51 ? _slots_14_io_out_uop_csr_addr : _GEN_50 ? _slots_13_io_out_uop_csr_addr : _GEN_49 ? _slots_12_io_out_uop_csr_addr : _slots_11_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_51 ? _slots_14_io_out_uop_rob_idx : _GEN_50 ? _slots_13_io_out_uop_rob_idx : _GEN_49 ? _slots_12_io_out_uop_rob_idx : _slots_11_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_51 ? _slots_14_io_out_uop_ldq_idx : _GEN_50 ? _slots_13_io_out_uop_ldq_idx : _GEN_49 ? _slots_12_io_out_uop_ldq_idx : _slots_11_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_51 ? _slots_14_io_out_uop_stq_idx : _GEN_50 ? _slots_13_io_out_uop_stq_idx : _GEN_49 ? _slots_12_io_out_uop_stq_idx : _slots_11_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_51 ? _slots_14_io_out_uop_rxq_idx : _GEN_50 ? _slots_13_io_out_uop_rxq_idx : _GEN_49 ? _slots_12_io_out_uop_rxq_idx : _slots_11_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_51 ? _slots_14_io_out_uop_pdst : _GEN_50 ? _slots_13_io_out_uop_pdst : _GEN_49 ? _slots_12_io_out_uop_pdst : _slots_11_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_51 ? _slots_14_io_out_uop_prs1 : _GEN_50 ? _slots_13_io_out_uop_prs1 : _GEN_49 ? _slots_12_io_out_uop_prs1 : _slots_11_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_51 ? _slots_14_io_out_uop_prs2 : _GEN_50 ? _slots_13_io_out_uop_prs2 : _GEN_49 ? _slots_12_io_out_uop_prs2 : _slots_11_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_51 ? _slots_14_io_out_uop_prs3 : _GEN_50 ? _slots_13_io_out_uop_prs3 : _GEN_49 ? _slots_12_io_out_uop_prs3 : _slots_11_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_51 ? _slots_14_io_out_uop_ppred : _GEN_50 ? _slots_13_io_out_uop_ppred : _GEN_49 ? _slots_12_io_out_uop_ppred : _slots_11_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_51 ? _slots_14_io_out_uop_prs1_busy : _GEN_50 ? _slots_13_io_out_uop_prs1_busy : _GEN_49 ? _slots_12_io_out_uop_prs1_busy : _slots_11_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_51 ? _slots_14_io_out_uop_prs2_busy : _GEN_50 ? _slots_13_io_out_uop_prs2_busy : _GEN_49 ? _slots_12_io_out_uop_prs2_busy : _slots_11_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_51 ? _slots_14_io_out_uop_prs3_busy : _GEN_50 ? _slots_13_io_out_uop_prs3_busy : _GEN_49 ? _slots_12_io_out_uop_prs3_busy : _slots_11_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_51 ? _slots_14_io_out_uop_ppred_busy : _GEN_50 ? _slots_13_io_out_uop_ppred_busy : _GEN_49 ? _slots_12_io_out_uop_ppred_busy : _slots_11_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_51 ? _slots_14_io_out_uop_stale_pdst : _GEN_50 ? _slots_13_io_out_uop_stale_pdst : _GEN_49 ? _slots_12_io_out_uop_stale_pdst : _slots_11_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_51 ? _slots_14_io_out_uop_exception : _GEN_50 ? _slots_13_io_out_uop_exception : _GEN_49 ? _slots_12_io_out_uop_exception : _slots_11_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_51 ? _slots_14_io_out_uop_exc_cause : _GEN_50 ? _slots_13_io_out_uop_exc_cause : _GEN_49 ? _slots_12_io_out_uop_exc_cause : _slots_11_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_51 ? _slots_14_io_out_uop_bypassable : _GEN_50 ? _slots_13_io_out_uop_bypassable : _GEN_49 ? _slots_12_io_out_uop_bypassable : _slots_11_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_51 ? _slots_14_io_out_uop_mem_cmd : _GEN_50 ? _slots_13_io_out_uop_mem_cmd : _GEN_49 ? _slots_12_io_out_uop_mem_cmd : _slots_11_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_51 ? _slots_14_io_out_uop_mem_size : _GEN_50 ? _slots_13_io_out_uop_mem_size : _GEN_49 ? _slots_12_io_out_uop_mem_size : _slots_11_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_51 ? _slots_14_io_out_uop_mem_signed : _GEN_50 ? _slots_13_io_out_uop_mem_signed : _GEN_49 ? _slots_12_io_out_uop_mem_signed : _slots_11_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_51 ? _slots_14_io_out_uop_is_fence : _GEN_50 ? _slots_13_io_out_uop_is_fence : _GEN_49 ? _slots_12_io_out_uop_is_fence : _slots_11_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_51 ? _slots_14_io_out_uop_is_fencei : _GEN_50 ? _slots_13_io_out_uop_is_fencei : _GEN_49 ? _slots_12_io_out_uop_is_fencei : _slots_11_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_51 ? _slots_14_io_out_uop_is_amo : _GEN_50 ? _slots_13_io_out_uop_is_amo : _GEN_49 ? _slots_12_io_out_uop_is_amo : _slots_11_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_51 ? _slots_14_io_out_uop_uses_ldq : _GEN_50 ? _slots_13_io_out_uop_uses_ldq : _GEN_49 ? _slots_12_io_out_uop_uses_ldq : _slots_11_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_51 ? _slots_14_io_out_uop_uses_stq : _GEN_50 ? _slots_13_io_out_uop_uses_stq : _GEN_49 ? _slots_12_io_out_uop_uses_stq : _slots_11_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_51 ? _slots_14_io_out_uop_is_sys_pc2epc : _GEN_50 ? _slots_13_io_out_uop_is_sys_pc2epc : _GEN_49 ? _slots_12_io_out_uop_is_sys_pc2epc : _slots_11_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_51 ? _slots_14_io_out_uop_is_unique : _GEN_50 ? _slots_13_io_out_uop_is_unique : _GEN_49 ? _slots_12_io_out_uop_is_unique : _slots_11_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_51 ? _slots_14_io_out_uop_flush_on_commit : _GEN_50 ? _slots_13_io_out_uop_flush_on_commit : _GEN_49 ? _slots_12_io_out_uop_flush_on_commit : _slots_11_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_51 ? _slots_14_io_out_uop_ldst_is_rs1 : _GEN_50 ? _slots_13_io_out_uop_ldst_is_rs1 : _GEN_49 ? _slots_12_io_out_uop_ldst_is_rs1 : _slots_11_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_51 ? _slots_14_io_out_uop_ldst : _GEN_50 ? _slots_13_io_out_uop_ldst : _GEN_49 ? _slots_12_io_out_uop_ldst : _slots_11_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_51 ? _slots_14_io_out_uop_lrs1 : _GEN_50 ? _slots_13_io_out_uop_lrs1 : _GEN_49 ? _slots_12_io_out_uop_lrs1 : _slots_11_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_51 ? _slots_14_io_out_uop_lrs2 : _GEN_50 ? _slots_13_io_out_uop_lrs2 : _GEN_49 ? _slots_12_io_out_uop_lrs2 : _slots_11_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_51 ? _slots_14_io_out_uop_lrs3 : _GEN_50 ? _slots_13_io_out_uop_lrs3 : _GEN_49 ? _slots_12_io_out_uop_lrs3 : _slots_11_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_51 ? _slots_14_io_out_uop_ldst_val : _GEN_50 ? _slots_13_io_out_uop_ldst_val : _GEN_49 ? _slots_12_io_out_uop_ldst_val : _slots_11_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_51 ? _slots_14_io_out_uop_dst_rtype : _GEN_50 ? _slots_13_io_out_uop_dst_rtype : _GEN_49 ? _slots_12_io_out_uop_dst_rtype : _slots_11_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_51 ? _slots_14_io_out_uop_lrs1_rtype : _GEN_50 ? _slots_13_io_out_uop_lrs1_rtype : _GEN_49 ? _slots_12_io_out_uop_lrs1_rtype : _slots_11_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_51 ? _slots_14_io_out_uop_lrs2_rtype : _GEN_50 ? _slots_13_io_out_uop_lrs2_rtype : _GEN_49 ? _slots_12_io_out_uop_lrs2_rtype : _slots_11_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_51 ? _slots_14_io_out_uop_frs3_en : _GEN_50 ? _slots_13_io_out_uop_frs3_en : _GEN_49 ? _slots_12_io_out_uop_frs3_en : _slots_11_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_51 ? _slots_14_io_out_uop_fp_val : _GEN_50 ? _slots_13_io_out_uop_fp_val : _GEN_49 ? _slots_12_io_out_uop_fp_val : _slots_11_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_51 ? _slots_14_io_out_uop_fp_single : _GEN_50 ? _slots_13_io_out_uop_fp_single : _GEN_49 ? _slots_12_io_out_uop_fp_single : _slots_11_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_51 ? _slots_14_io_out_uop_xcpt_pf_if : _GEN_50 ? _slots_13_io_out_uop_xcpt_pf_if : _GEN_49 ? _slots_12_io_out_uop_xcpt_pf_if : _slots_11_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_51 ? _slots_14_io_out_uop_xcpt_ae_if : _GEN_50 ? _slots_13_io_out_uop_xcpt_ae_if : _GEN_49 ? _slots_12_io_out_uop_xcpt_ae_if : _slots_11_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_51 ? _slots_14_io_out_uop_xcpt_ma_if : _GEN_50 ? _slots_13_io_out_uop_xcpt_ma_if : _GEN_49 ? _slots_12_io_out_uop_xcpt_ma_if : _slots_11_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_51 ? _slots_14_io_out_uop_bp_debug_if : _GEN_50 ? _slots_13_io_out_uop_bp_debug_if : _GEN_49 ? _slots_12_io_out_uop_bp_debug_if : _slots_11_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_51 ? _slots_14_io_out_uop_bp_xcpt_if : _GEN_50 ? _slots_13_io_out_uop_bp_xcpt_if : _GEN_49 ? _slots_12_io_out_uop_bp_xcpt_if : _slots_11_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_51 ? _slots_14_io_out_uop_debug_fsrc : _GEN_50 ? _slots_13_io_out_uop_debug_fsrc : _GEN_49 ? _slots_12_io_out_uop_debug_fsrc : _slots_11_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_51 ? _slots_14_io_out_uop_debug_tsrc : _GEN_50 ? _slots_13_io_out_uop_debug_tsrc : _GEN_49 ? _slots_12_io_out_uop_debug_tsrc : _slots_11_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_10_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_10_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_10_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_10_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_10_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_10_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_10_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_10_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_10_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_10_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_10_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_10_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_10_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_10_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_10_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_10_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_10_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_10_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_10_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_10_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_10_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_10_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_10_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_10_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_10_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_10_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_10_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_10_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_10_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_10_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_10_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_10_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_10_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_10_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_10_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_10_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_10_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_10_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_10_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_10_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_10_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_10_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_10_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_10_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_10_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_10_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_10_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_10_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_10_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_10_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_10_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_10_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_10_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_10_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_10_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_10_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_10_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_10_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_10_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_10_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_10_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_10_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_10_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_10_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_10_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_10_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_10_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_10_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_10_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_10_io_uop_uopc),
    .io_uop_inst                    (_slots_10_io_uop_inst),
    .io_uop_debug_inst              (_slots_10_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_10_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_10_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_10_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_10_io_uop_fu_code),
    .io_uop_iw_state                (_slots_10_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_10_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_10_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_10_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_10_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_10_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_10_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_10_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_10_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_10_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_10_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_10_io_uop_pc_lob),
    .io_uop_taken                   (_slots_10_io_uop_taken),
    .io_uop_imm_packed              (_slots_10_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_10_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_10_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_10_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_10_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_10_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_10_io_uop_pdst),
    .io_uop_prs1                    (_slots_10_io_uop_prs1),
    .io_uop_prs2                    (_slots_10_io_uop_prs2),
    .io_uop_prs3                    (_slots_10_io_uop_prs3),
    .io_uop_ppred                   (_slots_10_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_10_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_10_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_10_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_10_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_10_io_uop_stale_pdst),
    .io_uop_exception               (_slots_10_io_uop_exception),
    .io_uop_exc_cause               (_slots_10_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_10_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_10_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_10_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_10_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_10_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_10_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_10_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_10_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_10_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_10_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_10_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_10_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_10_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_10_io_uop_ldst),
    .io_uop_lrs1                    (_slots_10_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_10_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_10_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_10_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_10_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_10_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_10_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_10_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_10_io_uop_fp_val),
    .io_uop_fp_single               (_slots_10_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_10_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_10_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_10_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_10_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_10_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_10_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_10_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_11 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_11_io_valid),
    .io_will_be_valid               (_slots_11_io_will_be_valid),
    .io_request                     (_slots_11_io_request),
    .io_grant                       (issue_slots_11_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_10),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_11_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_54 ? _slots_15_io_out_uop_uopc : _GEN_53 ? _slots_14_io_out_uop_uopc : _GEN_52 ? _slots_13_io_out_uop_uopc : _slots_12_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_54 ? _slots_15_io_out_uop_inst : _GEN_53 ? _slots_14_io_out_uop_inst : _GEN_52 ? _slots_13_io_out_uop_inst : _slots_12_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_54 ? _slots_15_io_out_uop_debug_inst : _GEN_53 ? _slots_14_io_out_uop_debug_inst : _GEN_52 ? _slots_13_io_out_uop_debug_inst : _slots_12_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_54 ? _slots_15_io_out_uop_is_rvc : _GEN_53 ? _slots_14_io_out_uop_is_rvc : _GEN_52 ? _slots_13_io_out_uop_is_rvc : _slots_12_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_54 ? _slots_15_io_out_uop_debug_pc : _GEN_53 ? _slots_14_io_out_uop_debug_pc : _GEN_52 ? _slots_13_io_out_uop_debug_pc : _slots_12_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_54 ? _slots_15_io_out_uop_iq_type : _GEN_53 ? _slots_14_io_out_uop_iq_type : _GEN_52 ? _slots_13_io_out_uop_iq_type : _slots_12_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_54 ? _slots_15_io_out_uop_fu_code : _GEN_53 ? _slots_14_io_out_uop_fu_code : _GEN_52 ? _slots_13_io_out_uop_fu_code : _slots_12_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_54 ? _slots_15_io_out_uop_iw_state : _GEN_53 ? _slots_14_io_out_uop_iw_state : _GEN_52 ? _slots_13_io_out_uop_iw_state : _slots_12_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_54 ? _slots_15_io_out_uop_iw_p1_poisoned : _GEN_53 ? _slots_14_io_out_uop_iw_p1_poisoned : _GEN_52 ? _slots_13_io_out_uop_iw_p1_poisoned : _slots_12_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_54 ? _slots_15_io_out_uop_iw_p2_poisoned : _GEN_53 ? _slots_14_io_out_uop_iw_p2_poisoned : _GEN_52 ? _slots_13_io_out_uop_iw_p2_poisoned : _slots_12_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_54 ? _slots_15_io_out_uop_is_br : _GEN_53 ? _slots_14_io_out_uop_is_br : _GEN_52 ? _slots_13_io_out_uop_is_br : _slots_12_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_54 ? _slots_15_io_out_uop_is_jalr : _GEN_53 ? _slots_14_io_out_uop_is_jalr : _GEN_52 ? _slots_13_io_out_uop_is_jalr : _slots_12_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_54 ? _slots_15_io_out_uop_is_jal : _GEN_53 ? _slots_14_io_out_uop_is_jal : _GEN_52 ? _slots_13_io_out_uop_is_jal : _slots_12_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_54 ? _slots_15_io_out_uop_is_sfb : _GEN_53 ? _slots_14_io_out_uop_is_sfb : _GEN_52 ? _slots_13_io_out_uop_is_sfb : _slots_12_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_54 ? _slots_15_io_out_uop_br_mask : _GEN_53 ? _slots_14_io_out_uop_br_mask : _GEN_52 ? _slots_13_io_out_uop_br_mask : _slots_12_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_54 ? _slots_15_io_out_uop_br_tag : _GEN_53 ? _slots_14_io_out_uop_br_tag : _GEN_52 ? _slots_13_io_out_uop_br_tag : _slots_12_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_54 ? _slots_15_io_out_uop_ftq_idx : _GEN_53 ? _slots_14_io_out_uop_ftq_idx : _GEN_52 ? _slots_13_io_out_uop_ftq_idx : _slots_12_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_54 ? _slots_15_io_out_uop_edge_inst : _GEN_53 ? _slots_14_io_out_uop_edge_inst : _GEN_52 ? _slots_13_io_out_uop_edge_inst : _slots_12_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_54 ? _slots_15_io_out_uop_pc_lob : _GEN_53 ? _slots_14_io_out_uop_pc_lob : _GEN_52 ? _slots_13_io_out_uop_pc_lob : _slots_12_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_54 ? _slots_15_io_out_uop_taken : _GEN_53 ? _slots_14_io_out_uop_taken : _GEN_52 ? _slots_13_io_out_uop_taken : _slots_12_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_54 ? _slots_15_io_out_uop_imm_packed : _GEN_53 ? _slots_14_io_out_uop_imm_packed : _GEN_52 ? _slots_13_io_out_uop_imm_packed : _slots_12_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_54 ? _slots_15_io_out_uop_csr_addr : _GEN_53 ? _slots_14_io_out_uop_csr_addr : _GEN_52 ? _slots_13_io_out_uop_csr_addr : _slots_12_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_54 ? _slots_15_io_out_uop_rob_idx : _GEN_53 ? _slots_14_io_out_uop_rob_idx : _GEN_52 ? _slots_13_io_out_uop_rob_idx : _slots_12_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_54 ? _slots_15_io_out_uop_ldq_idx : _GEN_53 ? _slots_14_io_out_uop_ldq_idx : _GEN_52 ? _slots_13_io_out_uop_ldq_idx : _slots_12_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_54 ? _slots_15_io_out_uop_stq_idx : _GEN_53 ? _slots_14_io_out_uop_stq_idx : _GEN_52 ? _slots_13_io_out_uop_stq_idx : _slots_12_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_54 ? _slots_15_io_out_uop_rxq_idx : _GEN_53 ? _slots_14_io_out_uop_rxq_idx : _GEN_52 ? _slots_13_io_out_uop_rxq_idx : _slots_12_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_54 ? _slots_15_io_out_uop_pdst : _GEN_53 ? _slots_14_io_out_uop_pdst : _GEN_52 ? _slots_13_io_out_uop_pdst : _slots_12_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_54 ? _slots_15_io_out_uop_prs1 : _GEN_53 ? _slots_14_io_out_uop_prs1 : _GEN_52 ? _slots_13_io_out_uop_prs1 : _slots_12_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_54 ? _slots_15_io_out_uop_prs2 : _GEN_53 ? _slots_14_io_out_uop_prs2 : _GEN_52 ? _slots_13_io_out_uop_prs2 : _slots_12_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_54 ? _slots_15_io_out_uop_prs3 : _GEN_53 ? _slots_14_io_out_uop_prs3 : _GEN_52 ? _slots_13_io_out_uop_prs3 : _slots_12_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_54 ? _slots_15_io_out_uop_ppred : _GEN_53 ? _slots_14_io_out_uop_ppred : _GEN_52 ? _slots_13_io_out_uop_ppred : _slots_12_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_54 ? _slots_15_io_out_uop_prs1_busy : _GEN_53 ? _slots_14_io_out_uop_prs1_busy : _GEN_52 ? _slots_13_io_out_uop_prs1_busy : _slots_12_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_54 ? _slots_15_io_out_uop_prs2_busy : _GEN_53 ? _slots_14_io_out_uop_prs2_busy : _GEN_52 ? _slots_13_io_out_uop_prs2_busy : _slots_12_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_54 ? _slots_15_io_out_uop_prs3_busy : _GEN_53 ? _slots_14_io_out_uop_prs3_busy : _GEN_52 ? _slots_13_io_out_uop_prs3_busy : _slots_12_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_54 ? _slots_15_io_out_uop_ppred_busy : _GEN_53 ? _slots_14_io_out_uop_ppred_busy : _GEN_52 ? _slots_13_io_out_uop_ppred_busy : _slots_12_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_54 ? _slots_15_io_out_uop_stale_pdst : _GEN_53 ? _slots_14_io_out_uop_stale_pdst : _GEN_52 ? _slots_13_io_out_uop_stale_pdst : _slots_12_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_54 ? _slots_15_io_out_uop_exception : _GEN_53 ? _slots_14_io_out_uop_exception : _GEN_52 ? _slots_13_io_out_uop_exception : _slots_12_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_54 ? _slots_15_io_out_uop_exc_cause : _GEN_53 ? _slots_14_io_out_uop_exc_cause : _GEN_52 ? _slots_13_io_out_uop_exc_cause : _slots_12_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_54 ? _slots_15_io_out_uop_bypassable : _GEN_53 ? _slots_14_io_out_uop_bypassable : _GEN_52 ? _slots_13_io_out_uop_bypassable : _slots_12_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_54 ? _slots_15_io_out_uop_mem_cmd : _GEN_53 ? _slots_14_io_out_uop_mem_cmd : _GEN_52 ? _slots_13_io_out_uop_mem_cmd : _slots_12_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_54 ? _slots_15_io_out_uop_mem_size : _GEN_53 ? _slots_14_io_out_uop_mem_size : _GEN_52 ? _slots_13_io_out_uop_mem_size : _slots_12_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_54 ? _slots_15_io_out_uop_mem_signed : _GEN_53 ? _slots_14_io_out_uop_mem_signed : _GEN_52 ? _slots_13_io_out_uop_mem_signed : _slots_12_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_54 ? _slots_15_io_out_uop_is_fence : _GEN_53 ? _slots_14_io_out_uop_is_fence : _GEN_52 ? _slots_13_io_out_uop_is_fence : _slots_12_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_54 ? _slots_15_io_out_uop_is_fencei : _GEN_53 ? _slots_14_io_out_uop_is_fencei : _GEN_52 ? _slots_13_io_out_uop_is_fencei : _slots_12_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_54 ? _slots_15_io_out_uop_is_amo : _GEN_53 ? _slots_14_io_out_uop_is_amo : _GEN_52 ? _slots_13_io_out_uop_is_amo : _slots_12_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_54 ? _slots_15_io_out_uop_uses_ldq : _GEN_53 ? _slots_14_io_out_uop_uses_ldq : _GEN_52 ? _slots_13_io_out_uop_uses_ldq : _slots_12_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_54 ? _slots_15_io_out_uop_uses_stq : _GEN_53 ? _slots_14_io_out_uop_uses_stq : _GEN_52 ? _slots_13_io_out_uop_uses_stq : _slots_12_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_54 ? _slots_15_io_out_uop_is_sys_pc2epc : _GEN_53 ? _slots_14_io_out_uop_is_sys_pc2epc : _GEN_52 ? _slots_13_io_out_uop_is_sys_pc2epc : _slots_12_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_54 ? _slots_15_io_out_uop_is_unique : _GEN_53 ? _slots_14_io_out_uop_is_unique : _GEN_52 ? _slots_13_io_out_uop_is_unique : _slots_12_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_54 ? _slots_15_io_out_uop_flush_on_commit : _GEN_53 ? _slots_14_io_out_uop_flush_on_commit : _GEN_52 ? _slots_13_io_out_uop_flush_on_commit : _slots_12_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_54 ? _slots_15_io_out_uop_ldst_is_rs1 : _GEN_53 ? _slots_14_io_out_uop_ldst_is_rs1 : _GEN_52 ? _slots_13_io_out_uop_ldst_is_rs1 : _slots_12_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_54 ? _slots_15_io_out_uop_ldst : _GEN_53 ? _slots_14_io_out_uop_ldst : _GEN_52 ? _slots_13_io_out_uop_ldst : _slots_12_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_54 ? _slots_15_io_out_uop_lrs1 : _GEN_53 ? _slots_14_io_out_uop_lrs1 : _GEN_52 ? _slots_13_io_out_uop_lrs1 : _slots_12_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_54 ? _slots_15_io_out_uop_lrs2 : _GEN_53 ? _slots_14_io_out_uop_lrs2 : _GEN_52 ? _slots_13_io_out_uop_lrs2 : _slots_12_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_54 ? _slots_15_io_out_uop_lrs3 : _GEN_53 ? _slots_14_io_out_uop_lrs3 : _GEN_52 ? _slots_13_io_out_uop_lrs3 : _slots_12_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_54 ? _slots_15_io_out_uop_ldst_val : _GEN_53 ? _slots_14_io_out_uop_ldst_val : _GEN_52 ? _slots_13_io_out_uop_ldst_val : _slots_12_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_54 ? _slots_15_io_out_uop_dst_rtype : _GEN_53 ? _slots_14_io_out_uop_dst_rtype : _GEN_52 ? _slots_13_io_out_uop_dst_rtype : _slots_12_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_54 ? _slots_15_io_out_uop_lrs1_rtype : _GEN_53 ? _slots_14_io_out_uop_lrs1_rtype : _GEN_52 ? _slots_13_io_out_uop_lrs1_rtype : _slots_12_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_54 ? _slots_15_io_out_uop_lrs2_rtype : _GEN_53 ? _slots_14_io_out_uop_lrs2_rtype : _GEN_52 ? _slots_13_io_out_uop_lrs2_rtype : _slots_12_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_54 ? _slots_15_io_out_uop_frs3_en : _GEN_53 ? _slots_14_io_out_uop_frs3_en : _GEN_52 ? _slots_13_io_out_uop_frs3_en : _slots_12_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_54 ? _slots_15_io_out_uop_fp_val : _GEN_53 ? _slots_14_io_out_uop_fp_val : _GEN_52 ? _slots_13_io_out_uop_fp_val : _slots_12_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_54 ? _slots_15_io_out_uop_fp_single : _GEN_53 ? _slots_14_io_out_uop_fp_single : _GEN_52 ? _slots_13_io_out_uop_fp_single : _slots_12_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_54 ? _slots_15_io_out_uop_xcpt_pf_if : _GEN_53 ? _slots_14_io_out_uop_xcpt_pf_if : _GEN_52 ? _slots_13_io_out_uop_xcpt_pf_if : _slots_12_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_54 ? _slots_15_io_out_uop_xcpt_ae_if : _GEN_53 ? _slots_14_io_out_uop_xcpt_ae_if : _GEN_52 ? _slots_13_io_out_uop_xcpt_ae_if : _slots_12_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_54 ? _slots_15_io_out_uop_xcpt_ma_if : _GEN_53 ? _slots_14_io_out_uop_xcpt_ma_if : _GEN_52 ? _slots_13_io_out_uop_xcpt_ma_if : _slots_12_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_54 ? _slots_15_io_out_uop_bp_debug_if : _GEN_53 ? _slots_14_io_out_uop_bp_debug_if : _GEN_52 ? _slots_13_io_out_uop_bp_debug_if : _slots_12_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_54 ? _slots_15_io_out_uop_bp_xcpt_if : _GEN_53 ? _slots_14_io_out_uop_bp_xcpt_if : _GEN_52 ? _slots_13_io_out_uop_bp_xcpt_if : _slots_12_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_54 ? _slots_15_io_out_uop_debug_fsrc : _GEN_53 ? _slots_14_io_out_uop_debug_fsrc : _GEN_52 ? _slots_13_io_out_uop_debug_fsrc : _slots_12_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_54 ? _slots_15_io_out_uop_debug_tsrc : _GEN_53 ? _slots_14_io_out_uop_debug_tsrc : _GEN_52 ? _slots_13_io_out_uop_debug_tsrc : _slots_12_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_11_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_11_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_11_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_11_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_11_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_11_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_11_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_11_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_11_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_11_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_11_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_11_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_11_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_11_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_11_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_11_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_11_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_11_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_11_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_11_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_11_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_11_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_11_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_11_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_11_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_11_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_11_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_11_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_11_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_11_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_11_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_11_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_11_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_11_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_11_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_11_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_11_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_11_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_11_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_11_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_11_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_11_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_11_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_11_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_11_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_11_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_11_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_11_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_11_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_11_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_11_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_11_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_11_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_11_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_11_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_11_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_11_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_11_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_11_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_11_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_11_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_11_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_11_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_11_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_11_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_11_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_11_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_11_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_11_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_11_io_uop_uopc),
    .io_uop_inst                    (_slots_11_io_uop_inst),
    .io_uop_debug_inst              (_slots_11_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_11_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_11_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_11_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_11_io_uop_fu_code),
    .io_uop_iw_state                (_slots_11_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_11_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_11_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_11_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_11_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_11_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_11_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_11_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_11_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_11_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_11_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_11_io_uop_pc_lob),
    .io_uop_taken                   (_slots_11_io_uop_taken),
    .io_uop_imm_packed              (_slots_11_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_11_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_11_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_11_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_11_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_11_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_11_io_uop_pdst),
    .io_uop_prs1                    (_slots_11_io_uop_prs1),
    .io_uop_prs2                    (_slots_11_io_uop_prs2),
    .io_uop_prs3                    (_slots_11_io_uop_prs3),
    .io_uop_ppred                   (_slots_11_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_11_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_11_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_11_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_11_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_11_io_uop_stale_pdst),
    .io_uop_exception               (_slots_11_io_uop_exception),
    .io_uop_exc_cause               (_slots_11_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_11_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_11_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_11_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_11_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_11_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_11_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_11_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_11_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_11_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_11_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_11_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_11_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_11_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_11_io_uop_ldst),
    .io_uop_lrs1                    (_slots_11_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_11_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_11_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_11_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_11_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_11_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_11_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_11_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_11_io_uop_fp_val),
    .io_uop_fp_single               (_slots_11_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_11_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_11_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_11_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_11_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_11_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_11_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_11_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_12 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_12_io_valid),
    .io_will_be_valid               (_slots_12_io_will_be_valid),
    .io_request                     (_slots_12_io_request),
    .io_grant                       (issue_slots_12_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_11),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_12_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_57 ? _slots_16_io_out_uop_uopc : _GEN_56 ? _slots_15_io_out_uop_uopc : _GEN_55 ? _slots_14_io_out_uop_uopc : _slots_13_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_57 ? _slots_16_io_out_uop_inst : _GEN_56 ? _slots_15_io_out_uop_inst : _GEN_55 ? _slots_14_io_out_uop_inst : _slots_13_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_57 ? _slots_16_io_out_uop_debug_inst : _GEN_56 ? _slots_15_io_out_uop_debug_inst : _GEN_55 ? _slots_14_io_out_uop_debug_inst : _slots_13_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_57 ? _slots_16_io_out_uop_is_rvc : _GEN_56 ? _slots_15_io_out_uop_is_rvc : _GEN_55 ? _slots_14_io_out_uop_is_rvc : _slots_13_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_57 ? _slots_16_io_out_uop_debug_pc : _GEN_56 ? _slots_15_io_out_uop_debug_pc : _GEN_55 ? _slots_14_io_out_uop_debug_pc : _slots_13_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_57 ? _slots_16_io_out_uop_iq_type : _GEN_56 ? _slots_15_io_out_uop_iq_type : _GEN_55 ? _slots_14_io_out_uop_iq_type : _slots_13_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_57 ? _slots_16_io_out_uop_fu_code : _GEN_56 ? _slots_15_io_out_uop_fu_code : _GEN_55 ? _slots_14_io_out_uop_fu_code : _slots_13_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_57 ? _slots_16_io_out_uop_iw_state : _GEN_56 ? _slots_15_io_out_uop_iw_state : _GEN_55 ? _slots_14_io_out_uop_iw_state : _slots_13_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_57 ? _slots_16_io_out_uop_iw_p1_poisoned : _GEN_56 ? _slots_15_io_out_uop_iw_p1_poisoned : _GEN_55 ? _slots_14_io_out_uop_iw_p1_poisoned : _slots_13_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_57 ? _slots_16_io_out_uop_iw_p2_poisoned : _GEN_56 ? _slots_15_io_out_uop_iw_p2_poisoned : _GEN_55 ? _slots_14_io_out_uop_iw_p2_poisoned : _slots_13_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_57 ? _slots_16_io_out_uop_is_br : _GEN_56 ? _slots_15_io_out_uop_is_br : _GEN_55 ? _slots_14_io_out_uop_is_br : _slots_13_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_57 ? _slots_16_io_out_uop_is_jalr : _GEN_56 ? _slots_15_io_out_uop_is_jalr : _GEN_55 ? _slots_14_io_out_uop_is_jalr : _slots_13_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_57 ? _slots_16_io_out_uop_is_jal : _GEN_56 ? _slots_15_io_out_uop_is_jal : _GEN_55 ? _slots_14_io_out_uop_is_jal : _slots_13_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_57 ? _slots_16_io_out_uop_is_sfb : _GEN_56 ? _slots_15_io_out_uop_is_sfb : _GEN_55 ? _slots_14_io_out_uop_is_sfb : _slots_13_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_57 ? _slots_16_io_out_uop_br_mask : _GEN_56 ? _slots_15_io_out_uop_br_mask : _GEN_55 ? _slots_14_io_out_uop_br_mask : _slots_13_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_57 ? _slots_16_io_out_uop_br_tag : _GEN_56 ? _slots_15_io_out_uop_br_tag : _GEN_55 ? _slots_14_io_out_uop_br_tag : _slots_13_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_57 ? _slots_16_io_out_uop_ftq_idx : _GEN_56 ? _slots_15_io_out_uop_ftq_idx : _GEN_55 ? _slots_14_io_out_uop_ftq_idx : _slots_13_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_57 ? _slots_16_io_out_uop_edge_inst : _GEN_56 ? _slots_15_io_out_uop_edge_inst : _GEN_55 ? _slots_14_io_out_uop_edge_inst : _slots_13_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_57 ? _slots_16_io_out_uop_pc_lob : _GEN_56 ? _slots_15_io_out_uop_pc_lob : _GEN_55 ? _slots_14_io_out_uop_pc_lob : _slots_13_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_57 ? _slots_16_io_out_uop_taken : _GEN_56 ? _slots_15_io_out_uop_taken : _GEN_55 ? _slots_14_io_out_uop_taken : _slots_13_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_57 ? _slots_16_io_out_uop_imm_packed : _GEN_56 ? _slots_15_io_out_uop_imm_packed : _GEN_55 ? _slots_14_io_out_uop_imm_packed : _slots_13_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_57 ? _slots_16_io_out_uop_csr_addr : _GEN_56 ? _slots_15_io_out_uop_csr_addr : _GEN_55 ? _slots_14_io_out_uop_csr_addr : _slots_13_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_57 ? _slots_16_io_out_uop_rob_idx : _GEN_56 ? _slots_15_io_out_uop_rob_idx : _GEN_55 ? _slots_14_io_out_uop_rob_idx : _slots_13_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_57 ? _slots_16_io_out_uop_ldq_idx : _GEN_56 ? _slots_15_io_out_uop_ldq_idx : _GEN_55 ? _slots_14_io_out_uop_ldq_idx : _slots_13_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_57 ? _slots_16_io_out_uop_stq_idx : _GEN_56 ? _slots_15_io_out_uop_stq_idx : _GEN_55 ? _slots_14_io_out_uop_stq_idx : _slots_13_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_57 ? _slots_16_io_out_uop_rxq_idx : _GEN_56 ? _slots_15_io_out_uop_rxq_idx : _GEN_55 ? _slots_14_io_out_uop_rxq_idx : _slots_13_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_57 ? _slots_16_io_out_uop_pdst : _GEN_56 ? _slots_15_io_out_uop_pdst : _GEN_55 ? _slots_14_io_out_uop_pdst : _slots_13_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_57 ? _slots_16_io_out_uop_prs1 : _GEN_56 ? _slots_15_io_out_uop_prs1 : _GEN_55 ? _slots_14_io_out_uop_prs1 : _slots_13_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_57 ? _slots_16_io_out_uop_prs2 : _GEN_56 ? _slots_15_io_out_uop_prs2 : _GEN_55 ? _slots_14_io_out_uop_prs2 : _slots_13_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_57 ? _slots_16_io_out_uop_prs3 : _GEN_56 ? _slots_15_io_out_uop_prs3 : _GEN_55 ? _slots_14_io_out_uop_prs3 : _slots_13_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_57 ? _slots_16_io_out_uop_ppred : _GEN_56 ? _slots_15_io_out_uop_ppred : _GEN_55 ? _slots_14_io_out_uop_ppred : _slots_13_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_57 ? _slots_16_io_out_uop_prs1_busy : _GEN_56 ? _slots_15_io_out_uop_prs1_busy : _GEN_55 ? _slots_14_io_out_uop_prs1_busy : _slots_13_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_57 ? _slots_16_io_out_uop_prs2_busy : _GEN_56 ? _slots_15_io_out_uop_prs2_busy : _GEN_55 ? _slots_14_io_out_uop_prs2_busy : _slots_13_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_57 ? _slots_16_io_out_uop_prs3_busy : _GEN_56 ? _slots_15_io_out_uop_prs3_busy : _GEN_55 ? _slots_14_io_out_uop_prs3_busy : _slots_13_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_57 ? _slots_16_io_out_uop_ppred_busy : _GEN_56 ? _slots_15_io_out_uop_ppred_busy : _GEN_55 ? _slots_14_io_out_uop_ppred_busy : _slots_13_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_57 ? _slots_16_io_out_uop_stale_pdst : _GEN_56 ? _slots_15_io_out_uop_stale_pdst : _GEN_55 ? _slots_14_io_out_uop_stale_pdst : _slots_13_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_57 ? _slots_16_io_out_uop_exception : _GEN_56 ? _slots_15_io_out_uop_exception : _GEN_55 ? _slots_14_io_out_uop_exception : _slots_13_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_57 ? _slots_16_io_out_uop_exc_cause : _GEN_56 ? _slots_15_io_out_uop_exc_cause : _GEN_55 ? _slots_14_io_out_uop_exc_cause : _slots_13_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_57 ? _slots_16_io_out_uop_bypassable : _GEN_56 ? _slots_15_io_out_uop_bypassable : _GEN_55 ? _slots_14_io_out_uop_bypassable : _slots_13_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_57 ? _slots_16_io_out_uop_mem_cmd : _GEN_56 ? _slots_15_io_out_uop_mem_cmd : _GEN_55 ? _slots_14_io_out_uop_mem_cmd : _slots_13_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_57 ? _slots_16_io_out_uop_mem_size : _GEN_56 ? _slots_15_io_out_uop_mem_size : _GEN_55 ? _slots_14_io_out_uop_mem_size : _slots_13_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_57 ? _slots_16_io_out_uop_mem_signed : _GEN_56 ? _slots_15_io_out_uop_mem_signed : _GEN_55 ? _slots_14_io_out_uop_mem_signed : _slots_13_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_57 ? _slots_16_io_out_uop_is_fence : _GEN_56 ? _slots_15_io_out_uop_is_fence : _GEN_55 ? _slots_14_io_out_uop_is_fence : _slots_13_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_57 ? _slots_16_io_out_uop_is_fencei : _GEN_56 ? _slots_15_io_out_uop_is_fencei : _GEN_55 ? _slots_14_io_out_uop_is_fencei : _slots_13_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_57 ? _slots_16_io_out_uop_is_amo : _GEN_56 ? _slots_15_io_out_uop_is_amo : _GEN_55 ? _slots_14_io_out_uop_is_amo : _slots_13_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_57 ? _slots_16_io_out_uop_uses_ldq : _GEN_56 ? _slots_15_io_out_uop_uses_ldq : _GEN_55 ? _slots_14_io_out_uop_uses_ldq : _slots_13_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_57 ? _slots_16_io_out_uop_uses_stq : _GEN_56 ? _slots_15_io_out_uop_uses_stq : _GEN_55 ? _slots_14_io_out_uop_uses_stq : _slots_13_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_57 ? _slots_16_io_out_uop_is_sys_pc2epc : _GEN_56 ? _slots_15_io_out_uop_is_sys_pc2epc : _GEN_55 ? _slots_14_io_out_uop_is_sys_pc2epc : _slots_13_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_57 ? _slots_16_io_out_uop_is_unique : _GEN_56 ? _slots_15_io_out_uop_is_unique : _GEN_55 ? _slots_14_io_out_uop_is_unique : _slots_13_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_57 ? _slots_16_io_out_uop_flush_on_commit : _GEN_56 ? _slots_15_io_out_uop_flush_on_commit : _GEN_55 ? _slots_14_io_out_uop_flush_on_commit : _slots_13_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_57 ? _slots_16_io_out_uop_ldst_is_rs1 : _GEN_56 ? _slots_15_io_out_uop_ldst_is_rs1 : _GEN_55 ? _slots_14_io_out_uop_ldst_is_rs1 : _slots_13_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_57 ? _slots_16_io_out_uop_ldst : _GEN_56 ? _slots_15_io_out_uop_ldst : _GEN_55 ? _slots_14_io_out_uop_ldst : _slots_13_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_57 ? _slots_16_io_out_uop_lrs1 : _GEN_56 ? _slots_15_io_out_uop_lrs1 : _GEN_55 ? _slots_14_io_out_uop_lrs1 : _slots_13_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_57 ? _slots_16_io_out_uop_lrs2 : _GEN_56 ? _slots_15_io_out_uop_lrs2 : _GEN_55 ? _slots_14_io_out_uop_lrs2 : _slots_13_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_57 ? _slots_16_io_out_uop_lrs3 : _GEN_56 ? _slots_15_io_out_uop_lrs3 : _GEN_55 ? _slots_14_io_out_uop_lrs3 : _slots_13_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_57 ? _slots_16_io_out_uop_ldst_val : _GEN_56 ? _slots_15_io_out_uop_ldst_val : _GEN_55 ? _slots_14_io_out_uop_ldst_val : _slots_13_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_57 ? _slots_16_io_out_uop_dst_rtype : _GEN_56 ? _slots_15_io_out_uop_dst_rtype : _GEN_55 ? _slots_14_io_out_uop_dst_rtype : _slots_13_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_57 ? _slots_16_io_out_uop_lrs1_rtype : _GEN_56 ? _slots_15_io_out_uop_lrs1_rtype : _GEN_55 ? _slots_14_io_out_uop_lrs1_rtype : _slots_13_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_57 ? _slots_16_io_out_uop_lrs2_rtype : _GEN_56 ? _slots_15_io_out_uop_lrs2_rtype : _GEN_55 ? _slots_14_io_out_uop_lrs2_rtype : _slots_13_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_57 ? _slots_16_io_out_uop_frs3_en : _GEN_56 ? _slots_15_io_out_uop_frs3_en : _GEN_55 ? _slots_14_io_out_uop_frs3_en : _slots_13_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_57 ? _slots_16_io_out_uop_fp_val : _GEN_56 ? _slots_15_io_out_uop_fp_val : _GEN_55 ? _slots_14_io_out_uop_fp_val : _slots_13_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_57 ? _slots_16_io_out_uop_fp_single : _GEN_56 ? _slots_15_io_out_uop_fp_single : _GEN_55 ? _slots_14_io_out_uop_fp_single : _slots_13_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_57 ? _slots_16_io_out_uop_xcpt_pf_if : _GEN_56 ? _slots_15_io_out_uop_xcpt_pf_if : _GEN_55 ? _slots_14_io_out_uop_xcpt_pf_if : _slots_13_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_57 ? _slots_16_io_out_uop_xcpt_ae_if : _GEN_56 ? _slots_15_io_out_uop_xcpt_ae_if : _GEN_55 ? _slots_14_io_out_uop_xcpt_ae_if : _slots_13_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_57 ? _slots_16_io_out_uop_xcpt_ma_if : _GEN_56 ? _slots_15_io_out_uop_xcpt_ma_if : _GEN_55 ? _slots_14_io_out_uop_xcpt_ma_if : _slots_13_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_57 ? _slots_16_io_out_uop_bp_debug_if : _GEN_56 ? _slots_15_io_out_uop_bp_debug_if : _GEN_55 ? _slots_14_io_out_uop_bp_debug_if : _slots_13_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_57 ? _slots_16_io_out_uop_bp_xcpt_if : _GEN_56 ? _slots_15_io_out_uop_bp_xcpt_if : _GEN_55 ? _slots_14_io_out_uop_bp_xcpt_if : _slots_13_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_57 ? _slots_16_io_out_uop_debug_fsrc : _GEN_56 ? _slots_15_io_out_uop_debug_fsrc : _GEN_55 ? _slots_14_io_out_uop_debug_fsrc : _slots_13_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_57 ? _slots_16_io_out_uop_debug_tsrc : _GEN_56 ? _slots_15_io_out_uop_debug_tsrc : _GEN_55 ? _slots_14_io_out_uop_debug_tsrc : _slots_13_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_12_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_12_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_12_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_12_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_12_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_12_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_12_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_12_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_12_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_12_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_12_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_12_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_12_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_12_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_12_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_12_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_12_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_12_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_12_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_12_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_12_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_12_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_12_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_12_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_12_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_12_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_12_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_12_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_12_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_12_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_12_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_12_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_12_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_12_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_12_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_12_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_12_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_12_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_12_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_12_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_12_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_12_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_12_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_12_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_12_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_12_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_12_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_12_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_12_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_12_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_12_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_12_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_12_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_12_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_12_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_12_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_12_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_12_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_12_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_12_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_12_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_12_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_12_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_12_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_12_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_12_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_12_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_12_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_12_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_12_io_uop_uopc),
    .io_uop_inst                    (_slots_12_io_uop_inst),
    .io_uop_debug_inst              (_slots_12_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_12_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_12_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_12_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_12_io_uop_fu_code),
    .io_uop_iw_state                (_slots_12_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_12_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_12_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_12_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_12_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_12_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_12_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_12_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_12_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_12_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_12_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_12_io_uop_pc_lob),
    .io_uop_taken                   (_slots_12_io_uop_taken),
    .io_uop_imm_packed              (_slots_12_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_12_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_12_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_12_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_12_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_12_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_12_io_uop_pdst),
    .io_uop_prs1                    (_slots_12_io_uop_prs1),
    .io_uop_prs2                    (_slots_12_io_uop_prs2),
    .io_uop_prs3                    (_slots_12_io_uop_prs3),
    .io_uop_ppred                   (_slots_12_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_12_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_12_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_12_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_12_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_12_io_uop_stale_pdst),
    .io_uop_exception               (_slots_12_io_uop_exception),
    .io_uop_exc_cause               (_slots_12_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_12_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_12_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_12_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_12_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_12_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_12_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_12_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_12_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_12_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_12_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_12_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_12_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_12_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_12_io_uop_ldst),
    .io_uop_lrs1                    (_slots_12_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_12_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_12_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_12_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_12_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_12_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_12_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_12_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_12_io_uop_fp_val),
    .io_uop_fp_single               (_slots_12_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_12_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_12_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_12_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_12_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_12_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_12_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_12_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_13 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_13_io_valid),
    .io_will_be_valid               (_slots_13_io_will_be_valid),
    .io_request                     (_slots_13_io_request),
    .io_grant                       (issue_slots_13_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_12),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_13_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_60 ? _slots_17_io_out_uop_uopc : _GEN_59 ? _slots_16_io_out_uop_uopc : _GEN_58 ? _slots_15_io_out_uop_uopc : _slots_14_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_60 ? _slots_17_io_out_uop_inst : _GEN_59 ? _slots_16_io_out_uop_inst : _GEN_58 ? _slots_15_io_out_uop_inst : _slots_14_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_60 ? _slots_17_io_out_uop_debug_inst : _GEN_59 ? _slots_16_io_out_uop_debug_inst : _GEN_58 ? _slots_15_io_out_uop_debug_inst : _slots_14_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_60 ? _slots_17_io_out_uop_is_rvc : _GEN_59 ? _slots_16_io_out_uop_is_rvc : _GEN_58 ? _slots_15_io_out_uop_is_rvc : _slots_14_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_60 ? _slots_17_io_out_uop_debug_pc : _GEN_59 ? _slots_16_io_out_uop_debug_pc : _GEN_58 ? _slots_15_io_out_uop_debug_pc : _slots_14_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_60 ? _slots_17_io_out_uop_iq_type : _GEN_59 ? _slots_16_io_out_uop_iq_type : _GEN_58 ? _slots_15_io_out_uop_iq_type : _slots_14_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_60 ? _slots_17_io_out_uop_fu_code : _GEN_59 ? _slots_16_io_out_uop_fu_code : _GEN_58 ? _slots_15_io_out_uop_fu_code : _slots_14_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_60 ? _slots_17_io_out_uop_iw_state : _GEN_59 ? _slots_16_io_out_uop_iw_state : _GEN_58 ? _slots_15_io_out_uop_iw_state : _slots_14_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_60 ? _slots_17_io_out_uop_iw_p1_poisoned : _GEN_59 ? _slots_16_io_out_uop_iw_p1_poisoned : _GEN_58 ? _slots_15_io_out_uop_iw_p1_poisoned : _slots_14_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_60 ? _slots_17_io_out_uop_iw_p2_poisoned : _GEN_59 ? _slots_16_io_out_uop_iw_p2_poisoned : _GEN_58 ? _slots_15_io_out_uop_iw_p2_poisoned : _slots_14_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_60 ? _slots_17_io_out_uop_is_br : _GEN_59 ? _slots_16_io_out_uop_is_br : _GEN_58 ? _slots_15_io_out_uop_is_br : _slots_14_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_60 ? _slots_17_io_out_uop_is_jalr : _GEN_59 ? _slots_16_io_out_uop_is_jalr : _GEN_58 ? _slots_15_io_out_uop_is_jalr : _slots_14_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_60 ? _slots_17_io_out_uop_is_jal : _GEN_59 ? _slots_16_io_out_uop_is_jal : _GEN_58 ? _slots_15_io_out_uop_is_jal : _slots_14_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_60 ? _slots_17_io_out_uop_is_sfb : _GEN_59 ? _slots_16_io_out_uop_is_sfb : _GEN_58 ? _slots_15_io_out_uop_is_sfb : _slots_14_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_60 ? _slots_17_io_out_uop_br_mask : _GEN_59 ? _slots_16_io_out_uop_br_mask : _GEN_58 ? _slots_15_io_out_uop_br_mask : _slots_14_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_60 ? _slots_17_io_out_uop_br_tag : _GEN_59 ? _slots_16_io_out_uop_br_tag : _GEN_58 ? _slots_15_io_out_uop_br_tag : _slots_14_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_60 ? _slots_17_io_out_uop_ftq_idx : _GEN_59 ? _slots_16_io_out_uop_ftq_idx : _GEN_58 ? _slots_15_io_out_uop_ftq_idx : _slots_14_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_60 ? _slots_17_io_out_uop_edge_inst : _GEN_59 ? _slots_16_io_out_uop_edge_inst : _GEN_58 ? _slots_15_io_out_uop_edge_inst : _slots_14_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_60 ? _slots_17_io_out_uop_pc_lob : _GEN_59 ? _slots_16_io_out_uop_pc_lob : _GEN_58 ? _slots_15_io_out_uop_pc_lob : _slots_14_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_60 ? _slots_17_io_out_uop_taken : _GEN_59 ? _slots_16_io_out_uop_taken : _GEN_58 ? _slots_15_io_out_uop_taken : _slots_14_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_60 ? _slots_17_io_out_uop_imm_packed : _GEN_59 ? _slots_16_io_out_uop_imm_packed : _GEN_58 ? _slots_15_io_out_uop_imm_packed : _slots_14_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_60 ? _slots_17_io_out_uop_csr_addr : _GEN_59 ? _slots_16_io_out_uop_csr_addr : _GEN_58 ? _slots_15_io_out_uop_csr_addr : _slots_14_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_60 ? _slots_17_io_out_uop_rob_idx : _GEN_59 ? _slots_16_io_out_uop_rob_idx : _GEN_58 ? _slots_15_io_out_uop_rob_idx : _slots_14_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_60 ? _slots_17_io_out_uop_ldq_idx : _GEN_59 ? _slots_16_io_out_uop_ldq_idx : _GEN_58 ? _slots_15_io_out_uop_ldq_idx : _slots_14_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_60 ? _slots_17_io_out_uop_stq_idx : _GEN_59 ? _slots_16_io_out_uop_stq_idx : _GEN_58 ? _slots_15_io_out_uop_stq_idx : _slots_14_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_60 ? _slots_17_io_out_uop_rxq_idx : _GEN_59 ? _slots_16_io_out_uop_rxq_idx : _GEN_58 ? _slots_15_io_out_uop_rxq_idx : _slots_14_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_60 ? _slots_17_io_out_uop_pdst : _GEN_59 ? _slots_16_io_out_uop_pdst : _GEN_58 ? _slots_15_io_out_uop_pdst : _slots_14_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_60 ? _slots_17_io_out_uop_prs1 : _GEN_59 ? _slots_16_io_out_uop_prs1 : _GEN_58 ? _slots_15_io_out_uop_prs1 : _slots_14_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_60 ? _slots_17_io_out_uop_prs2 : _GEN_59 ? _slots_16_io_out_uop_prs2 : _GEN_58 ? _slots_15_io_out_uop_prs2 : _slots_14_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_60 ? _slots_17_io_out_uop_prs3 : _GEN_59 ? _slots_16_io_out_uop_prs3 : _GEN_58 ? _slots_15_io_out_uop_prs3 : _slots_14_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_60 ? _slots_17_io_out_uop_ppred : _GEN_59 ? _slots_16_io_out_uop_ppred : _GEN_58 ? _slots_15_io_out_uop_ppred : _slots_14_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_60 ? _slots_17_io_out_uop_prs1_busy : _GEN_59 ? _slots_16_io_out_uop_prs1_busy : _GEN_58 ? _slots_15_io_out_uop_prs1_busy : _slots_14_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_60 ? _slots_17_io_out_uop_prs2_busy : _GEN_59 ? _slots_16_io_out_uop_prs2_busy : _GEN_58 ? _slots_15_io_out_uop_prs2_busy : _slots_14_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_60 ? _slots_17_io_out_uop_prs3_busy : _GEN_59 ? _slots_16_io_out_uop_prs3_busy : _GEN_58 ? _slots_15_io_out_uop_prs3_busy : _slots_14_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_60 ? _slots_17_io_out_uop_ppred_busy : _GEN_59 ? _slots_16_io_out_uop_ppred_busy : _GEN_58 ? _slots_15_io_out_uop_ppred_busy : _slots_14_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_60 ? _slots_17_io_out_uop_stale_pdst : _GEN_59 ? _slots_16_io_out_uop_stale_pdst : _GEN_58 ? _slots_15_io_out_uop_stale_pdst : _slots_14_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_60 ? _slots_17_io_out_uop_exception : _GEN_59 ? _slots_16_io_out_uop_exception : _GEN_58 ? _slots_15_io_out_uop_exception : _slots_14_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_60 ? _slots_17_io_out_uop_exc_cause : _GEN_59 ? _slots_16_io_out_uop_exc_cause : _GEN_58 ? _slots_15_io_out_uop_exc_cause : _slots_14_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_60 ? _slots_17_io_out_uop_bypassable : _GEN_59 ? _slots_16_io_out_uop_bypassable : _GEN_58 ? _slots_15_io_out_uop_bypassable : _slots_14_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_60 ? _slots_17_io_out_uop_mem_cmd : _GEN_59 ? _slots_16_io_out_uop_mem_cmd : _GEN_58 ? _slots_15_io_out_uop_mem_cmd : _slots_14_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_60 ? _slots_17_io_out_uop_mem_size : _GEN_59 ? _slots_16_io_out_uop_mem_size : _GEN_58 ? _slots_15_io_out_uop_mem_size : _slots_14_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_60 ? _slots_17_io_out_uop_mem_signed : _GEN_59 ? _slots_16_io_out_uop_mem_signed : _GEN_58 ? _slots_15_io_out_uop_mem_signed : _slots_14_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_60 ? _slots_17_io_out_uop_is_fence : _GEN_59 ? _slots_16_io_out_uop_is_fence : _GEN_58 ? _slots_15_io_out_uop_is_fence : _slots_14_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_60 ? _slots_17_io_out_uop_is_fencei : _GEN_59 ? _slots_16_io_out_uop_is_fencei : _GEN_58 ? _slots_15_io_out_uop_is_fencei : _slots_14_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_60 ? _slots_17_io_out_uop_is_amo : _GEN_59 ? _slots_16_io_out_uop_is_amo : _GEN_58 ? _slots_15_io_out_uop_is_amo : _slots_14_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_60 ? _slots_17_io_out_uop_uses_ldq : _GEN_59 ? _slots_16_io_out_uop_uses_ldq : _GEN_58 ? _slots_15_io_out_uop_uses_ldq : _slots_14_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_60 ? _slots_17_io_out_uop_uses_stq : _GEN_59 ? _slots_16_io_out_uop_uses_stq : _GEN_58 ? _slots_15_io_out_uop_uses_stq : _slots_14_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_60 ? _slots_17_io_out_uop_is_sys_pc2epc : _GEN_59 ? _slots_16_io_out_uop_is_sys_pc2epc : _GEN_58 ? _slots_15_io_out_uop_is_sys_pc2epc : _slots_14_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_60 ? _slots_17_io_out_uop_is_unique : _GEN_59 ? _slots_16_io_out_uop_is_unique : _GEN_58 ? _slots_15_io_out_uop_is_unique : _slots_14_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_60 ? _slots_17_io_out_uop_flush_on_commit : _GEN_59 ? _slots_16_io_out_uop_flush_on_commit : _GEN_58 ? _slots_15_io_out_uop_flush_on_commit : _slots_14_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_60 ? _slots_17_io_out_uop_ldst_is_rs1 : _GEN_59 ? _slots_16_io_out_uop_ldst_is_rs1 : _GEN_58 ? _slots_15_io_out_uop_ldst_is_rs1 : _slots_14_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_60 ? _slots_17_io_out_uop_ldst : _GEN_59 ? _slots_16_io_out_uop_ldst : _GEN_58 ? _slots_15_io_out_uop_ldst : _slots_14_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_60 ? _slots_17_io_out_uop_lrs1 : _GEN_59 ? _slots_16_io_out_uop_lrs1 : _GEN_58 ? _slots_15_io_out_uop_lrs1 : _slots_14_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_60 ? _slots_17_io_out_uop_lrs2 : _GEN_59 ? _slots_16_io_out_uop_lrs2 : _GEN_58 ? _slots_15_io_out_uop_lrs2 : _slots_14_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_60 ? _slots_17_io_out_uop_lrs3 : _GEN_59 ? _slots_16_io_out_uop_lrs3 : _GEN_58 ? _slots_15_io_out_uop_lrs3 : _slots_14_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_60 ? _slots_17_io_out_uop_ldst_val : _GEN_59 ? _slots_16_io_out_uop_ldst_val : _GEN_58 ? _slots_15_io_out_uop_ldst_val : _slots_14_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_60 ? _slots_17_io_out_uop_dst_rtype : _GEN_59 ? _slots_16_io_out_uop_dst_rtype : _GEN_58 ? _slots_15_io_out_uop_dst_rtype : _slots_14_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_60 ? _slots_17_io_out_uop_lrs1_rtype : _GEN_59 ? _slots_16_io_out_uop_lrs1_rtype : _GEN_58 ? _slots_15_io_out_uop_lrs1_rtype : _slots_14_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_60 ? _slots_17_io_out_uop_lrs2_rtype : _GEN_59 ? _slots_16_io_out_uop_lrs2_rtype : _GEN_58 ? _slots_15_io_out_uop_lrs2_rtype : _slots_14_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_60 ? _slots_17_io_out_uop_frs3_en : _GEN_59 ? _slots_16_io_out_uop_frs3_en : _GEN_58 ? _slots_15_io_out_uop_frs3_en : _slots_14_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_60 ? _slots_17_io_out_uop_fp_val : _GEN_59 ? _slots_16_io_out_uop_fp_val : _GEN_58 ? _slots_15_io_out_uop_fp_val : _slots_14_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_60 ? _slots_17_io_out_uop_fp_single : _GEN_59 ? _slots_16_io_out_uop_fp_single : _GEN_58 ? _slots_15_io_out_uop_fp_single : _slots_14_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_60 ? _slots_17_io_out_uop_xcpt_pf_if : _GEN_59 ? _slots_16_io_out_uop_xcpt_pf_if : _GEN_58 ? _slots_15_io_out_uop_xcpt_pf_if : _slots_14_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_60 ? _slots_17_io_out_uop_xcpt_ae_if : _GEN_59 ? _slots_16_io_out_uop_xcpt_ae_if : _GEN_58 ? _slots_15_io_out_uop_xcpt_ae_if : _slots_14_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_60 ? _slots_17_io_out_uop_xcpt_ma_if : _GEN_59 ? _slots_16_io_out_uop_xcpt_ma_if : _GEN_58 ? _slots_15_io_out_uop_xcpt_ma_if : _slots_14_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_60 ? _slots_17_io_out_uop_bp_debug_if : _GEN_59 ? _slots_16_io_out_uop_bp_debug_if : _GEN_58 ? _slots_15_io_out_uop_bp_debug_if : _slots_14_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_60 ? _slots_17_io_out_uop_bp_xcpt_if : _GEN_59 ? _slots_16_io_out_uop_bp_xcpt_if : _GEN_58 ? _slots_15_io_out_uop_bp_xcpt_if : _slots_14_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_60 ? _slots_17_io_out_uop_debug_fsrc : _GEN_59 ? _slots_16_io_out_uop_debug_fsrc : _GEN_58 ? _slots_15_io_out_uop_debug_fsrc : _slots_14_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_60 ? _slots_17_io_out_uop_debug_tsrc : _GEN_59 ? _slots_16_io_out_uop_debug_tsrc : _GEN_58 ? _slots_15_io_out_uop_debug_tsrc : _slots_14_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_13_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_13_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_13_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_13_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_13_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_13_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_13_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_13_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_13_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_13_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_13_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_13_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_13_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_13_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_13_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_13_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_13_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_13_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_13_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_13_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_13_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_13_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_13_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_13_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_13_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_13_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_13_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_13_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_13_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_13_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_13_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_13_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_13_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_13_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_13_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_13_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_13_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_13_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_13_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_13_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_13_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_13_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_13_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_13_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_13_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_13_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_13_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_13_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_13_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_13_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_13_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_13_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_13_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_13_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_13_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_13_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_13_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_13_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_13_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_13_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_13_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_13_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_13_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_13_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_13_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_13_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_13_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_13_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_13_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_13_io_uop_uopc),
    .io_uop_inst                    (_slots_13_io_uop_inst),
    .io_uop_debug_inst              (_slots_13_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_13_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_13_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_13_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_13_io_uop_fu_code),
    .io_uop_iw_state                (_slots_13_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_13_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_13_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_13_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_13_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_13_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_13_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_13_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_13_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_13_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_13_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_13_io_uop_pc_lob),
    .io_uop_taken                   (_slots_13_io_uop_taken),
    .io_uop_imm_packed              (_slots_13_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_13_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_13_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_13_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_13_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_13_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_13_io_uop_pdst),
    .io_uop_prs1                    (_slots_13_io_uop_prs1),
    .io_uop_prs2                    (_slots_13_io_uop_prs2),
    .io_uop_prs3                    (_slots_13_io_uop_prs3),
    .io_uop_ppred                   (_slots_13_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_13_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_13_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_13_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_13_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_13_io_uop_stale_pdst),
    .io_uop_exception               (_slots_13_io_uop_exception),
    .io_uop_exc_cause               (_slots_13_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_13_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_13_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_13_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_13_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_13_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_13_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_13_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_13_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_13_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_13_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_13_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_13_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_13_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_13_io_uop_ldst),
    .io_uop_lrs1                    (_slots_13_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_13_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_13_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_13_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_13_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_13_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_13_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_13_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_13_io_uop_fp_val),
    .io_uop_fp_single               (_slots_13_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_13_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_13_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_13_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_13_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_13_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_13_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_13_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_14 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_14_io_valid),
    .io_will_be_valid               (_slots_14_io_will_be_valid),
    .io_request                     (_slots_14_io_request),
    .io_grant                       (issue_slots_14_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_13),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_14_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_63 ? _slots_18_io_out_uop_uopc : _GEN_62 ? _slots_17_io_out_uop_uopc : _GEN_61 ? _slots_16_io_out_uop_uopc : _slots_15_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_63 ? _slots_18_io_out_uop_inst : _GEN_62 ? _slots_17_io_out_uop_inst : _GEN_61 ? _slots_16_io_out_uop_inst : _slots_15_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_63 ? _slots_18_io_out_uop_debug_inst : _GEN_62 ? _slots_17_io_out_uop_debug_inst : _GEN_61 ? _slots_16_io_out_uop_debug_inst : _slots_15_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_63 ? _slots_18_io_out_uop_is_rvc : _GEN_62 ? _slots_17_io_out_uop_is_rvc : _GEN_61 ? _slots_16_io_out_uop_is_rvc : _slots_15_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_63 ? _slots_18_io_out_uop_debug_pc : _GEN_62 ? _slots_17_io_out_uop_debug_pc : _GEN_61 ? _slots_16_io_out_uop_debug_pc : _slots_15_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_63 ? _slots_18_io_out_uop_iq_type : _GEN_62 ? _slots_17_io_out_uop_iq_type : _GEN_61 ? _slots_16_io_out_uop_iq_type : _slots_15_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_63 ? _slots_18_io_out_uop_fu_code : _GEN_62 ? _slots_17_io_out_uop_fu_code : _GEN_61 ? _slots_16_io_out_uop_fu_code : _slots_15_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_63 ? _slots_18_io_out_uop_iw_state : _GEN_62 ? _slots_17_io_out_uop_iw_state : _GEN_61 ? _slots_16_io_out_uop_iw_state : _slots_15_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_63 ? _slots_18_io_out_uop_iw_p1_poisoned : _GEN_62 ? _slots_17_io_out_uop_iw_p1_poisoned : _GEN_61 ? _slots_16_io_out_uop_iw_p1_poisoned : _slots_15_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_63 ? _slots_18_io_out_uop_iw_p2_poisoned : _GEN_62 ? _slots_17_io_out_uop_iw_p2_poisoned : _GEN_61 ? _slots_16_io_out_uop_iw_p2_poisoned : _slots_15_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_63 ? _slots_18_io_out_uop_is_br : _GEN_62 ? _slots_17_io_out_uop_is_br : _GEN_61 ? _slots_16_io_out_uop_is_br : _slots_15_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_63 ? _slots_18_io_out_uop_is_jalr : _GEN_62 ? _slots_17_io_out_uop_is_jalr : _GEN_61 ? _slots_16_io_out_uop_is_jalr : _slots_15_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_63 ? _slots_18_io_out_uop_is_jal : _GEN_62 ? _slots_17_io_out_uop_is_jal : _GEN_61 ? _slots_16_io_out_uop_is_jal : _slots_15_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_63 ? _slots_18_io_out_uop_is_sfb : _GEN_62 ? _slots_17_io_out_uop_is_sfb : _GEN_61 ? _slots_16_io_out_uop_is_sfb : _slots_15_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_63 ? _slots_18_io_out_uop_br_mask : _GEN_62 ? _slots_17_io_out_uop_br_mask : _GEN_61 ? _slots_16_io_out_uop_br_mask : _slots_15_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_63 ? _slots_18_io_out_uop_br_tag : _GEN_62 ? _slots_17_io_out_uop_br_tag : _GEN_61 ? _slots_16_io_out_uop_br_tag : _slots_15_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_63 ? _slots_18_io_out_uop_ftq_idx : _GEN_62 ? _slots_17_io_out_uop_ftq_idx : _GEN_61 ? _slots_16_io_out_uop_ftq_idx : _slots_15_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_63 ? _slots_18_io_out_uop_edge_inst : _GEN_62 ? _slots_17_io_out_uop_edge_inst : _GEN_61 ? _slots_16_io_out_uop_edge_inst : _slots_15_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_63 ? _slots_18_io_out_uop_pc_lob : _GEN_62 ? _slots_17_io_out_uop_pc_lob : _GEN_61 ? _slots_16_io_out_uop_pc_lob : _slots_15_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_63 ? _slots_18_io_out_uop_taken : _GEN_62 ? _slots_17_io_out_uop_taken : _GEN_61 ? _slots_16_io_out_uop_taken : _slots_15_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_63 ? _slots_18_io_out_uop_imm_packed : _GEN_62 ? _slots_17_io_out_uop_imm_packed : _GEN_61 ? _slots_16_io_out_uop_imm_packed : _slots_15_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_63 ? _slots_18_io_out_uop_csr_addr : _GEN_62 ? _slots_17_io_out_uop_csr_addr : _GEN_61 ? _slots_16_io_out_uop_csr_addr : _slots_15_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_63 ? _slots_18_io_out_uop_rob_idx : _GEN_62 ? _slots_17_io_out_uop_rob_idx : _GEN_61 ? _slots_16_io_out_uop_rob_idx : _slots_15_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_63 ? _slots_18_io_out_uop_ldq_idx : _GEN_62 ? _slots_17_io_out_uop_ldq_idx : _GEN_61 ? _slots_16_io_out_uop_ldq_idx : _slots_15_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_63 ? _slots_18_io_out_uop_stq_idx : _GEN_62 ? _slots_17_io_out_uop_stq_idx : _GEN_61 ? _slots_16_io_out_uop_stq_idx : _slots_15_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_63 ? _slots_18_io_out_uop_rxq_idx : _GEN_62 ? _slots_17_io_out_uop_rxq_idx : _GEN_61 ? _slots_16_io_out_uop_rxq_idx : _slots_15_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_63 ? _slots_18_io_out_uop_pdst : _GEN_62 ? _slots_17_io_out_uop_pdst : _GEN_61 ? _slots_16_io_out_uop_pdst : _slots_15_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_63 ? _slots_18_io_out_uop_prs1 : _GEN_62 ? _slots_17_io_out_uop_prs1 : _GEN_61 ? _slots_16_io_out_uop_prs1 : _slots_15_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_63 ? _slots_18_io_out_uop_prs2 : _GEN_62 ? _slots_17_io_out_uop_prs2 : _GEN_61 ? _slots_16_io_out_uop_prs2 : _slots_15_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_63 ? _slots_18_io_out_uop_prs3 : _GEN_62 ? _slots_17_io_out_uop_prs3 : _GEN_61 ? _slots_16_io_out_uop_prs3 : _slots_15_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_63 ? _slots_18_io_out_uop_ppred : _GEN_62 ? _slots_17_io_out_uop_ppred : _GEN_61 ? _slots_16_io_out_uop_ppred : _slots_15_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_63 ? _slots_18_io_out_uop_prs1_busy : _GEN_62 ? _slots_17_io_out_uop_prs1_busy : _GEN_61 ? _slots_16_io_out_uop_prs1_busy : _slots_15_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_63 ? _slots_18_io_out_uop_prs2_busy : _GEN_62 ? _slots_17_io_out_uop_prs2_busy : _GEN_61 ? _slots_16_io_out_uop_prs2_busy : _slots_15_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_63 ? _slots_18_io_out_uop_prs3_busy : _GEN_62 ? _slots_17_io_out_uop_prs3_busy : _GEN_61 ? _slots_16_io_out_uop_prs3_busy : _slots_15_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_63 ? _slots_18_io_out_uop_ppred_busy : _GEN_62 ? _slots_17_io_out_uop_ppred_busy : _GEN_61 ? _slots_16_io_out_uop_ppred_busy : _slots_15_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_63 ? _slots_18_io_out_uop_stale_pdst : _GEN_62 ? _slots_17_io_out_uop_stale_pdst : _GEN_61 ? _slots_16_io_out_uop_stale_pdst : _slots_15_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_63 ? _slots_18_io_out_uop_exception : _GEN_62 ? _slots_17_io_out_uop_exception : _GEN_61 ? _slots_16_io_out_uop_exception : _slots_15_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_63 ? _slots_18_io_out_uop_exc_cause : _GEN_62 ? _slots_17_io_out_uop_exc_cause : _GEN_61 ? _slots_16_io_out_uop_exc_cause : _slots_15_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_63 ? _slots_18_io_out_uop_bypassable : _GEN_62 ? _slots_17_io_out_uop_bypassable : _GEN_61 ? _slots_16_io_out_uop_bypassable : _slots_15_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_63 ? _slots_18_io_out_uop_mem_cmd : _GEN_62 ? _slots_17_io_out_uop_mem_cmd : _GEN_61 ? _slots_16_io_out_uop_mem_cmd : _slots_15_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_63 ? _slots_18_io_out_uop_mem_size : _GEN_62 ? _slots_17_io_out_uop_mem_size : _GEN_61 ? _slots_16_io_out_uop_mem_size : _slots_15_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_63 ? _slots_18_io_out_uop_mem_signed : _GEN_62 ? _slots_17_io_out_uop_mem_signed : _GEN_61 ? _slots_16_io_out_uop_mem_signed : _slots_15_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_63 ? _slots_18_io_out_uop_is_fence : _GEN_62 ? _slots_17_io_out_uop_is_fence : _GEN_61 ? _slots_16_io_out_uop_is_fence : _slots_15_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_63 ? _slots_18_io_out_uop_is_fencei : _GEN_62 ? _slots_17_io_out_uop_is_fencei : _GEN_61 ? _slots_16_io_out_uop_is_fencei : _slots_15_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_63 ? _slots_18_io_out_uop_is_amo : _GEN_62 ? _slots_17_io_out_uop_is_amo : _GEN_61 ? _slots_16_io_out_uop_is_amo : _slots_15_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_63 ? _slots_18_io_out_uop_uses_ldq : _GEN_62 ? _slots_17_io_out_uop_uses_ldq : _GEN_61 ? _slots_16_io_out_uop_uses_ldq : _slots_15_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_63 ? _slots_18_io_out_uop_uses_stq : _GEN_62 ? _slots_17_io_out_uop_uses_stq : _GEN_61 ? _slots_16_io_out_uop_uses_stq : _slots_15_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_63 ? _slots_18_io_out_uop_is_sys_pc2epc : _GEN_62 ? _slots_17_io_out_uop_is_sys_pc2epc : _GEN_61 ? _slots_16_io_out_uop_is_sys_pc2epc : _slots_15_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_63 ? _slots_18_io_out_uop_is_unique : _GEN_62 ? _slots_17_io_out_uop_is_unique : _GEN_61 ? _slots_16_io_out_uop_is_unique : _slots_15_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_63 ? _slots_18_io_out_uop_flush_on_commit : _GEN_62 ? _slots_17_io_out_uop_flush_on_commit : _GEN_61 ? _slots_16_io_out_uop_flush_on_commit : _slots_15_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_63 ? _slots_18_io_out_uop_ldst_is_rs1 : _GEN_62 ? _slots_17_io_out_uop_ldst_is_rs1 : _GEN_61 ? _slots_16_io_out_uop_ldst_is_rs1 : _slots_15_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_63 ? _slots_18_io_out_uop_ldst : _GEN_62 ? _slots_17_io_out_uop_ldst : _GEN_61 ? _slots_16_io_out_uop_ldst : _slots_15_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_63 ? _slots_18_io_out_uop_lrs1 : _GEN_62 ? _slots_17_io_out_uop_lrs1 : _GEN_61 ? _slots_16_io_out_uop_lrs1 : _slots_15_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_63 ? _slots_18_io_out_uop_lrs2 : _GEN_62 ? _slots_17_io_out_uop_lrs2 : _GEN_61 ? _slots_16_io_out_uop_lrs2 : _slots_15_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_63 ? _slots_18_io_out_uop_lrs3 : _GEN_62 ? _slots_17_io_out_uop_lrs3 : _GEN_61 ? _slots_16_io_out_uop_lrs3 : _slots_15_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_63 ? _slots_18_io_out_uop_ldst_val : _GEN_62 ? _slots_17_io_out_uop_ldst_val : _GEN_61 ? _slots_16_io_out_uop_ldst_val : _slots_15_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_63 ? _slots_18_io_out_uop_dst_rtype : _GEN_62 ? _slots_17_io_out_uop_dst_rtype : _GEN_61 ? _slots_16_io_out_uop_dst_rtype : _slots_15_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_63 ? _slots_18_io_out_uop_lrs1_rtype : _GEN_62 ? _slots_17_io_out_uop_lrs1_rtype : _GEN_61 ? _slots_16_io_out_uop_lrs1_rtype : _slots_15_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_63 ? _slots_18_io_out_uop_lrs2_rtype : _GEN_62 ? _slots_17_io_out_uop_lrs2_rtype : _GEN_61 ? _slots_16_io_out_uop_lrs2_rtype : _slots_15_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_63 ? _slots_18_io_out_uop_frs3_en : _GEN_62 ? _slots_17_io_out_uop_frs3_en : _GEN_61 ? _slots_16_io_out_uop_frs3_en : _slots_15_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_63 ? _slots_18_io_out_uop_fp_val : _GEN_62 ? _slots_17_io_out_uop_fp_val : _GEN_61 ? _slots_16_io_out_uop_fp_val : _slots_15_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_63 ? _slots_18_io_out_uop_fp_single : _GEN_62 ? _slots_17_io_out_uop_fp_single : _GEN_61 ? _slots_16_io_out_uop_fp_single : _slots_15_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_63 ? _slots_18_io_out_uop_xcpt_pf_if : _GEN_62 ? _slots_17_io_out_uop_xcpt_pf_if : _GEN_61 ? _slots_16_io_out_uop_xcpt_pf_if : _slots_15_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_63 ? _slots_18_io_out_uop_xcpt_ae_if : _GEN_62 ? _slots_17_io_out_uop_xcpt_ae_if : _GEN_61 ? _slots_16_io_out_uop_xcpt_ae_if : _slots_15_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_63 ? _slots_18_io_out_uop_xcpt_ma_if : _GEN_62 ? _slots_17_io_out_uop_xcpt_ma_if : _GEN_61 ? _slots_16_io_out_uop_xcpt_ma_if : _slots_15_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_63 ? _slots_18_io_out_uop_bp_debug_if : _GEN_62 ? _slots_17_io_out_uop_bp_debug_if : _GEN_61 ? _slots_16_io_out_uop_bp_debug_if : _slots_15_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_63 ? _slots_18_io_out_uop_bp_xcpt_if : _GEN_62 ? _slots_17_io_out_uop_bp_xcpt_if : _GEN_61 ? _slots_16_io_out_uop_bp_xcpt_if : _slots_15_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_63 ? _slots_18_io_out_uop_debug_fsrc : _GEN_62 ? _slots_17_io_out_uop_debug_fsrc : _GEN_61 ? _slots_16_io_out_uop_debug_fsrc : _slots_15_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_63 ? _slots_18_io_out_uop_debug_tsrc : _GEN_62 ? _slots_17_io_out_uop_debug_tsrc : _GEN_61 ? _slots_16_io_out_uop_debug_tsrc : _slots_15_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_14_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_14_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_14_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_14_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_14_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_14_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_14_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_14_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_14_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_14_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_14_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_14_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_14_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_14_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_14_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_14_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_14_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_14_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_14_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_14_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_14_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_14_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_14_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_14_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_14_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_14_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_14_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_14_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_14_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_14_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_14_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_14_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_14_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_14_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_14_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_14_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_14_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_14_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_14_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_14_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_14_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_14_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_14_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_14_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_14_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_14_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_14_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_14_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_14_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_14_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_14_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_14_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_14_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_14_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_14_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_14_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_14_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_14_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_14_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_14_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_14_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_14_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_14_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_14_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_14_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_14_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_14_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_14_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_14_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_14_io_uop_uopc),
    .io_uop_inst                    (_slots_14_io_uop_inst),
    .io_uop_debug_inst              (_slots_14_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_14_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_14_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_14_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_14_io_uop_fu_code),
    .io_uop_iw_state                (_slots_14_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_14_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_14_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_14_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_14_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_14_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_14_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_14_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_14_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_14_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_14_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_14_io_uop_pc_lob),
    .io_uop_taken                   (_slots_14_io_uop_taken),
    .io_uop_imm_packed              (_slots_14_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_14_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_14_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_14_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_14_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_14_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_14_io_uop_pdst),
    .io_uop_prs1                    (_slots_14_io_uop_prs1),
    .io_uop_prs2                    (_slots_14_io_uop_prs2),
    .io_uop_prs3                    (_slots_14_io_uop_prs3),
    .io_uop_ppred                   (_slots_14_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_14_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_14_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_14_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_14_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_14_io_uop_stale_pdst),
    .io_uop_exception               (_slots_14_io_uop_exception),
    .io_uop_exc_cause               (_slots_14_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_14_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_14_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_14_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_14_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_14_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_14_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_14_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_14_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_14_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_14_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_14_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_14_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_14_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_14_io_uop_ldst),
    .io_uop_lrs1                    (_slots_14_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_14_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_14_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_14_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_14_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_14_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_14_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_14_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_14_io_uop_fp_val),
    .io_uop_fp_single               (_slots_14_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_14_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_14_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_14_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_14_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_14_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_14_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_14_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_15 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_15_io_valid),
    .io_will_be_valid               (_slots_15_io_will_be_valid),
    .io_request                     (_slots_15_io_request),
    .io_grant                       (issue_slots_15_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_14),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_15_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_66 ? _slots_19_io_out_uop_uopc : _GEN_65 ? _slots_18_io_out_uop_uopc : _GEN_64 ? _slots_17_io_out_uop_uopc : _slots_16_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_66 ? _slots_19_io_out_uop_inst : _GEN_65 ? _slots_18_io_out_uop_inst : _GEN_64 ? _slots_17_io_out_uop_inst : _slots_16_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_66 ? _slots_19_io_out_uop_debug_inst : _GEN_65 ? _slots_18_io_out_uop_debug_inst : _GEN_64 ? _slots_17_io_out_uop_debug_inst : _slots_16_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_66 ? _slots_19_io_out_uop_is_rvc : _GEN_65 ? _slots_18_io_out_uop_is_rvc : _GEN_64 ? _slots_17_io_out_uop_is_rvc : _slots_16_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_66 ? _slots_19_io_out_uop_debug_pc : _GEN_65 ? _slots_18_io_out_uop_debug_pc : _GEN_64 ? _slots_17_io_out_uop_debug_pc : _slots_16_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_66 ? _slots_19_io_out_uop_iq_type : _GEN_65 ? _slots_18_io_out_uop_iq_type : _GEN_64 ? _slots_17_io_out_uop_iq_type : _slots_16_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_66 ? _slots_19_io_out_uop_fu_code : _GEN_65 ? _slots_18_io_out_uop_fu_code : _GEN_64 ? _slots_17_io_out_uop_fu_code : _slots_16_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_66 ? _slots_19_io_out_uop_iw_state : _GEN_65 ? _slots_18_io_out_uop_iw_state : _GEN_64 ? _slots_17_io_out_uop_iw_state : _slots_16_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_66 ? _slots_19_io_out_uop_iw_p1_poisoned : _GEN_65 ? _slots_18_io_out_uop_iw_p1_poisoned : _GEN_64 ? _slots_17_io_out_uop_iw_p1_poisoned : _slots_16_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_66 ? _slots_19_io_out_uop_iw_p2_poisoned : _GEN_65 ? _slots_18_io_out_uop_iw_p2_poisoned : _GEN_64 ? _slots_17_io_out_uop_iw_p2_poisoned : _slots_16_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_66 ? _slots_19_io_out_uop_is_br : _GEN_65 ? _slots_18_io_out_uop_is_br : _GEN_64 ? _slots_17_io_out_uop_is_br : _slots_16_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_66 ? _slots_19_io_out_uop_is_jalr : _GEN_65 ? _slots_18_io_out_uop_is_jalr : _GEN_64 ? _slots_17_io_out_uop_is_jalr : _slots_16_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_66 ? _slots_19_io_out_uop_is_jal : _GEN_65 ? _slots_18_io_out_uop_is_jal : _GEN_64 ? _slots_17_io_out_uop_is_jal : _slots_16_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_66 ? _slots_19_io_out_uop_is_sfb : _GEN_65 ? _slots_18_io_out_uop_is_sfb : _GEN_64 ? _slots_17_io_out_uop_is_sfb : _slots_16_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_66 ? _slots_19_io_out_uop_br_mask : _GEN_65 ? _slots_18_io_out_uop_br_mask : _GEN_64 ? _slots_17_io_out_uop_br_mask : _slots_16_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_66 ? _slots_19_io_out_uop_br_tag : _GEN_65 ? _slots_18_io_out_uop_br_tag : _GEN_64 ? _slots_17_io_out_uop_br_tag : _slots_16_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_66 ? _slots_19_io_out_uop_ftq_idx : _GEN_65 ? _slots_18_io_out_uop_ftq_idx : _GEN_64 ? _slots_17_io_out_uop_ftq_idx : _slots_16_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_66 ? _slots_19_io_out_uop_edge_inst : _GEN_65 ? _slots_18_io_out_uop_edge_inst : _GEN_64 ? _slots_17_io_out_uop_edge_inst : _slots_16_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_66 ? _slots_19_io_out_uop_pc_lob : _GEN_65 ? _slots_18_io_out_uop_pc_lob : _GEN_64 ? _slots_17_io_out_uop_pc_lob : _slots_16_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_66 ? _slots_19_io_out_uop_taken : _GEN_65 ? _slots_18_io_out_uop_taken : _GEN_64 ? _slots_17_io_out_uop_taken : _slots_16_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_66 ? _slots_19_io_out_uop_imm_packed : _GEN_65 ? _slots_18_io_out_uop_imm_packed : _GEN_64 ? _slots_17_io_out_uop_imm_packed : _slots_16_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_66 ? _slots_19_io_out_uop_csr_addr : _GEN_65 ? _slots_18_io_out_uop_csr_addr : _GEN_64 ? _slots_17_io_out_uop_csr_addr : _slots_16_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_66 ? _slots_19_io_out_uop_rob_idx : _GEN_65 ? _slots_18_io_out_uop_rob_idx : _GEN_64 ? _slots_17_io_out_uop_rob_idx : _slots_16_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_66 ? _slots_19_io_out_uop_ldq_idx : _GEN_65 ? _slots_18_io_out_uop_ldq_idx : _GEN_64 ? _slots_17_io_out_uop_ldq_idx : _slots_16_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_66 ? _slots_19_io_out_uop_stq_idx : _GEN_65 ? _slots_18_io_out_uop_stq_idx : _GEN_64 ? _slots_17_io_out_uop_stq_idx : _slots_16_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_66 ? _slots_19_io_out_uop_rxq_idx : _GEN_65 ? _slots_18_io_out_uop_rxq_idx : _GEN_64 ? _slots_17_io_out_uop_rxq_idx : _slots_16_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_66 ? _slots_19_io_out_uop_pdst : _GEN_65 ? _slots_18_io_out_uop_pdst : _GEN_64 ? _slots_17_io_out_uop_pdst : _slots_16_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_66 ? _slots_19_io_out_uop_prs1 : _GEN_65 ? _slots_18_io_out_uop_prs1 : _GEN_64 ? _slots_17_io_out_uop_prs1 : _slots_16_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_66 ? _slots_19_io_out_uop_prs2 : _GEN_65 ? _slots_18_io_out_uop_prs2 : _GEN_64 ? _slots_17_io_out_uop_prs2 : _slots_16_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_66 ? _slots_19_io_out_uop_prs3 : _GEN_65 ? _slots_18_io_out_uop_prs3 : _GEN_64 ? _slots_17_io_out_uop_prs3 : _slots_16_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_66 ? _slots_19_io_out_uop_ppred : _GEN_65 ? _slots_18_io_out_uop_ppred : _GEN_64 ? _slots_17_io_out_uop_ppred : _slots_16_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_66 ? _slots_19_io_out_uop_prs1_busy : _GEN_65 ? _slots_18_io_out_uop_prs1_busy : _GEN_64 ? _slots_17_io_out_uop_prs1_busy : _slots_16_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_66 ? _slots_19_io_out_uop_prs2_busy : _GEN_65 ? _slots_18_io_out_uop_prs2_busy : _GEN_64 ? _slots_17_io_out_uop_prs2_busy : _slots_16_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_66 ? _slots_19_io_out_uop_prs3_busy : _GEN_65 ? _slots_18_io_out_uop_prs3_busy : _GEN_64 ? _slots_17_io_out_uop_prs3_busy : _slots_16_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_66 ? _slots_19_io_out_uop_ppred_busy : _GEN_65 ? _slots_18_io_out_uop_ppred_busy : _GEN_64 ? _slots_17_io_out_uop_ppred_busy : _slots_16_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_66 ? _slots_19_io_out_uop_stale_pdst : _GEN_65 ? _slots_18_io_out_uop_stale_pdst : _GEN_64 ? _slots_17_io_out_uop_stale_pdst : _slots_16_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_66 ? _slots_19_io_out_uop_exception : _GEN_65 ? _slots_18_io_out_uop_exception : _GEN_64 ? _slots_17_io_out_uop_exception : _slots_16_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_66 ? _slots_19_io_out_uop_exc_cause : _GEN_65 ? _slots_18_io_out_uop_exc_cause : _GEN_64 ? _slots_17_io_out_uop_exc_cause : _slots_16_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_66 ? _slots_19_io_out_uop_bypassable : _GEN_65 ? _slots_18_io_out_uop_bypassable : _GEN_64 ? _slots_17_io_out_uop_bypassable : _slots_16_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_66 ? _slots_19_io_out_uop_mem_cmd : _GEN_65 ? _slots_18_io_out_uop_mem_cmd : _GEN_64 ? _slots_17_io_out_uop_mem_cmd : _slots_16_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_66 ? _slots_19_io_out_uop_mem_size : _GEN_65 ? _slots_18_io_out_uop_mem_size : _GEN_64 ? _slots_17_io_out_uop_mem_size : _slots_16_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_66 ? _slots_19_io_out_uop_mem_signed : _GEN_65 ? _slots_18_io_out_uop_mem_signed : _GEN_64 ? _slots_17_io_out_uop_mem_signed : _slots_16_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_66 ? _slots_19_io_out_uop_is_fence : _GEN_65 ? _slots_18_io_out_uop_is_fence : _GEN_64 ? _slots_17_io_out_uop_is_fence : _slots_16_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_66 ? _slots_19_io_out_uop_is_fencei : _GEN_65 ? _slots_18_io_out_uop_is_fencei : _GEN_64 ? _slots_17_io_out_uop_is_fencei : _slots_16_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_66 ? _slots_19_io_out_uop_is_amo : _GEN_65 ? _slots_18_io_out_uop_is_amo : _GEN_64 ? _slots_17_io_out_uop_is_amo : _slots_16_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_66 ? _slots_19_io_out_uop_uses_ldq : _GEN_65 ? _slots_18_io_out_uop_uses_ldq : _GEN_64 ? _slots_17_io_out_uop_uses_ldq : _slots_16_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_66 ? _slots_19_io_out_uop_uses_stq : _GEN_65 ? _slots_18_io_out_uop_uses_stq : _GEN_64 ? _slots_17_io_out_uop_uses_stq : _slots_16_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_66 ? _slots_19_io_out_uop_is_sys_pc2epc : _GEN_65 ? _slots_18_io_out_uop_is_sys_pc2epc : _GEN_64 ? _slots_17_io_out_uop_is_sys_pc2epc : _slots_16_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_66 ? _slots_19_io_out_uop_is_unique : _GEN_65 ? _slots_18_io_out_uop_is_unique : _GEN_64 ? _slots_17_io_out_uop_is_unique : _slots_16_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_66 ? _slots_19_io_out_uop_flush_on_commit : _GEN_65 ? _slots_18_io_out_uop_flush_on_commit : _GEN_64 ? _slots_17_io_out_uop_flush_on_commit : _slots_16_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_66 ? _slots_19_io_out_uop_ldst_is_rs1 : _GEN_65 ? _slots_18_io_out_uop_ldst_is_rs1 : _GEN_64 ? _slots_17_io_out_uop_ldst_is_rs1 : _slots_16_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_66 ? _slots_19_io_out_uop_ldst : _GEN_65 ? _slots_18_io_out_uop_ldst : _GEN_64 ? _slots_17_io_out_uop_ldst : _slots_16_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_66 ? _slots_19_io_out_uop_lrs1 : _GEN_65 ? _slots_18_io_out_uop_lrs1 : _GEN_64 ? _slots_17_io_out_uop_lrs1 : _slots_16_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_66 ? _slots_19_io_out_uop_lrs2 : _GEN_65 ? _slots_18_io_out_uop_lrs2 : _GEN_64 ? _slots_17_io_out_uop_lrs2 : _slots_16_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_66 ? _slots_19_io_out_uop_lrs3 : _GEN_65 ? _slots_18_io_out_uop_lrs3 : _GEN_64 ? _slots_17_io_out_uop_lrs3 : _slots_16_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_66 ? _slots_19_io_out_uop_ldst_val : _GEN_65 ? _slots_18_io_out_uop_ldst_val : _GEN_64 ? _slots_17_io_out_uop_ldst_val : _slots_16_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_66 ? _slots_19_io_out_uop_dst_rtype : _GEN_65 ? _slots_18_io_out_uop_dst_rtype : _GEN_64 ? _slots_17_io_out_uop_dst_rtype : _slots_16_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_66 ? _slots_19_io_out_uop_lrs1_rtype : _GEN_65 ? _slots_18_io_out_uop_lrs1_rtype : _GEN_64 ? _slots_17_io_out_uop_lrs1_rtype : _slots_16_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_66 ? _slots_19_io_out_uop_lrs2_rtype : _GEN_65 ? _slots_18_io_out_uop_lrs2_rtype : _GEN_64 ? _slots_17_io_out_uop_lrs2_rtype : _slots_16_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_66 ? _slots_19_io_out_uop_frs3_en : _GEN_65 ? _slots_18_io_out_uop_frs3_en : _GEN_64 ? _slots_17_io_out_uop_frs3_en : _slots_16_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_66 ? _slots_19_io_out_uop_fp_val : _GEN_65 ? _slots_18_io_out_uop_fp_val : _GEN_64 ? _slots_17_io_out_uop_fp_val : _slots_16_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_66 ? _slots_19_io_out_uop_fp_single : _GEN_65 ? _slots_18_io_out_uop_fp_single : _GEN_64 ? _slots_17_io_out_uop_fp_single : _slots_16_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_66 ? _slots_19_io_out_uop_xcpt_pf_if : _GEN_65 ? _slots_18_io_out_uop_xcpt_pf_if : _GEN_64 ? _slots_17_io_out_uop_xcpt_pf_if : _slots_16_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_66 ? _slots_19_io_out_uop_xcpt_ae_if : _GEN_65 ? _slots_18_io_out_uop_xcpt_ae_if : _GEN_64 ? _slots_17_io_out_uop_xcpt_ae_if : _slots_16_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_66 ? _slots_19_io_out_uop_xcpt_ma_if : _GEN_65 ? _slots_18_io_out_uop_xcpt_ma_if : _GEN_64 ? _slots_17_io_out_uop_xcpt_ma_if : _slots_16_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_66 ? _slots_19_io_out_uop_bp_debug_if : _GEN_65 ? _slots_18_io_out_uop_bp_debug_if : _GEN_64 ? _slots_17_io_out_uop_bp_debug_if : _slots_16_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_66 ? _slots_19_io_out_uop_bp_xcpt_if : _GEN_65 ? _slots_18_io_out_uop_bp_xcpt_if : _GEN_64 ? _slots_17_io_out_uop_bp_xcpt_if : _slots_16_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_66 ? _slots_19_io_out_uop_debug_fsrc : _GEN_65 ? _slots_18_io_out_uop_debug_fsrc : _GEN_64 ? _slots_17_io_out_uop_debug_fsrc : _slots_16_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_66 ? _slots_19_io_out_uop_debug_tsrc : _GEN_65 ? _slots_18_io_out_uop_debug_tsrc : _GEN_64 ? _slots_17_io_out_uop_debug_tsrc : _slots_16_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_15_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_15_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_15_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_15_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_15_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_15_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_15_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_15_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_15_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_15_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_15_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_15_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_15_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_15_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_15_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_15_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_15_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_15_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_15_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_15_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_15_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_15_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_15_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_15_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_15_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_15_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_15_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_15_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_15_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_15_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_15_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_15_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_15_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_15_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_15_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_15_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_15_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_15_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_15_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_15_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_15_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_15_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_15_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_15_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_15_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_15_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_15_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_15_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_15_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_15_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_15_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_15_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_15_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_15_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_15_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_15_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_15_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_15_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_15_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_15_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_15_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_15_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_15_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_15_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_15_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_15_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_15_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_15_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_15_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_15_io_uop_uopc),
    .io_uop_inst                    (_slots_15_io_uop_inst),
    .io_uop_debug_inst              (_slots_15_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_15_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_15_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_15_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_15_io_uop_fu_code),
    .io_uop_iw_state                (_slots_15_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_15_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_15_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_15_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_15_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_15_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_15_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_15_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_15_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_15_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_15_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_15_io_uop_pc_lob),
    .io_uop_taken                   (_slots_15_io_uop_taken),
    .io_uop_imm_packed              (_slots_15_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_15_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_15_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_15_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_15_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_15_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_15_io_uop_pdst),
    .io_uop_prs1                    (_slots_15_io_uop_prs1),
    .io_uop_prs2                    (_slots_15_io_uop_prs2),
    .io_uop_prs3                    (_slots_15_io_uop_prs3),
    .io_uop_ppred                   (_slots_15_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_15_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_15_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_15_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_15_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_15_io_uop_stale_pdst),
    .io_uop_exception               (_slots_15_io_uop_exception),
    .io_uop_exc_cause               (_slots_15_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_15_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_15_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_15_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_15_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_15_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_15_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_15_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_15_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_15_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_15_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_15_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_15_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_15_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_15_io_uop_ldst),
    .io_uop_lrs1                    (_slots_15_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_15_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_15_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_15_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_15_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_15_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_15_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_15_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_15_io_uop_fp_val),
    .io_uop_fp_single               (_slots_15_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_15_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_15_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_15_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_15_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_15_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_15_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_15_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_16 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_16_io_valid),
    .io_will_be_valid               (_slots_16_io_will_be_valid),
    .io_request                     (_slots_16_io_request),
    .io_grant                       (issue_slots_16_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_15),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_16_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_69 ? _slots_20_io_out_uop_uopc : _GEN_68 ? _slots_19_io_out_uop_uopc : _GEN_67 ? _slots_18_io_out_uop_uopc : _slots_17_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_69 ? _slots_20_io_out_uop_inst : _GEN_68 ? _slots_19_io_out_uop_inst : _GEN_67 ? _slots_18_io_out_uop_inst : _slots_17_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_69 ? _slots_20_io_out_uop_debug_inst : _GEN_68 ? _slots_19_io_out_uop_debug_inst : _GEN_67 ? _slots_18_io_out_uop_debug_inst : _slots_17_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_69 ? _slots_20_io_out_uop_is_rvc : _GEN_68 ? _slots_19_io_out_uop_is_rvc : _GEN_67 ? _slots_18_io_out_uop_is_rvc : _slots_17_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_69 ? _slots_20_io_out_uop_debug_pc : _GEN_68 ? _slots_19_io_out_uop_debug_pc : _GEN_67 ? _slots_18_io_out_uop_debug_pc : _slots_17_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_69 ? _slots_20_io_out_uop_iq_type : _GEN_68 ? _slots_19_io_out_uop_iq_type : _GEN_67 ? _slots_18_io_out_uop_iq_type : _slots_17_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_69 ? _slots_20_io_out_uop_fu_code : _GEN_68 ? _slots_19_io_out_uop_fu_code : _GEN_67 ? _slots_18_io_out_uop_fu_code : _slots_17_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_69 ? _slots_20_io_out_uop_iw_state : _GEN_68 ? _slots_19_io_out_uop_iw_state : _GEN_67 ? _slots_18_io_out_uop_iw_state : _slots_17_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_69 ? _slots_20_io_out_uop_iw_p1_poisoned : _GEN_68 ? _slots_19_io_out_uop_iw_p1_poisoned : _GEN_67 ? _slots_18_io_out_uop_iw_p1_poisoned : _slots_17_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_69 ? _slots_20_io_out_uop_iw_p2_poisoned : _GEN_68 ? _slots_19_io_out_uop_iw_p2_poisoned : _GEN_67 ? _slots_18_io_out_uop_iw_p2_poisoned : _slots_17_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_69 ? _slots_20_io_out_uop_is_br : _GEN_68 ? _slots_19_io_out_uop_is_br : _GEN_67 ? _slots_18_io_out_uop_is_br : _slots_17_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_69 ? _slots_20_io_out_uop_is_jalr : _GEN_68 ? _slots_19_io_out_uop_is_jalr : _GEN_67 ? _slots_18_io_out_uop_is_jalr : _slots_17_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_69 ? _slots_20_io_out_uop_is_jal : _GEN_68 ? _slots_19_io_out_uop_is_jal : _GEN_67 ? _slots_18_io_out_uop_is_jal : _slots_17_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_69 ? _slots_20_io_out_uop_is_sfb : _GEN_68 ? _slots_19_io_out_uop_is_sfb : _GEN_67 ? _slots_18_io_out_uop_is_sfb : _slots_17_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_69 ? _slots_20_io_out_uop_br_mask : _GEN_68 ? _slots_19_io_out_uop_br_mask : _GEN_67 ? _slots_18_io_out_uop_br_mask : _slots_17_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_69 ? _slots_20_io_out_uop_br_tag : _GEN_68 ? _slots_19_io_out_uop_br_tag : _GEN_67 ? _slots_18_io_out_uop_br_tag : _slots_17_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_69 ? _slots_20_io_out_uop_ftq_idx : _GEN_68 ? _slots_19_io_out_uop_ftq_idx : _GEN_67 ? _slots_18_io_out_uop_ftq_idx : _slots_17_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_69 ? _slots_20_io_out_uop_edge_inst : _GEN_68 ? _slots_19_io_out_uop_edge_inst : _GEN_67 ? _slots_18_io_out_uop_edge_inst : _slots_17_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_69 ? _slots_20_io_out_uop_pc_lob : _GEN_68 ? _slots_19_io_out_uop_pc_lob : _GEN_67 ? _slots_18_io_out_uop_pc_lob : _slots_17_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_69 ? _slots_20_io_out_uop_taken : _GEN_68 ? _slots_19_io_out_uop_taken : _GEN_67 ? _slots_18_io_out_uop_taken : _slots_17_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_69 ? _slots_20_io_out_uop_imm_packed : _GEN_68 ? _slots_19_io_out_uop_imm_packed : _GEN_67 ? _slots_18_io_out_uop_imm_packed : _slots_17_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_69 ? _slots_20_io_out_uop_csr_addr : _GEN_68 ? _slots_19_io_out_uop_csr_addr : _GEN_67 ? _slots_18_io_out_uop_csr_addr : _slots_17_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_69 ? _slots_20_io_out_uop_rob_idx : _GEN_68 ? _slots_19_io_out_uop_rob_idx : _GEN_67 ? _slots_18_io_out_uop_rob_idx : _slots_17_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_69 ? _slots_20_io_out_uop_ldq_idx : _GEN_68 ? _slots_19_io_out_uop_ldq_idx : _GEN_67 ? _slots_18_io_out_uop_ldq_idx : _slots_17_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_69 ? _slots_20_io_out_uop_stq_idx : _GEN_68 ? _slots_19_io_out_uop_stq_idx : _GEN_67 ? _slots_18_io_out_uop_stq_idx : _slots_17_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_69 ? _slots_20_io_out_uop_rxq_idx : _GEN_68 ? _slots_19_io_out_uop_rxq_idx : _GEN_67 ? _slots_18_io_out_uop_rxq_idx : _slots_17_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_69 ? _slots_20_io_out_uop_pdst : _GEN_68 ? _slots_19_io_out_uop_pdst : _GEN_67 ? _slots_18_io_out_uop_pdst : _slots_17_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_69 ? _slots_20_io_out_uop_prs1 : _GEN_68 ? _slots_19_io_out_uop_prs1 : _GEN_67 ? _slots_18_io_out_uop_prs1 : _slots_17_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_69 ? _slots_20_io_out_uop_prs2 : _GEN_68 ? _slots_19_io_out_uop_prs2 : _GEN_67 ? _slots_18_io_out_uop_prs2 : _slots_17_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_69 ? _slots_20_io_out_uop_prs3 : _GEN_68 ? _slots_19_io_out_uop_prs3 : _GEN_67 ? _slots_18_io_out_uop_prs3 : _slots_17_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_69 ? _slots_20_io_out_uop_ppred : _GEN_68 ? _slots_19_io_out_uop_ppred : _GEN_67 ? _slots_18_io_out_uop_ppred : _slots_17_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_69 ? _slots_20_io_out_uop_prs1_busy : _GEN_68 ? _slots_19_io_out_uop_prs1_busy : _GEN_67 ? _slots_18_io_out_uop_prs1_busy : _slots_17_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_69 ? _slots_20_io_out_uop_prs2_busy : _GEN_68 ? _slots_19_io_out_uop_prs2_busy : _GEN_67 ? _slots_18_io_out_uop_prs2_busy : _slots_17_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_69 ? _slots_20_io_out_uop_prs3_busy : _GEN_68 ? _slots_19_io_out_uop_prs3_busy : _GEN_67 ? _slots_18_io_out_uop_prs3_busy : _slots_17_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_69 ? _slots_20_io_out_uop_ppred_busy : _GEN_68 ? _slots_19_io_out_uop_ppred_busy : _GEN_67 ? _slots_18_io_out_uop_ppred_busy : _slots_17_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_69 ? _slots_20_io_out_uop_stale_pdst : _GEN_68 ? _slots_19_io_out_uop_stale_pdst : _GEN_67 ? _slots_18_io_out_uop_stale_pdst : _slots_17_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_69 ? _slots_20_io_out_uop_exception : _GEN_68 ? _slots_19_io_out_uop_exception : _GEN_67 ? _slots_18_io_out_uop_exception : _slots_17_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_69 ? _slots_20_io_out_uop_exc_cause : _GEN_68 ? _slots_19_io_out_uop_exc_cause : _GEN_67 ? _slots_18_io_out_uop_exc_cause : _slots_17_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_69 ? _slots_20_io_out_uop_bypassable : _GEN_68 ? _slots_19_io_out_uop_bypassable : _GEN_67 ? _slots_18_io_out_uop_bypassable : _slots_17_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_69 ? _slots_20_io_out_uop_mem_cmd : _GEN_68 ? _slots_19_io_out_uop_mem_cmd : _GEN_67 ? _slots_18_io_out_uop_mem_cmd : _slots_17_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_69 ? _slots_20_io_out_uop_mem_size : _GEN_68 ? _slots_19_io_out_uop_mem_size : _GEN_67 ? _slots_18_io_out_uop_mem_size : _slots_17_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_69 ? _slots_20_io_out_uop_mem_signed : _GEN_68 ? _slots_19_io_out_uop_mem_signed : _GEN_67 ? _slots_18_io_out_uop_mem_signed : _slots_17_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_69 ? _slots_20_io_out_uop_is_fence : _GEN_68 ? _slots_19_io_out_uop_is_fence : _GEN_67 ? _slots_18_io_out_uop_is_fence : _slots_17_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_69 ? _slots_20_io_out_uop_is_fencei : _GEN_68 ? _slots_19_io_out_uop_is_fencei : _GEN_67 ? _slots_18_io_out_uop_is_fencei : _slots_17_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_69 ? _slots_20_io_out_uop_is_amo : _GEN_68 ? _slots_19_io_out_uop_is_amo : _GEN_67 ? _slots_18_io_out_uop_is_amo : _slots_17_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_69 ? _slots_20_io_out_uop_uses_ldq : _GEN_68 ? _slots_19_io_out_uop_uses_ldq : _GEN_67 ? _slots_18_io_out_uop_uses_ldq : _slots_17_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_69 ? _slots_20_io_out_uop_uses_stq : _GEN_68 ? _slots_19_io_out_uop_uses_stq : _GEN_67 ? _slots_18_io_out_uop_uses_stq : _slots_17_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_69 ? _slots_20_io_out_uop_is_sys_pc2epc : _GEN_68 ? _slots_19_io_out_uop_is_sys_pc2epc : _GEN_67 ? _slots_18_io_out_uop_is_sys_pc2epc : _slots_17_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_69 ? _slots_20_io_out_uop_is_unique : _GEN_68 ? _slots_19_io_out_uop_is_unique : _GEN_67 ? _slots_18_io_out_uop_is_unique : _slots_17_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_69 ? _slots_20_io_out_uop_flush_on_commit : _GEN_68 ? _slots_19_io_out_uop_flush_on_commit : _GEN_67 ? _slots_18_io_out_uop_flush_on_commit : _slots_17_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_69 ? _slots_20_io_out_uop_ldst_is_rs1 : _GEN_68 ? _slots_19_io_out_uop_ldst_is_rs1 : _GEN_67 ? _slots_18_io_out_uop_ldst_is_rs1 : _slots_17_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_69 ? _slots_20_io_out_uop_ldst : _GEN_68 ? _slots_19_io_out_uop_ldst : _GEN_67 ? _slots_18_io_out_uop_ldst : _slots_17_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_69 ? _slots_20_io_out_uop_lrs1 : _GEN_68 ? _slots_19_io_out_uop_lrs1 : _GEN_67 ? _slots_18_io_out_uop_lrs1 : _slots_17_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_69 ? _slots_20_io_out_uop_lrs2 : _GEN_68 ? _slots_19_io_out_uop_lrs2 : _GEN_67 ? _slots_18_io_out_uop_lrs2 : _slots_17_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_69 ? _slots_20_io_out_uop_lrs3 : _GEN_68 ? _slots_19_io_out_uop_lrs3 : _GEN_67 ? _slots_18_io_out_uop_lrs3 : _slots_17_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_69 ? _slots_20_io_out_uop_ldst_val : _GEN_68 ? _slots_19_io_out_uop_ldst_val : _GEN_67 ? _slots_18_io_out_uop_ldst_val : _slots_17_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_69 ? _slots_20_io_out_uop_dst_rtype : _GEN_68 ? _slots_19_io_out_uop_dst_rtype : _GEN_67 ? _slots_18_io_out_uop_dst_rtype : _slots_17_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_69 ? _slots_20_io_out_uop_lrs1_rtype : _GEN_68 ? _slots_19_io_out_uop_lrs1_rtype : _GEN_67 ? _slots_18_io_out_uop_lrs1_rtype : _slots_17_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_69 ? _slots_20_io_out_uop_lrs2_rtype : _GEN_68 ? _slots_19_io_out_uop_lrs2_rtype : _GEN_67 ? _slots_18_io_out_uop_lrs2_rtype : _slots_17_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_69 ? _slots_20_io_out_uop_frs3_en : _GEN_68 ? _slots_19_io_out_uop_frs3_en : _GEN_67 ? _slots_18_io_out_uop_frs3_en : _slots_17_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_69 ? _slots_20_io_out_uop_fp_val : _GEN_68 ? _slots_19_io_out_uop_fp_val : _GEN_67 ? _slots_18_io_out_uop_fp_val : _slots_17_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_69 ? _slots_20_io_out_uop_fp_single : _GEN_68 ? _slots_19_io_out_uop_fp_single : _GEN_67 ? _slots_18_io_out_uop_fp_single : _slots_17_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_69 ? _slots_20_io_out_uop_xcpt_pf_if : _GEN_68 ? _slots_19_io_out_uop_xcpt_pf_if : _GEN_67 ? _slots_18_io_out_uop_xcpt_pf_if : _slots_17_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_69 ? _slots_20_io_out_uop_xcpt_ae_if : _GEN_68 ? _slots_19_io_out_uop_xcpt_ae_if : _GEN_67 ? _slots_18_io_out_uop_xcpt_ae_if : _slots_17_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_69 ? _slots_20_io_out_uop_xcpt_ma_if : _GEN_68 ? _slots_19_io_out_uop_xcpt_ma_if : _GEN_67 ? _slots_18_io_out_uop_xcpt_ma_if : _slots_17_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_69 ? _slots_20_io_out_uop_bp_debug_if : _GEN_68 ? _slots_19_io_out_uop_bp_debug_if : _GEN_67 ? _slots_18_io_out_uop_bp_debug_if : _slots_17_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_69 ? _slots_20_io_out_uop_bp_xcpt_if : _GEN_68 ? _slots_19_io_out_uop_bp_xcpt_if : _GEN_67 ? _slots_18_io_out_uop_bp_xcpt_if : _slots_17_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_69 ? _slots_20_io_out_uop_debug_fsrc : _GEN_68 ? _slots_19_io_out_uop_debug_fsrc : _GEN_67 ? _slots_18_io_out_uop_debug_fsrc : _slots_17_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_69 ? _slots_20_io_out_uop_debug_tsrc : _GEN_68 ? _slots_19_io_out_uop_debug_tsrc : _GEN_67 ? _slots_18_io_out_uop_debug_tsrc : _slots_17_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_16_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_16_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_16_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_16_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_16_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_16_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_16_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_16_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_16_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_16_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_16_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_16_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_16_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_16_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_16_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_16_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_16_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_16_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_16_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_16_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_16_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_16_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_16_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_16_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_16_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_16_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_16_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_16_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_16_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_16_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_16_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_16_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_16_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_16_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_16_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_16_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_16_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_16_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_16_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_16_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_16_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_16_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_16_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_16_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_16_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_16_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_16_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_16_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_16_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_16_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_16_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_16_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_16_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_16_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_16_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_16_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_16_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_16_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_16_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_16_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_16_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_16_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_16_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_16_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_16_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_16_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_16_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_16_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_16_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_16_io_uop_uopc),
    .io_uop_inst                    (_slots_16_io_uop_inst),
    .io_uop_debug_inst              (_slots_16_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_16_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_16_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_16_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_16_io_uop_fu_code),
    .io_uop_iw_state                (_slots_16_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_16_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_16_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_16_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_16_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_16_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_16_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_16_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_16_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_16_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_16_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_16_io_uop_pc_lob),
    .io_uop_taken                   (_slots_16_io_uop_taken),
    .io_uop_imm_packed              (_slots_16_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_16_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_16_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_16_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_16_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_16_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_16_io_uop_pdst),
    .io_uop_prs1                    (_slots_16_io_uop_prs1),
    .io_uop_prs2                    (_slots_16_io_uop_prs2),
    .io_uop_prs3                    (_slots_16_io_uop_prs3),
    .io_uop_ppred                   (_slots_16_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_16_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_16_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_16_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_16_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_16_io_uop_stale_pdst),
    .io_uop_exception               (_slots_16_io_uop_exception),
    .io_uop_exc_cause               (_slots_16_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_16_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_16_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_16_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_16_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_16_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_16_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_16_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_16_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_16_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_16_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_16_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_16_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_16_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_16_io_uop_ldst),
    .io_uop_lrs1                    (_slots_16_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_16_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_16_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_16_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_16_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_16_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_16_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_16_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_16_io_uop_fp_val),
    .io_uop_fp_single               (_slots_16_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_16_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_16_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_16_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_16_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_16_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_16_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_16_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_17 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_17_io_valid),
    .io_will_be_valid               (_slots_17_io_will_be_valid),
    .io_request                     (_slots_17_io_request),
    .io_grant                       (issue_slots_17_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_16),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_17_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_72 ? _slots_21_io_out_uop_uopc : _GEN_71 ? _slots_20_io_out_uop_uopc : _GEN_70 ? _slots_19_io_out_uop_uopc : _slots_18_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_72 ? _slots_21_io_out_uop_inst : _GEN_71 ? _slots_20_io_out_uop_inst : _GEN_70 ? _slots_19_io_out_uop_inst : _slots_18_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_72 ? _slots_21_io_out_uop_debug_inst : _GEN_71 ? _slots_20_io_out_uop_debug_inst : _GEN_70 ? _slots_19_io_out_uop_debug_inst : _slots_18_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_72 ? _slots_21_io_out_uop_is_rvc : _GEN_71 ? _slots_20_io_out_uop_is_rvc : _GEN_70 ? _slots_19_io_out_uop_is_rvc : _slots_18_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_72 ? _slots_21_io_out_uop_debug_pc : _GEN_71 ? _slots_20_io_out_uop_debug_pc : _GEN_70 ? _slots_19_io_out_uop_debug_pc : _slots_18_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_72 ? _slots_21_io_out_uop_iq_type : _GEN_71 ? _slots_20_io_out_uop_iq_type : _GEN_70 ? _slots_19_io_out_uop_iq_type : _slots_18_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_72 ? _slots_21_io_out_uop_fu_code : _GEN_71 ? _slots_20_io_out_uop_fu_code : _GEN_70 ? _slots_19_io_out_uop_fu_code : _slots_18_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_72 ? _slots_21_io_out_uop_iw_state : _GEN_71 ? _slots_20_io_out_uop_iw_state : _GEN_70 ? _slots_19_io_out_uop_iw_state : _slots_18_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_72 ? _slots_21_io_out_uop_iw_p1_poisoned : _GEN_71 ? _slots_20_io_out_uop_iw_p1_poisoned : _GEN_70 ? _slots_19_io_out_uop_iw_p1_poisoned : _slots_18_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_72 ? _slots_21_io_out_uop_iw_p2_poisoned : _GEN_71 ? _slots_20_io_out_uop_iw_p2_poisoned : _GEN_70 ? _slots_19_io_out_uop_iw_p2_poisoned : _slots_18_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_72 ? _slots_21_io_out_uop_is_br : _GEN_71 ? _slots_20_io_out_uop_is_br : _GEN_70 ? _slots_19_io_out_uop_is_br : _slots_18_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_72 ? _slots_21_io_out_uop_is_jalr : _GEN_71 ? _slots_20_io_out_uop_is_jalr : _GEN_70 ? _slots_19_io_out_uop_is_jalr : _slots_18_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_72 ? _slots_21_io_out_uop_is_jal : _GEN_71 ? _slots_20_io_out_uop_is_jal : _GEN_70 ? _slots_19_io_out_uop_is_jal : _slots_18_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_72 ? _slots_21_io_out_uop_is_sfb : _GEN_71 ? _slots_20_io_out_uop_is_sfb : _GEN_70 ? _slots_19_io_out_uop_is_sfb : _slots_18_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_72 ? _slots_21_io_out_uop_br_mask : _GEN_71 ? _slots_20_io_out_uop_br_mask : _GEN_70 ? _slots_19_io_out_uop_br_mask : _slots_18_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_72 ? _slots_21_io_out_uop_br_tag : _GEN_71 ? _slots_20_io_out_uop_br_tag : _GEN_70 ? _slots_19_io_out_uop_br_tag : _slots_18_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_72 ? _slots_21_io_out_uop_ftq_idx : _GEN_71 ? _slots_20_io_out_uop_ftq_idx : _GEN_70 ? _slots_19_io_out_uop_ftq_idx : _slots_18_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_72 ? _slots_21_io_out_uop_edge_inst : _GEN_71 ? _slots_20_io_out_uop_edge_inst : _GEN_70 ? _slots_19_io_out_uop_edge_inst : _slots_18_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_72 ? _slots_21_io_out_uop_pc_lob : _GEN_71 ? _slots_20_io_out_uop_pc_lob : _GEN_70 ? _slots_19_io_out_uop_pc_lob : _slots_18_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_72 ? _slots_21_io_out_uop_taken : _GEN_71 ? _slots_20_io_out_uop_taken : _GEN_70 ? _slots_19_io_out_uop_taken : _slots_18_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_72 ? _slots_21_io_out_uop_imm_packed : _GEN_71 ? _slots_20_io_out_uop_imm_packed : _GEN_70 ? _slots_19_io_out_uop_imm_packed : _slots_18_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_72 ? _slots_21_io_out_uop_csr_addr : _GEN_71 ? _slots_20_io_out_uop_csr_addr : _GEN_70 ? _slots_19_io_out_uop_csr_addr : _slots_18_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_72 ? _slots_21_io_out_uop_rob_idx : _GEN_71 ? _slots_20_io_out_uop_rob_idx : _GEN_70 ? _slots_19_io_out_uop_rob_idx : _slots_18_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_72 ? _slots_21_io_out_uop_ldq_idx : _GEN_71 ? _slots_20_io_out_uop_ldq_idx : _GEN_70 ? _slots_19_io_out_uop_ldq_idx : _slots_18_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_72 ? _slots_21_io_out_uop_stq_idx : _GEN_71 ? _slots_20_io_out_uop_stq_idx : _GEN_70 ? _slots_19_io_out_uop_stq_idx : _slots_18_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_72 ? _slots_21_io_out_uop_rxq_idx : _GEN_71 ? _slots_20_io_out_uop_rxq_idx : _GEN_70 ? _slots_19_io_out_uop_rxq_idx : _slots_18_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_72 ? _slots_21_io_out_uop_pdst : _GEN_71 ? _slots_20_io_out_uop_pdst : _GEN_70 ? _slots_19_io_out_uop_pdst : _slots_18_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_72 ? _slots_21_io_out_uop_prs1 : _GEN_71 ? _slots_20_io_out_uop_prs1 : _GEN_70 ? _slots_19_io_out_uop_prs1 : _slots_18_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_72 ? _slots_21_io_out_uop_prs2 : _GEN_71 ? _slots_20_io_out_uop_prs2 : _GEN_70 ? _slots_19_io_out_uop_prs2 : _slots_18_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_72 ? _slots_21_io_out_uop_prs3 : _GEN_71 ? _slots_20_io_out_uop_prs3 : _GEN_70 ? _slots_19_io_out_uop_prs3 : _slots_18_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_72 ? _slots_21_io_out_uop_ppred : _GEN_71 ? _slots_20_io_out_uop_ppred : _GEN_70 ? _slots_19_io_out_uop_ppred : _slots_18_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_72 ? _slots_21_io_out_uop_prs1_busy : _GEN_71 ? _slots_20_io_out_uop_prs1_busy : _GEN_70 ? _slots_19_io_out_uop_prs1_busy : _slots_18_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_72 ? _slots_21_io_out_uop_prs2_busy : _GEN_71 ? _slots_20_io_out_uop_prs2_busy : _GEN_70 ? _slots_19_io_out_uop_prs2_busy : _slots_18_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_72 ? _slots_21_io_out_uop_prs3_busy : _GEN_71 ? _slots_20_io_out_uop_prs3_busy : _GEN_70 ? _slots_19_io_out_uop_prs3_busy : _slots_18_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_72 ? _slots_21_io_out_uop_ppred_busy : _GEN_71 ? _slots_20_io_out_uop_ppred_busy : _GEN_70 ? _slots_19_io_out_uop_ppred_busy : _slots_18_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_72 ? _slots_21_io_out_uop_stale_pdst : _GEN_71 ? _slots_20_io_out_uop_stale_pdst : _GEN_70 ? _slots_19_io_out_uop_stale_pdst : _slots_18_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_72 ? _slots_21_io_out_uop_exception : _GEN_71 ? _slots_20_io_out_uop_exception : _GEN_70 ? _slots_19_io_out_uop_exception : _slots_18_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_72 ? _slots_21_io_out_uop_exc_cause : _GEN_71 ? _slots_20_io_out_uop_exc_cause : _GEN_70 ? _slots_19_io_out_uop_exc_cause : _slots_18_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_72 ? _slots_21_io_out_uop_bypassable : _GEN_71 ? _slots_20_io_out_uop_bypassable : _GEN_70 ? _slots_19_io_out_uop_bypassable : _slots_18_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_72 ? _slots_21_io_out_uop_mem_cmd : _GEN_71 ? _slots_20_io_out_uop_mem_cmd : _GEN_70 ? _slots_19_io_out_uop_mem_cmd : _slots_18_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_72 ? _slots_21_io_out_uop_mem_size : _GEN_71 ? _slots_20_io_out_uop_mem_size : _GEN_70 ? _slots_19_io_out_uop_mem_size : _slots_18_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_72 ? _slots_21_io_out_uop_mem_signed : _GEN_71 ? _slots_20_io_out_uop_mem_signed : _GEN_70 ? _slots_19_io_out_uop_mem_signed : _slots_18_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_72 ? _slots_21_io_out_uop_is_fence : _GEN_71 ? _slots_20_io_out_uop_is_fence : _GEN_70 ? _slots_19_io_out_uop_is_fence : _slots_18_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_72 ? _slots_21_io_out_uop_is_fencei : _GEN_71 ? _slots_20_io_out_uop_is_fencei : _GEN_70 ? _slots_19_io_out_uop_is_fencei : _slots_18_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_72 ? _slots_21_io_out_uop_is_amo : _GEN_71 ? _slots_20_io_out_uop_is_amo : _GEN_70 ? _slots_19_io_out_uop_is_amo : _slots_18_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_72 ? _slots_21_io_out_uop_uses_ldq : _GEN_71 ? _slots_20_io_out_uop_uses_ldq : _GEN_70 ? _slots_19_io_out_uop_uses_ldq : _slots_18_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_72 ? _slots_21_io_out_uop_uses_stq : _GEN_71 ? _slots_20_io_out_uop_uses_stq : _GEN_70 ? _slots_19_io_out_uop_uses_stq : _slots_18_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_72 ? _slots_21_io_out_uop_is_sys_pc2epc : _GEN_71 ? _slots_20_io_out_uop_is_sys_pc2epc : _GEN_70 ? _slots_19_io_out_uop_is_sys_pc2epc : _slots_18_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_72 ? _slots_21_io_out_uop_is_unique : _GEN_71 ? _slots_20_io_out_uop_is_unique : _GEN_70 ? _slots_19_io_out_uop_is_unique : _slots_18_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_72 ? _slots_21_io_out_uop_flush_on_commit : _GEN_71 ? _slots_20_io_out_uop_flush_on_commit : _GEN_70 ? _slots_19_io_out_uop_flush_on_commit : _slots_18_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_72 ? _slots_21_io_out_uop_ldst_is_rs1 : _GEN_71 ? _slots_20_io_out_uop_ldst_is_rs1 : _GEN_70 ? _slots_19_io_out_uop_ldst_is_rs1 : _slots_18_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_72 ? _slots_21_io_out_uop_ldst : _GEN_71 ? _slots_20_io_out_uop_ldst : _GEN_70 ? _slots_19_io_out_uop_ldst : _slots_18_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_72 ? _slots_21_io_out_uop_lrs1 : _GEN_71 ? _slots_20_io_out_uop_lrs1 : _GEN_70 ? _slots_19_io_out_uop_lrs1 : _slots_18_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_72 ? _slots_21_io_out_uop_lrs2 : _GEN_71 ? _slots_20_io_out_uop_lrs2 : _GEN_70 ? _slots_19_io_out_uop_lrs2 : _slots_18_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_72 ? _slots_21_io_out_uop_lrs3 : _GEN_71 ? _slots_20_io_out_uop_lrs3 : _GEN_70 ? _slots_19_io_out_uop_lrs3 : _slots_18_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_72 ? _slots_21_io_out_uop_ldst_val : _GEN_71 ? _slots_20_io_out_uop_ldst_val : _GEN_70 ? _slots_19_io_out_uop_ldst_val : _slots_18_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_72 ? _slots_21_io_out_uop_dst_rtype : _GEN_71 ? _slots_20_io_out_uop_dst_rtype : _GEN_70 ? _slots_19_io_out_uop_dst_rtype : _slots_18_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_72 ? _slots_21_io_out_uop_lrs1_rtype : _GEN_71 ? _slots_20_io_out_uop_lrs1_rtype : _GEN_70 ? _slots_19_io_out_uop_lrs1_rtype : _slots_18_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_72 ? _slots_21_io_out_uop_lrs2_rtype : _GEN_71 ? _slots_20_io_out_uop_lrs2_rtype : _GEN_70 ? _slots_19_io_out_uop_lrs2_rtype : _slots_18_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_72 ? _slots_21_io_out_uop_frs3_en : _GEN_71 ? _slots_20_io_out_uop_frs3_en : _GEN_70 ? _slots_19_io_out_uop_frs3_en : _slots_18_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_72 ? _slots_21_io_out_uop_fp_val : _GEN_71 ? _slots_20_io_out_uop_fp_val : _GEN_70 ? _slots_19_io_out_uop_fp_val : _slots_18_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_72 ? _slots_21_io_out_uop_fp_single : _GEN_71 ? _slots_20_io_out_uop_fp_single : _GEN_70 ? _slots_19_io_out_uop_fp_single : _slots_18_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_72 ? _slots_21_io_out_uop_xcpt_pf_if : _GEN_71 ? _slots_20_io_out_uop_xcpt_pf_if : _GEN_70 ? _slots_19_io_out_uop_xcpt_pf_if : _slots_18_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_72 ? _slots_21_io_out_uop_xcpt_ae_if : _GEN_71 ? _slots_20_io_out_uop_xcpt_ae_if : _GEN_70 ? _slots_19_io_out_uop_xcpt_ae_if : _slots_18_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_72 ? _slots_21_io_out_uop_xcpt_ma_if : _GEN_71 ? _slots_20_io_out_uop_xcpt_ma_if : _GEN_70 ? _slots_19_io_out_uop_xcpt_ma_if : _slots_18_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_72 ? _slots_21_io_out_uop_bp_debug_if : _GEN_71 ? _slots_20_io_out_uop_bp_debug_if : _GEN_70 ? _slots_19_io_out_uop_bp_debug_if : _slots_18_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_72 ? _slots_21_io_out_uop_bp_xcpt_if : _GEN_71 ? _slots_20_io_out_uop_bp_xcpt_if : _GEN_70 ? _slots_19_io_out_uop_bp_xcpt_if : _slots_18_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_72 ? _slots_21_io_out_uop_debug_fsrc : _GEN_71 ? _slots_20_io_out_uop_debug_fsrc : _GEN_70 ? _slots_19_io_out_uop_debug_fsrc : _slots_18_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_72 ? _slots_21_io_out_uop_debug_tsrc : _GEN_71 ? _slots_20_io_out_uop_debug_tsrc : _GEN_70 ? _slots_19_io_out_uop_debug_tsrc : _slots_18_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_17_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_17_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_17_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_17_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_17_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_17_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_17_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_17_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_17_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_17_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_17_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_17_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_17_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_17_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_17_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_17_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_17_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_17_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_17_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_17_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_17_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_17_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_17_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_17_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_17_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_17_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_17_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_17_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_17_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_17_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_17_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_17_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_17_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_17_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_17_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_17_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_17_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_17_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_17_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_17_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_17_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_17_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_17_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_17_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_17_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_17_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_17_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_17_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_17_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_17_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_17_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_17_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_17_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_17_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_17_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_17_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_17_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_17_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_17_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_17_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_17_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_17_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_17_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_17_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_17_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_17_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_17_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_17_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_17_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_17_io_uop_uopc),
    .io_uop_inst                    (_slots_17_io_uop_inst),
    .io_uop_debug_inst              (_slots_17_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_17_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_17_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_17_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_17_io_uop_fu_code),
    .io_uop_iw_state                (_slots_17_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_17_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_17_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_17_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_17_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_17_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_17_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_17_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_17_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_17_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_17_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_17_io_uop_pc_lob),
    .io_uop_taken                   (_slots_17_io_uop_taken),
    .io_uop_imm_packed              (_slots_17_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_17_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_17_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_17_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_17_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_17_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_17_io_uop_pdst),
    .io_uop_prs1                    (_slots_17_io_uop_prs1),
    .io_uop_prs2                    (_slots_17_io_uop_prs2),
    .io_uop_prs3                    (_slots_17_io_uop_prs3),
    .io_uop_ppred                   (_slots_17_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_17_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_17_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_17_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_17_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_17_io_uop_stale_pdst),
    .io_uop_exception               (_slots_17_io_uop_exception),
    .io_uop_exc_cause               (_slots_17_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_17_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_17_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_17_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_17_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_17_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_17_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_17_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_17_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_17_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_17_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_17_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_17_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_17_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_17_io_uop_ldst),
    .io_uop_lrs1                    (_slots_17_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_17_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_17_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_17_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_17_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_17_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_17_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_17_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_17_io_uop_fp_val),
    .io_uop_fp_single               (_slots_17_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_17_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_17_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_17_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_17_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_17_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_17_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_17_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_18 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_18_io_valid),
    .io_will_be_valid               (_slots_18_io_will_be_valid),
    .io_request                     (_slots_18_io_request),
    .io_grant                       (issue_slots_18_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_17),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_18_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_75 ? _slots_22_io_out_uop_uopc : _GEN_74 ? _slots_21_io_out_uop_uopc : _GEN_73 ? _slots_20_io_out_uop_uopc : _slots_19_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_75 ? _slots_22_io_out_uop_inst : _GEN_74 ? _slots_21_io_out_uop_inst : _GEN_73 ? _slots_20_io_out_uop_inst : _slots_19_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_75 ? _slots_22_io_out_uop_debug_inst : _GEN_74 ? _slots_21_io_out_uop_debug_inst : _GEN_73 ? _slots_20_io_out_uop_debug_inst : _slots_19_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_75 ? _slots_22_io_out_uop_is_rvc : _GEN_74 ? _slots_21_io_out_uop_is_rvc : _GEN_73 ? _slots_20_io_out_uop_is_rvc : _slots_19_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_75 ? _slots_22_io_out_uop_debug_pc : _GEN_74 ? _slots_21_io_out_uop_debug_pc : _GEN_73 ? _slots_20_io_out_uop_debug_pc : _slots_19_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_75 ? _slots_22_io_out_uop_iq_type : _GEN_74 ? _slots_21_io_out_uop_iq_type : _GEN_73 ? _slots_20_io_out_uop_iq_type : _slots_19_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_75 ? _slots_22_io_out_uop_fu_code : _GEN_74 ? _slots_21_io_out_uop_fu_code : _GEN_73 ? _slots_20_io_out_uop_fu_code : _slots_19_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_75 ? _slots_22_io_out_uop_iw_state : _GEN_74 ? _slots_21_io_out_uop_iw_state : _GEN_73 ? _slots_20_io_out_uop_iw_state : _slots_19_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_75 ? _slots_22_io_out_uop_iw_p1_poisoned : _GEN_74 ? _slots_21_io_out_uop_iw_p1_poisoned : _GEN_73 ? _slots_20_io_out_uop_iw_p1_poisoned : _slots_19_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_75 ? _slots_22_io_out_uop_iw_p2_poisoned : _GEN_74 ? _slots_21_io_out_uop_iw_p2_poisoned : _GEN_73 ? _slots_20_io_out_uop_iw_p2_poisoned : _slots_19_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_75 ? _slots_22_io_out_uop_is_br : _GEN_74 ? _slots_21_io_out_uop_is_br : _GEN_73 ? _slots_20_io_out_uop_is_br : _slots_19_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_75 ? _slots_22_io_out_uop_is_jalr : _GEN_74 ? _slots_21_io_out_uop_is_jalr : _GEN_73 ? _slots_20_io_out_uop_is_jalr : _slots_19_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_75 ? _slots_22_io_out_uop_is_jal : _GEN_74 ? _slots_21_io_out_uop_is_jal : _GEN_73 ? _slots_20_io_out_uop_is_jal : _slots_19_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_75 ? _slots_22_io_out_uop_is_sfb : _GEN_74 ? _slots_21_io_out_uop_is_sfb : _GEN_73 ? _slots_20_io_out_uop_is_sfb : _slots_19_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_75 ? _slots_22_io_out_uop_br_mask : _GEN_74 ? _slots_21_io_out_uop_br_mask : _GEN_73 ? _slots_20_io_out_uop_br_mask : _slots_19_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_75 ? _slots_22_io_out_uop_br_tag : _GEN_74 ? _slots_21_io_out_uop_br_tag : _GEN_73 ? _slots_20_io_out_uop_br_tag : _slots_19_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_75 ? _slots_22_io_out_uop_ftq_idx : _GEN_74 ? _slots_21_io_out_uop_ftq_idx : _GEN_73 ? _slots_20_io_out_uop_ftq_idx : _slots_19_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_75 ? _slots_22_io_out_uop_edge_inst : _GEN_74 ? _slots_21_io_out_uop_edge_inst : _GEN_73 ? _slots_20_io_out_uop_edge_inst : _slots_19_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_75 ? _slots_22_io_out_uop_pc_lob : _GEN_74 ? _slots_21_io_out_uop_pc_lob : _GEN_73 ? _slots_20_io_out_uop_pc_lob : _slots_19_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_75 ? _slots_22_io_out_uop_taken : _GEN_74 ? _slots_21_io_out_uop_taken : _GEN_73 ? _slots_20_io_out_uop_taken : _slots_19_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_75 ? _slots_22_io_out_uop_imm_packed : _GEN_74 ? _slots_21_io_out_uop_imm_packed : _GEN_73 ? _slots_20_io_out_uop_imm_packed : _slots_19_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_75 ? _slots_22_io_out_uop_csr_addr : _GEN_74 ? _slots_21_io_out_uop_csr_addr : _GEN_73 ? _slots_20_io_out_uop_csr_addr : _slots_19_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_75 ? _slots_22_io_out_uop_rob_idx : _GEN_74 ? _slots_21_io_out_uop_rob_idx : _GEN_73 ? _slots_20_io_out_uop_rob_idx : _slots_19_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_75 ? _slots_22_io_out_uop_ldq_idx : _GEN_74 ? _slots_21_io_out_uop_ldq_idx : _GEN_73 ? _slots_20_io_out_uop_ldq_idx : _slots_19_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_75 ? _slots_22_io_out_uop_stq_idx : _GEN_74 ? _slots_21_io_out_uop_stq_idx : _GEN_73 ? _slots_20_io_out_uop_stq_idx : _slots_19_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_75 ? _slots_22_io_out_uop_rxq_idx : _GEN_74 ? _slots_21_io_out_uop_rxq_idx : _GEN_73 ? _slots_20_io_out_uop_rxq_idx : _slots_19_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_75 ? _slots_22_io_out_uop_pdst : _GEN_74 ? _slots_21_io_out_uop_pdst : _GEN_73 ? _slots_20_io_out_uop_pdst : _slots_19_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_75 ? _slots_22_io_out_uop_prs1 : _GEN_74 ? _slots_21_io_out_uop_prs1 : _GEN_73 ? _slots_20_io_out_uop_prs1 : _slots_19_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_75 ? _slots_22_io_out_uop_prs2 : _GEN_74 ? _slots_21_io_out_uop_prs2 : _GEN_73 ? _slots_20_io_out_uop_prs2 : _slots_19_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_75 ? _slots_22_io_out_uop_prs3 : _GEN_74 ? _slots_21_io_out_uop_prs3 : _GEN_73 ? _slots_20_io_out_uop_prs3 : _slots_19_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_75 ? _slots_22_io_out_uop_ppred : _GEN_74 ? _slots_21_io_out_uop_ppred : _GEN_73 ? _slots_20_io_out_uop_ppred : _slots_19_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_75 ? _slots_22_io_out_uop_prs1_busy : _GEN_74 ? _slots_21_io_out_uop_prs1_busy : _GEN_73 ? _slots_20_io_out_uop_prs1_busy : _slots_19_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_75 ? _slots_22_io_out_uop_prs2_busy : _GEN_74 ? _slots_21_io_out_uop_prs2_busy : _GEN_73 ? _slots_20_io_out_uop_prs2_busy : _slots_19_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_75 ? _slots_22_io_out_uop_prs3_busy : _GEN_74 ? _slots_21_io_out_uop_prs3_busy : _GEN_73 ? _slots_20_io_out_uop_prs3_busy : _slots_19_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_75 ? _slots_22_io_out_uop_ppred_busy : _GEN_74 ? _slots_21_io_out_uop_ppred_busy : _GEN_73 ? _slots_20_io_out_uop_ppred_busy : _slots_19_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_75 ? _slots_22_io_out_uop_stale_pdst : _GEN_74 ? _slots_21_io_out_uop_stale_pdst : _GEN_73 ? _slots_20_io_out_uop_stale_pdst : _slots_19_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_75 ? _slots_22_io_out_uop_exception : _GEN_74 ? _slots_21_io_out_uop_exception : _GEN_73 ? _slots_20_io_out_uop_exception : _slots_19_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_75 ? _slots_22_io_out_uop_exc_cause : _GEN_74 ? _slots_21_io_out_uop_exc_cause : _GEN_73 ? _slots_20_io_out_uop_exc_cause : _slots_19_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_75 ? _slots_22_io_out_uop_bypassable : _GEN_74 ? _slots_21_io_out_uop_bypassable : _GEN_73 ? _slots_20_io_out_uop_bypassable : _slots_19_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_75 ? _slots_22_io_out_uop_mem_cmd : _GEN_74 ? _slots_21_io_out_uop_mem_cmd : _GEN_73 ? _slots_20_io_out_uop_mem_cmd : _slots_19_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_75 ? _slots_22_io_out_uop_mem_size : _GEN_74 ? _slots_21_io_out_uop_mem_size : _GEN_73 ? _slots_20_io_out_uop_mem_size : _slots_19_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_75 ? _slots_22_io_out_uop_mem_signed : _GEN_74 ? _slots_21_io_out_uop_mem_signed : _GEN_73 ? _slots_20_io_out_uop_mem_signed : _slots_19_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_75 ? _slots_22_io_out_uop_is_fence : _GEN_74 ? _slots_21_io_out_uop_is_fence : _GEN_73 ? _slots_20_io_out_uop_is_fence : _slots_19_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_75 ? _slots_22_io_out_uop_is_fencei : _GEN_74 ? _slots_21_io_out_uop_is_fencei : _GEN_73 ? _slots_20_io_out_uop_is_fencei : _slots_19_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_75 ? _slots_22_io_out_uop_is_amo : _GEN_74 ? _slots_21_io_out_uop_is_amo : _GEN_73 ? _slots_20_io_out_uop_is_amo : _slots_19_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_75 ? _slots_22_io_out_uop_uses_ldq : _GEN_74 ? _slots_21_io_out_uop_uses_ldq : _GEN_73 ? _slots_20_io_out_uop_uses_ldq : _slots_19_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_75 ? _slots_22_io_out_uop_uses_stq : _GEN_74 ? _slots_21_io_out_uop_uses_stq : _GEN_73 ? _slots_20_io_out_uop_uses_stq : _slots_19_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_75 ? _slots_22_io_out_uop_is_sys_pc2epc : _GEN_74 ? _slots_21_io_out_uop_is_sys_pc2epc : _GEN_73 ? _slots_20_io_out_uop_is_sys_pc2epc : _slots_19_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_75 ? _slots_22_io_out_uop_is_unique : _GEN_74 ? _slots_21_io_out_uop_is_unique : _GEN_73 ? _slots_20_io_out_uop_is_unique : _slots_19_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_75 ? _slots_22_io_out_uop_flush_on_commit : _GEN_74 ? _slots_21_io_out_uop_flush_on_commit : _GEN_73 ? _slots_20_io_out_uop_flush_on_commit : _slots_19_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_75 ? _slots_22_io_out_uop_ldst_is_rs1 : _GEN_74 ? _slots_21_io_out_uop_ldst_is_rs1 : _GEN_73 ? _slots_20_io_out_uop_ldst_is_rs1 : _slots_19_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_75 ? _slots_22_io_out_uop_ldst : _GEN_74 ? _slots_21_io_out_uop_ldst : _GEN_73 ? _slots_20_io_out_uop_ldst : _slots_19_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_75 ? _slots_22_io_out_uop_lrs1 : _GEN_74 ? _slots_21_io_out_uop_lrs1 : _GEN_73 ? _slots_20_io_out_uop_lrs1 : _slots_19_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_75 ? _slots_22_io_out_uop_lrs2 : _GEN_74 ? _slots_21_io_out_uop_lrs2 : _GEN_73 ? _slots_20_io_out_uop_lrs2 : _slots_19_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_75 ? _slots_22_io_out_uop_lrs3 : _GEN_74 ? _slots_21_io_out_uop_lrs3 : _GEN_73 ? _slots_20_io_out_uop_lrs3 : _slots_19_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_75 ? _slots_22_io_out_uop_ldst_val : _GEN_74 ? _slots_21_io_out_uop_ldst_val : _GEN_73 ? _slots_20_io_out_uop_ldst_val : _slots_19_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_75 ? _slots_22_io_out_uop_dst_rtype : _GEN_74 ? _slots_21_io_out_uop_dst_rtype : _GEN_73 ? _slots_20_io_out_uop_dst_rtype : _slots_19_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_75 ? _slots_22_io_out_uop_lrs1_rtype : _GEN_74 ? _slots_21_io_out_uop_lrs1_rtype : _GEN_73 ? _slots_20_io_out_uop_lrs1_rtype : _slots_19_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_75 ? _slots_22_io_out_uop_lrs2_rtype : _GEN_74 ? _slots_21_io_out_uop_lrs2_rtype : _GEN_73 ? _slots_20_io_out_uop_lrs2_rtype : _slots_19_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_75 ? _slots_22_io_out_uop_frs3_en : _GEN_74 ? _slots_21_io_out_uop_frs3_en : _GEN_73 ? _slots_20_io_out_uop_frs3_en : _slots_19_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_75 ? _slots_22_io_out_uop_fp_val : _GEN_74 ? _slots_21_io_out_uop_fp_val : _GEN_73 ? _slots_20_io_out_uop_fp_val : _slots_19_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_75 ? _slots_22_io_out_uop_fp_single : _GEN_74 ? _slots_21_io_out_uop_fp_single : _GEN_73 ? _slots_20_io_out_uop_fp_single : _slots_19_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_75 ? _slots_22_io_out_uop_xcpt_pf_if : _GEN_74 ? _slots_21_io_out_uop_xcpt_pf_if : _GEN_73 ? _slots_20_io_out_uop_xcpt_pf_if : _slots_19_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_75 ? _slots_22_io_out_uop_xcpt_ae_if : _GEN_74 ? _slots_21_io_out_uop_xcpt_ae_if : _GEN_73 ? _slots_20_io_out_uop_xcpt_ae_if : _slots_19_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_75 ? _slots_22_io_out_uop_xcpt_ma_if : _GEN_74 ? _slots_21_io_out_uop_xcpt_ma_if : _GEN_73 ? _slots_20_io_out_uop_xcpt_ma_if : _slots_19_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_75 ? _slots_22_io_out_uop_bp_debug_if : _GEN_74 ? _slots_21_io_out_uop_bp_debug_if : _GEN_73 ? _slots_20_io_out_uop_bp_debug_if : _slots_19_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_75 ? _slots_22_io_out_uop_bp_xcpt_if : _GEN_74 ? _slots_21_io_out_uop_bp_xcpt_if : _GEN_73 ? _slots_20_io_out_uop_bp_xcpt_if : _slots_19_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_75 ? _slots_22_io_out_uop_debug_fsrc : _GEN_74 ? _slots_21_io_out_uop_debug_fsrc : _GEN_73 ? _slots_20_io_out_uop_debug_fsrc : _slots_19_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_75 ? _slots_22_io_out_uop_debug_tsrc : _GEN_74 ? _slots_21_io_out_uop_debug_tsrc : _GEN_73 ? _slots_20_io_out_uop_debug_tsrc : _slots_19_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_18_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_18_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_18_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_18_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_18_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_18_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_18_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_18_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_18_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_18_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_18_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_18_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_18_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_18_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_18_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_18_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_18_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_18_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_18_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_18_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_18_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_18_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_18_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_18_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_18_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_18_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_18_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_18_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_18_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_18_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_18_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_18_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_18_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_18_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_18_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_18_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_18_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_18_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_18_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_18_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_18_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_18_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_18_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_18_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_18_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_18_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_18_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_18_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_18_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_18_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_18_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_18_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_18_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_18_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_18_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_18_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_18_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_18_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_18_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_18_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_18_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_18_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_18_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_18_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_18_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_18_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_18_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_18_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_18_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_18_io_uop_uopc),
    .io_uop_inst                    (_slots_18_io_uop_inst),
    .io_uop_debug_inst              (_slots_18_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_18_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_18_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_18_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_18_io_uop_fu_code),
    .io_uop_iw_state                (_slots_18_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_18_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_18_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_18_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_18_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_18_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_18_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_18_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_18_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_18_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_18_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_18_io_uop_pc_lob),
    .io_uop_taken                   (_slots_18_io_uop_taken),
    .io_uop_imm_packed              (_slots_18_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_18_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_18_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_18_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_18_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_18_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_18_io_uop_pdst),
    .io_uop_prs1                    (_slots_18_io_uop_prs1),
    .io_uop_prs2                    (_slots_18_io_uop_prs2),
    .io_uop_prs3                    (_slots_18_io_uop_prs3),
    .io_uop_ppred                   (_slots_18_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_18_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_18_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_18_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_18_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_18_io_uop_stale_pdst),
    .io_uop_exception               (_slots_18_io_uop_exception),
    .io_uop_exc_cause               (_slots_18_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_18_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_18_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_18_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_18_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_18_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_18_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_18_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_18_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_18_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_18_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_18_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_18_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_18_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_18_io_uop_ldst),
    .io_uop_lrs1                    (_slots_18_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_18_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_18_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_18_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_18_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_18_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_18_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_18_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_18_io_uop_fp_val),
    .io_uop_fp_single               (_slots_18_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_18_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_18_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_18_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_18_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_18_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_18_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_18_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_19 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_19_io_valid),
    .io_will_be_valid               (_slots_19_io_will_be_valid),
    .io_request                     (_slots_19_io_request),
    .io_grant                       (issue_slots_19_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_18),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_19_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_78 ? _slots_23_io_out_uop_uopc : _GEN_77 ? _slots_22_io_out_uop_uopc : _GEN_76 ? _slots_21_io_out_uop_uopc : _slots_20_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_78 ? _slots_23_io_out_uop_inst : _GEN_77 ? _slots_22_io_out_uop_inst : _GEN_76 ? _slots_21_io_out_uop_inst : _slots_20_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_78 ? _slots_23_io_out_uop_debug_inst : _GEN_77 ? _slots_22_io_out_uop_debug_inst : _GEN_76 ? _slots_21_io_out_uop_debug_inst : _slots_20_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_78 ? _slots_23_io_out_uop_is_rvc : _GEN_77 ? _slots_22_io_out_uop_is_rvc : _GEN_76 ? _slots_21_io_out_uop_is_rvc : _slots_20_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_78 ? _slots_23_io_out_uop_debug_pc : _GEN_77 ? _slots_22_io_out_uop_debug_pc : _GEN_76 ? _slots_21_io_out_uop_debug_pc : _slots_20_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_78 ? _slots_23_io_out_uop_iq_type : _GEN_77 ? _slots_22_io_out_uop_iq_type : _GEN_76 ? _slots_21_io_out_uop_iq_type : _slots_20_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_78 ? _slots_23_io_out_uop_fu_code : _GEN_77 ? _slots_22_io_out_uop_fu_code : _GEN_76 ? _slots_21_io_out_uop_fu_code : _slots_20_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_78 ? _slots_23_io_out_uop_iw_state : _GEN_77 ? _slots_22_io_out_uop_iw_state : _GEN_76 ? _slots_21_io_out_uop_iw_state : _slots_20_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_78 ? _slots_23_io_out_uop_iw_p1_poisoned : _GEN_77 ? _slots_22_io_out_uop_iw_p1_poisoned : _GEN_76 ? _slots_21_io_out_uop_iw_p1_poisoned : _slots_20_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_78 ? _slots_23_io_out_uop_iw_p2_poisoned : _GEN_77 ? _slots_22_io_out_uop_iw_p2_poisoned : _GEN_76 ? _slots_21_io_out_uop_iw_p2_poisoned : _slots_20_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_78 ? _slots_23_io_out_uop_is_br : _GEN_77 ? _slots_22_io_out_uop_is_br : _GEN_76 ? _slots_21_io_out_uop_is_br : _slots_20_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_78 ? _slots_23_io_out_uop_is_jalr : _GEN_77 ? _slots_22_io_out_uop_is_jalr : _GEN_76 ? _slots_21_io_out_uop_is_jalr : _slots_20_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_78 ? _slots_23_io_out_uop_is_jal : _GEN_77 ? _slots_22_io_out_uop_is_jal : _GEN_76 ? _slots_21_io_out_uop_is_jal : _slots_20_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_78 ? _slots_23_io_out_uop_is_sfb : _GEN_77 ? _slots_22_io_out_uop_is_sfb : _GEN_76 ? _slots_21_io_out_uop_is_sfb : _slots_20_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_78 ? _slots_23_io_out_uop_br_mask : _GEN_77 ? _slots_22_io_out_uop_br_mask : _GEN_76 ? _slots_21_io_out_uop_br_mask : _slots_20_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_78 ? _slots_23_io_out_uop_br_tag : _GEN_77 ? _slots_22_io_out_uop_br_tag : _GEN_76 ? _slots_21_io_out_uop_br_tag : _slots_20_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_78 ? _slots_23_io_out_uop_ftq_idx : _GEN_77 ? _slots_22_io_out_uop_ftq_idx : _GEN_76 ? _slots_21_io_out_uop_ftq_idx : _slots_20_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_78 ? _slots_23_io_out_uop_edge_inst : _GEN_77 ? _slots_22_io_out_uop_edge_inst : _GEN_76 ? _slots_21_io_out_uop_edge_inst : _slots_20_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_78 ? _slots_23_io_out_uop_pc_lob : _GEN_77 ? _slots_22_io_out_uop_pc_lob : _GEN_76 ? _slots_21_io_out_uop_pc_lob : _slots_20_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_78 ? _slots_23_io_out_uop_taken : _GEN_77 ? _slots_22_io_out_uop_taken : _GEN_76 ? _slots_21_io_out_uop_taken : _slots_20_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_78 ? _slots_23_io_out_uop_imm_packed : _GEN_77 ? _slots_22_io_out_uop_imm_packed : _GEN_76 ? _slots_21_io_out_uop_imm_packed : _slots_20_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_78 ? _slots_23_io_out_uop_csr_addr : _GEN_77 ? _slots_22_io_out_uop_csr_addr : _GEN_76 ? _slots_21_io_out_uop_csr_addr : _slots_20_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_78 ? _slots_23_io_out_uop_rob_idx : _GEN_77 ? _slots_22_io_out_uop_rob_idx : _GEN_76 ? _slots_21_io_out_uop_rob_idx : _slots_20_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_78 ? _slots_23_io_out_uop_ldq_idx : _GEN_77 ? _slots_22_io_out_uop_ldq_idx : _GEN_76 ? _slots_21_io_out_uop_ldq_idx : _slots_20_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_78 ? _slots_23_io_out_uop_stq_idx : _GEN_77 ? _slots_22_io_out_uop_stq_idx : _GEN_76 ? _slots_21_io_out_uop_stq_idx : _slots_20_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_78 ? _slots_23_io_out_uop_rxq_idx : _GEN_77 ? _slots_22_io_out_uop_rxq_idx : _GEN_76 ? _slots_21_io_out_uop_rxq_idx : _slots_20_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_78 ? _slots_23_io_out_uop_pdst : _GEN_77 ? _slots_22_io_out_uop_pdst : _GEN_76 ? _slots_21_io_out_uop_pdst : _slots_20_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_78 ? _slots_23_io_out_uop_prs1 : _GEN_77 ? _slots_22_io_out_uop_prs1 : _GEN_76 ? _slots_21_io_out_uop_prs1 : _slots_20_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_78 ? _slots_23_io_out_uop_prs2 : _GEN_77 ? _slots_22_io_out_uop_prs2 : _GEN_76 ? _slots_21_io_out_uop_prs2 : _slots_20_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_78 ? _slots_23_io_out_uop_prs3 : _GEN_77 ? _slots_22_io_out_uop_prs3 : _GEN_76 ? _slots_21_io_out_uop_prs3 : _slots_20_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_78 ? _slots_23_io_out_uop_ppred : _GEN_77 ? _slots_22_io_out_uop_ppred : _GEN_76 ? _slots_21_io_out_uop_ppred : _slots_20_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_78 ? _slots_23_io_out_uop_prs1_busy : _GEN_77 ? _slots_22_io_out_uop_prs1_busy : _GEN_76 ? _slots_21_io_out_uop_prs1_busy : _slots_20_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_78 ? _slots_23_io_out_uop_prs2_busy : _GEN_77 ? _slots_22_io_out_uop_prs2_busy : _GEN_76 ? _slots_21_io_out_uop_prs2_busy : _slots_20_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_78 ? _slots_23_io_out_uop_prs3_busy : _GEN_77 ? _slots_22_io_out_uop_prs3_busy : _GEN_76 ? _slots_21_io_out_uop_prs3_busy : _slots_20_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_78 ? _slots_23_io_out_uop_ppred_busy : _GEN_77 ? _slots_22_io_out_uop_ppred_busy : _GEN_76 ? _slots_21_io_out_uop_ppred_busy : _slots_20_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_78 ? _slots_23_io_out_uop_stale_pdst : _GEN_77 ? _slots_22_io_out_uop_stale_pdst : _GEN_76 ? _slots_21_io_out_uop_stale_pdst : _slots_20_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_78 ? _slots_23_io_out_uop_exception : _GEN_77 ? _slots_22_io_out_uop_exception : _GEN_76 ? _slots_21_io_out_uop_exception : _slots_20_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_78 ? _slots_23_io_out_uop_exc_cause : _GEN_77 ? _slots_22_io_out_uop_exc_cause : _GEN_76 ? _slots_21_io_out_uop_exc_cause : _slots_20_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_78 ? _slots_23_io_out_uop_bypassable : _GEN_77 ? _slots_22_io_out_uop_bypassable : _GEN_76 ? _slots_21_io_out_uop_bypassable : _slots_20_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_78 ? _slots_23_io_out_uop_mem_cmd : _GEN_77 ? _slots_22_io_out_uop_mem_cmd : _GEN_76 ? _slots_21_io_out_uop_mem_cmd : _slots_20_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_78 ? _slots_23_io_out_uop_mem_size : _GEN_77 ? _slots_22_io_out_uop_mem_size : _GEN_76 ? _slots_21_io_out_uop_mem_size : _slots_20_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_78 ? _slots_23_io_out_uop_mem_signed : _GEN_77 ? _slots_22_io_out_uop_mem_signed : _GEN_76 ? _slots_21_io_out_uop_mem_signed : _slots_20_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_78 ? _slots_23_io_out_uop_is_fence : _GEN_77 ? _slots_22_io_out_uop_is_fence : _GEN_76 ? _slots_21_io_out_uop_is_fence : _slots_20_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_78 ? _slots_23_io_out_uop_is_fencei : _GEN_77 ? _slots_22_io_out_uop_is_fencei : _GEN_76 ? _slots_21_io_out_uop_is_fencei : _slots_20_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_78 ? _slots_23_io_out_uop_is_amo : _GEN_77 ? _slots_22_io_out_uop_is_amo : _GEN_76 ? _slots_21_io_out_uop_is_amo : _slots_20_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_78 ? _slots_23_io_out_uop_uses_ldq : _GEN_77 ? _slots_22_io_out_uop_uses_ldq : _GEN_76 ? _slots_21_io_out_uop_uses_ldq : _slots_20_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_78 ? _slots_23_io_out_uop_uses_stq : _GEN_77 ? _slots_22_io_out_uop_uses_stq : _GEN_76 ? _slots_21_io_out_uop_uses_stq : _slots_20_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_78 ? _slots_23_io_out_uop_is_sys_pc2epc : _GEN_77 ? _slots_22_io_out_uop_is_sys_pc2epc : _GEN_76 ? _slots_21_io_out_uop_is_sys_pc2epc : _slots_20_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_78 ? _slots_23_io_out_uop_is_unique : _GEN_77 ? _slots_22_io_out_uop_is_unique : _GEN_76 ? _slots_21_io_out_uop_is_unique : _slots_20_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_78 ? _slots_23_io_out_uop_flush_on_commit : _GEN_77 ? _slots_22_io_out_uop_flush_on_commit : _GEN_76 ? _slots_21_io_out_uop_flush_on_commit : _slots_20_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_78 ? _slots_23_io_out_uop_ldst_is_rs1 : _GEN_77 ? _slots_22_io_out_uop_ldst_is_rs1 : _GEN_76 ? _slots_21_io_out_uop_ldst_is_rs1 : _slots_20_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_78 ? _slots_23_io_out_uop_ldst : _GEN_77 ? _slots_22_io_out_uop_ldst : _GEN_76 ? _slots_21_io_out_uop_ldst : _slots_20_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_78 ? _slots_23_io_out_uop_lrs1 : _GEN_77 ? _slots_22_io_out_uop_lrs1 : _GEN_76 ? _slots_21_io_out_uop_lrs1 : _slots_20_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_78 ? _slots_23_io_out_uop_lrs2 : _GEN_77 ? _slots_22_io_out_uop_lrs2 : _GEN_76 ? _slots_21_io_out_uop_lrs2 : _slots_20_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_78 ? _slots_23_io_out_uop_lrs3 : _GEN_77 ? _slots_22_io_out_uop_lrs3 : _GEN_76 ? _slots_21_io_out_uop_lrs3 : _slots_20_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_78 ? _slots_23_io_out_uop_ldst_val : _GEN_77 ? _slots_22_io_out_uop_ldst_val : _GEN_76 ? _slots_21_io_out_uop_ldst_val : _slots_20_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_78 ? _slots_23_io_out_uop_dst_rtype : _GEN_77 ? _slots_22_io_out_uop_dst_rtype : _GEN_76 ? _slots_21_io_out_uop_dst_rtype : _slots_20_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_78 ? _slots_23_io_out_uop_lrs1_rtype : _GEN_77 ? _slots_22_io_out_uop_lrs1_rtype : _GEN_76 ? _slots_21_io_out_uop_lrs1_rtype : _slots_20_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_78 ? _slots_23_io_out_uop_lrs2_rtype : _GEN_77 ? _slots_22_io_out_uop_lrs2_rtype : _GEN_76 ? _slots_21_io_out_uop_lrs2_rtype : _slots_20_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_78 ? _slots_23_io_out_uop_frs3_en : _GEN_77 ? _slots_22_io_out_uop_frs3_en : _GEN_76 ? _slots_21_io_out_uop_frs3_en : _slots_20_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_78 ? _slots_23_io_out_uop_fp_val : _GEN_77 ? _slots_22_io_out_uop_fp_val : _GEN_76 ? _slots_21_io_out_uop_fp_val : _slots_20_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_78 ? _slots_23_io_out_uop_fp_single : _GEN_77 ? _slots_22_io_out_uop_fp_single : _GEN_76 ? _slots_21_io_out_uop_fp_single : _slots_20_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_78 ? _slots_23_io_out_uop_xcpt_pf_if : _GEN_77 ? _slots_22_io_out_uop_xcpt_pf_if : _GEN_76 ? _slots_21_io_out_uop_xcpt_pf_if : _slots_20_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_78 ? _slots_23_io_out_uop_xcpt_ae_if : _GEN_77 ? _slots_22_io_out_uop_xcpt_ae_if : _GEN_76 ? _slots_21_io_out_uop_xcpt_ae_if : _slots_20_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_78 ? _slots_23_io_out_uop_xcpt_ma_if : _GEN_77 ? _slots_22_io_out_uop_xcpt_ma_if : _GEN_76 ? _slots_21_io_out_uop_xcpt_ma_if : _slots_20_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_78 ? _slots_23_io_out_uop_bp_debug_if : _GEN_77 ? _slots_22_io_out_uop_bp_debug_if : _GEN_76 ? _slots_21_io_out_uop_bp_debug_if : _slots_20_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_78 ? _slots_23_io_out_uop_bp_xcpt_if : _GEN_77 ? _slots_22_io_out_uop_bp_xcpt_if : _GEN_76 ? _slots_21_io_out_uop_bp_xcpt_if : _slots_20_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_78 ? _slots_23_io_out_uop_debug_fsrc : _GEN_77 ? _slots_22_io_out_uop_debug_fsrc : _GEN_76 ? _slots_21_io_out_uop_debug_fsrc : _slots_20_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_78 ? _slots_23_io_out_uop_debug_tsrc : _GEN_77 ? _slots_22_io_out_uop_debug_tsrc : _GEN_76 ? _slots_21_io_out_uop_debug_tsrc : _slots_20_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_19_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_19_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_19_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_19_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_19_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_19_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_19_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_19_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_19_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_19_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_19_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_19_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_19_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_19_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_19_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_19_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_19_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_19_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_19_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_19_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_19_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_19_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_19_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_19_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_19_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_19_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_19_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_19_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_19_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_19_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_19_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_19_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_19_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_19_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_19_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_19_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_19_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_19_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_19_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_19_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_19_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_19_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_19_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_19_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_19_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_19_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_19_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_19_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_19_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_19_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_19_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_19_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_19_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_19_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_19_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_19_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_19_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_19_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_19_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_19_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_19_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_19_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_19_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_19_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_19_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_19_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_19_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_19_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_19_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_19_io_uop_uopc),
    .io_uop_inst                    (_slots_19_io_uop_inst),
    .io_uop_debug_inst              (_slots_19_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_19_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_19_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_19_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_19_io_uop_fu_code),
    .io_uop_iw_state                (_slots_19_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_19_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_19_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_19_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_19_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_19_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_19_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_19_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_19_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_19_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_19_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_19_io_uop_pc_lob),
    .io_uop_taken                   (_slots_19_io_uop_taken),
    .io_uop_imm_packed              (_slots_19_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_19_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_19_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_19_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_19_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_19_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_19_io_uop_pdst),
    .io_uop_prs1                    (_slots_19_io_uop_prs1),
    .io_uop_prs2                    (_slots_19_io_uop_prs2),
    .io_uop_prs3                    (_slots_19_io_uop_prs3),
    .io_uop_ppred                   (_slots_19_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_19_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_19_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_19_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_19_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_19_io_uop_stale_pdst),
    .io_uop_exception               (_slots_19_io_uop_exception),
    .io_uop_exc_cause               (_slots_19_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_19_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_19_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_19_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_19_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_19_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_19_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_19_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_19_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_19_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_19_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_19_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_19_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_19_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_19_io_uop_ldst),
    .io_uop_lrs1                    (_slots_19_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_19_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_19_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_19_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_19_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_19_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_19_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_19_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_19_io_uop_fp_val),
    .io_uop_fp_single               (_slots_19_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_19_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_19_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_19_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_19_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_19_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_19_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_19_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_20 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_20_io_valid),
    .io_will_be_valid               (_slots_20_io_will_be_valid),
    .io_request                     (_slots_20_io_request),
    .io_grant                       (issue_slots_20_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_19),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_20_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_81 ? io_dis_uops_0_bits_uopc : _GEN_80 ? _slots_23_io_out_uop_uopc : _GEN_79 ? _slots_22_io_out_uop_uopc : _slots_21_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_81 ? io_dis_uops_0_bits_inst : _GEN_80 ? _slots_23_io_out_uop_inst : _GEN_79 ? _slots_22_io_out_uop_inst : _slots_21_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_81 ? io_dis_uops_0_bits_debug_inst : _GEN_80 ? _slots_23_io_out_uop_debug_inst : _GEN_79 ? _slots_22_io_out_uop_debug_inst : _slots_21_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_81 ? io_dis_uops_0_bits_is_rvc : _GEN_80 ? _slots_23_io_out_uop_is_rvc : _GEN_79 ? _slots_22_io_out_uop_is_rvc : _slots_21_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_81 ? io_dis_uops_0_bits_debug_pc : _GEN_80 ? _slots_23_io_out_uop_debug_pc : _GEN_79 ? _slots_22_io_out_uop_debug_pc : _slots_21_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_81 ? io_dis_uops_0_bits_iq_type : _GEN_80 ? _slots_23_io_out_uop_iq_type : _GEN_79 ? _slots_22_io_out_uop_iq_type : _slots_21_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_81 ? io_dis_uops_0_bits_fu_code : _GEN_80 ? _slots_23_io_out_uop_fu_code : _GEN_79 ? _slots_22_io_out_uop_fu_code : _slots_21_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_81 ? _GEN_1 : _GEN_80 ? _slots_23_io_out_uop_iw_state : _GEN_79 ? _slots_22_io_out_uop_iw_state : _slots_21_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_81 & (_GEN_80 ? _slots_23_io_out_uop_iw_p1_poisoned : _GEN_79 ? _slots_22_io_out_uop_iw_p1_poisoned : _slots_21_io_out_uop_iw_p1_poisoned)),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_81 & (_GEN_80 ? _slots_23_io_out_uop_iw_p2_poisoned : _GEN_79 ? _slots_22_io_out_uop_iw_p2_poisoned : _slots_21_io_out_uop_iw_p2_poisoned)),
    .io_in_uop_bits_is_br           (_GEN_81 ? io_dis_uops_0_bits_is_br : _GEN_80 ? _slots_23_io_out_uop_is_br : _GEN_79 ? _slots_22_io_out_uop_is_br : _slots_21_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_81 ? io_dis_uops_0_bits_is_jalr : _GEN_80 ? _slots_23_io_out_uop_is_jalr : _GEN_79 ? _slots_22_io_out_uop_is_jalr : _slots_21_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_81 ? io_dis_uops_0_bits_is_jal : _GEN_80 ? _slots_23_io_out_uop_is_jal : _GEN_79 ? _slots_22_io_out_uop_is_jal : _slots_21_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_81 ? io_dis_uops_0_bits_is_sfb : _GEN_80 ? _slots_23_io_out_uop_is_sfb : _GEN_79 ? _slots_22_io_out_uop_is_sfb : _slots_21_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_81 ? io_dis_uops_0_bits_br_mask : _GEN_80 ? _slots_23_io_out_uop_br_mask : _GEN_79 ? _slots_22_io_out_uop_br_mask : _slots_21_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_81 ? io_dis_uops_0_bits_br_tag : _GEN_80 ? _slots_23_io_out_uop_br_tag : _GEN_79 ? _slots_22_io_out_uop_br_tag : _slots_21_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_81 ? io_dis_uops_0_bits_ftq_idx : _GEN_80 ? _slots_23_io_out_uop_ftq_idx : _GEN_79 ? _slots_22_io_out_uop_ftq_idx : _slots_21_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_81 ? io_dis_uops_0_bits_edge_inst : _GEN_80 ? _slots_23_io_out_uop_edge_inst : _GEN_79 ? _slots_22_io_out_uop_edge_inst : _slots_21_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_81 ? io_dis_uops_0_bits_pc_lob : _GEN_80 ? _slots_23_io_out_uop_pc_lob : _GEN_79 ? _slots_22_io_out_uop_pc_lob : _slots_21_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_81 ? io_dis_uops_0_bits_taken : _GEN_80 ? _slots_23_io_out_uop_taken : _GEN_79 ? _slots_22_io_out_uop_taken : _slots_21_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_81 ? io_dis_uops_0_bits_imm_packed : _GEN_80 ? _slots_23_io_out_uop_imm_packed : _GEN_79 ? _slots_22_io_out_uop_imm_packed : _slots_21_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_81 ? io_dis_uops_0_bits_csr_addr : _GEN_80 ? _slots_23_io_out_uop_csr_addr : _GEN_79 ? _slots_22_io_out_uop_csr_addr : _slots_21_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_81 ? io_dis_uops_0_bits_rob_idx : _GEN_80 ? _slots_23_io_out_uop_rob_idx : _GEN_79 ? _slots_22_io_out_uop_rob_idx : _slots_21_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_81 ? io_dis_uops_0_bits_ldq_idx : _GEN_80 ? _slots_23_io_out_uop_ldq_idx : _GEN_79 ? _slots_22_io_out_uop_ldq_idx : _slots_21_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_81 ? io_dis_uops_0_bits_stq_idx : _GEN_80 ? _slots_23_io_out_uop_stq_idx : _GEN_79 ? _slots_22_io_out_uop_stq_idx : _slots_21_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_81 ? io_dis_uops_0_bits_rxq_idx : _GEN_80 ? _slots_23_io_out_uop_rxq_idx : _GEN_79 ? _slots_22_io_out_uop_rxq_idx : _slots_21_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_81 ? io_dis_uops_0_bits_pdst : _GEN_80 ? _slots_23_io_out_uop_pdst : _GEN_79 ? _slots_22_io_out_uop_pdst : _slots_21_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_81 ? io_dis_uops_0_bits_prs1 : _GEN_80 ? _slots_23_io_out_uop_prs1 : _GEN_79 ? _slots_22_io_out_uop_prs1 : _slots_21_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_81 ? io_dis_uops_0_bits_prs2 : _GEN_80 ? _slots_23_io_out_uop_prs2 : _GEN_79 ? _slots_22_io_out_uop_prs2 : _slots_21_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_81 ? io_dis_uops_0_bits_prs3 : _GEN_80 ? _slots_23_io_out_uop_prs3 : _GEN_79 ? _slots_22_io_out_uop_prs3 : _slots_21_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_81 ? 6'h0 : _GEN_80 ? _slots_23_io_out_uop_ppred : _GEN_79 ? _slots_22_io_out_uop_ppred : _slots_21_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_81 ? io_dis_uops_0_bits_prs1_busy : _GEN_80 ? _slots_23_io_out_uop_prs1_busy : _GEN_79 ? _slots_22_io_out_uop_prs1_busy : _slots_21_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_81 ? _GEN_4 : _GEN_80 ? _slots_23_io_out_uop_prs2_busy : _GEN_79 ? _slots_22_io_out_uop_prs2_busy : _slots_21_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_81 & (_GEN_80 ? _slots_23_io_out_uop_prs3_busy : _GEN_79 ? _slots_22_io_out_uop_prs3_busy : _slots_21_io_out_uop_prs3_busy)),
    .io_in_uop_bits_ppred_busy      (~_GEN_81 & (_GEN_80 ? _slots_23_io_out_uop_ppred_busy : _GEN_79 ? _slots_22_io_out_uop_ppred_busy : _slots_21_io_out_uop_ppred_busy)),
    .io_in_uop_bits_stale_pdst      (_GEN_81 ? io_dis_uops_0_bits_stale_pdst : _GEN_80 ? _slots_23_io_out_uop_stale_pdst : _GEN_79 ? _slots_22_io_out_uop_stale_pdst : _slots_21_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_81 ? io_dis_uops_0_bits_exception : _GEN_80 ? _slots_23_io_out_uop_exception : _GEN_79 ? _slots_22_io_out_uop_exception : _slots_21_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_81 ? io_dis_uops_0_bits_exc_cause : _GEN_80 ? _slots_23_io_out_uop_exc_cause : _GEN_79 ? _slots_22_io_out_uop_exc_cause : _slots_21_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_81 ? io_dis_uops_0_bits_bypassable : _GEN_80 ? _slots_23_io_out_uop_bypassable : _GEN_79 ? _slots_22_io_out_uop_bypassable : _slots_21_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_81 ? io_dis_uops_0_bits_mem_cmd : _GEN_80 ? _slots_23_io_out_uop_mem_cmd : _GEN_79 ? _slots_22_io_out_uop_mem_cmd : _slots_21_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_81 ? io_dis_uops_0_bits_mem_size : _GEN_80 ? _slots_23_io_out_uop_mem_size : _GEN_79 ? _slots_22_io_out_uop_mem_size : _slots_21_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_81 ? io_dis_uops_0_bits_mem_signed : _GEN_80 ? _slots_23_io_out_uop_mem_signed : _GEN_79 ? _slots_22_io_out_uop_mem_signed : _slots_21_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_81 ? io_dis_uops_0_bits_is_fence : _GEN_80 ? _slots_23_io_out_uop_is_fence : _GEN_79 ? _slots_22_io_out_uop_is_fence : _slots_21_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_81 ? io_dis_uops_0_bits_is_fencei : _GEN_80 ? _slots_23_io_out_uop_is_fencei : _GEN_79 ? _slots_22_io_out_uop_is_fencei : _slots_21_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_81 ? io_dis_uops_0_bits_is_amo : _GEN_80 ? _slots_23_io_out_uop_is_amo : _GEN_79 ? _slots_22_io_out_uop_is_amo : _slots_21_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_81 ? io_dis_uops_0_bits_uses_ldq : _GEN_80 ? _slots_23_io_out_uop_uses_ldq : _GEN_79 ? _slots_22_io_out_uop_uses_ldq : _slots_21_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_81 ? io_dis_uops_0_bits_uses_stq : _GEN_80 ? _slots_23_io_out_uop_uses_stq : _GEN_79 ? _slots_22_io_out_uop_uses_stq : _slots_21_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_81 ? io_dis_uops_0_bits_is_sys_pc2epc : _GEN_80 ? _slots_23_io_out_uop_is_sys_pc2epc : _GEN_79 ? _slots_22_io_out_uop_is_sys_pc2epc : _slots_21_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_81 ? io_dis_uops_0_bits_is_unique : _GEN_80 ? _slots_23_io_out_uop_is_unique : _GEN_79 ? _slots_22_io_out_uop_is_unique : _slots_21_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_81 ? io_dis_uops_0_bits_flush_on_commit : _GEN_80 ? _slots_23_io_out_uop_flush_on_commit : _GEN_79 ? _slots_22_io_out_uop_flush_on_commit : _slots_21_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_81 ? io_dis_uops_0_bits_ldst_is_rs1 : _GEN_80 ? _slots_23_io_out_uop_ldst_is_rs1 : _GEN_79 ? _slots_22_io_out_uop_ldst_is_rs1 : _slots_21_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_81 ? io_dis_uops_0_bits_ldst : _GEN_80 ? _slots_23_io_out_uop_ldst : _GEN_79 ? _slots_22_io_out_uop_ldst : _slots_21_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_81 ? io_dis_uops_0_bits_lrs1 : _GEN_80 ? _slots_23_io_out_uop_lrs1 : _GEN_79 ? _slots_22_io_out_uop_lrs1 : _slots_21_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_81 ? io_dis_uops_0_bits_lrs2 : _GEN_80 ? _slots_23_io_out_uop_lrs2 : _GEN_79 ? _slots_22_io_out_uop_lrs2 : _slots_21_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_81 ? io_dis_uops_0_bits_lrs3 : _GEN_80 ? _slots_23_io_out_uop_lrs3 : _GEN_79 ? _slots_22_io_out_uop_lrs3 : _slots_21_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_81 ? io_dis_uops_0_bits_ldst_val : _GEN_80 ? _slots_23_io_out_uop_ldst_val : _GEN_79 ? _slots_22_io_out_uop_ldst_val : _slots_21_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_81 ? io_dis_uops_0_bits_dst_rtype : _GEN_80 ? _slots_23_io_out_uop_dst_rtype : _GEN_79 ? _slots_22_io_out_uop_dst_rtype : _slots_21_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_81 ? io_dis_uops_0_bits_lrs1_rtype : _GEN_80 ? _slots_23_io_out_uop_lrs1_rtype : _GEN_79 ? _slots_22_io_out_uop_lrs1_rtype : _slots_21_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_81 ? _GEN_3 : _GEN_80 ? _slots_23_io_out_uop_lrs2_rtype : _GEN_79 ? _slots_22_io_out_uop_lrs2_rtype : _slots_21_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_81 ? io_dis_uops_0_bits_frs3_en : _GEN_80 ? _slots_23_io_out_uop_frs3_en : _GEN_79 ? _slots_22_io_out_uop_frs3_en : _slots_21_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_81 ? io_dis_uops_0_bits_fp_val : _GEN_80 ? _slots_23_io_out_uop_fp_val : _GEN_79 ? _slots_22_io_out_uop_fp_val : _slots_21_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_81 ? io_dis_uops_0_bits_fp_single : _GEN_80 ? _slots_23_io_out_uop_fp_single : _GEN_79 ? _slots_22_io_out_uop_fp_single : _slots_21_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_81 ? io_dis_uops_0_bits_xcpt_pf_if : _GEN_80 ? _slots_23_io_out_uop_xcpt_pf_if : _GEN_79 ? _slots_22_io_out_uop_xcpt_pf_if : _slots_21_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_81 ? io_dis_uops_0_bits_xcpt_ae_if : _GEN_80 ? _slots_23_io_out_uop_xcpt_ae_if : _GEN_79 ? _slots_22_io_out_uop_xcpt_ae_if : _slots_21_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_81 ? io_dis_uops_0_bits_xcpt_ma_if : _GEN_80 ? _slots_23_io_out_uop_xcpt_ma_if : _GEN_79 ? _slots_22_io_out_uop_xcpt_ma_if : _slots_21_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_81 ? io_dis_uops_0_bits_bp_debug_if : _GEN_80 ? _slots_23_io_out_uop_bp_debug_if : _GEN_79 ? _slots_22_io_out_uop_bp_debug_if : _slots_21_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_81 ? io_dis_uops_0_bits_bp_xcpt_if : _GEN_80 ? _slots_23_io_out_uop_bp_xcpt_if : _GEN_79 ? _slots_22_io_out_uop_bp_xcpt_if : _slots_21_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_81 ? io_dis_uops_0_bits_debug_fsrc : _GEN_80 ? _slots_23_io_out_uop_debug_fsrc : _GEN_79 ? _slots_22_io_out_uop_debug_fsrc : _slots_21_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_81 ? io_dis_uops_0_bits_debug_tsrc : _GEN_80 ? _slots_23_io_out_uop_debug_tsrc : _GEN_79 ? _slots_22_io_out_uop_debug_tsrc : _slots_21_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_20_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_20_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_20_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_20_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_20_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_20_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_20_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_20_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_20_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_20_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_20_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_20_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_20_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_20_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_20_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_20_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_20_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_20_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_20_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_20_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_20_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_20_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_20_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_20_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_20_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_20_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_20_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_20_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_20_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_20_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_20_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_20_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_20_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_20_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_20_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_20_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_20_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_20_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_20_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_20_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_20_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_20_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_20_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_20_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_20_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_20_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_20_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_20_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_20_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_20_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_20_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_20_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_20_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_20_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_20_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_20_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_20_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_20_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_20_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_20_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_20_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_20_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_20_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_20_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_20_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_20_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_20_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_20_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_20_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_20_io_uop_uopc),
    .io_uop_inst                    (_slots_20_io_uop_inst),
    .io_uop_debug_inst              (_slots_20_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_20_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_20_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_20_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_20_io_uop_fu_code),
    .io_uop_iw_state                (_slots_20_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_20_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_20_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_20_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_20_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_20_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_20_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_20_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_20_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_20_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_20_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_20_io_uop_pc_lob),
    .io_uop_taken                   (_slots_20_io_uop_taken),
    .io_uop_imm_packed              (_slots_20_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_20_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_20_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_20_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_20_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_20_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_20_io_uop_pdst),
    .io_uop_prs1                    (_slots_20_io_uop_prs1),
    .io_uop_prs2                    (_slots_20_io_uop_prs2),
    .io_uop_prs3                    (_slots_20_io_uop_prs3),
    .io_uop_ppred                   (_slots_20_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_20_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_20_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_20_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_20_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_20_io_uop_stale_pdst),
    .io_uop_exception               (_slots_20_io_uop_exception),
    .io_uop_exc_cause               (_slots_20_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_20_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_20_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_20_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_20_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_20_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_20_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_20_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_20_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_20_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_20_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_20_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_20_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_20_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_20_io_uop_ldst),
    .io_uop_lrs1                    (_slots_20_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_20_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_20_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_20_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_20_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_20_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_20_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_20_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_20_io_uop_fp_val),
    .io_uop_fp_single               (_slots_20_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_20_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_20_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_20_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_20_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_20_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_20_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_20_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_21 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_21_io_valid),
    .io_will_be_valid               (_slots_21_io_will_be_valid),
    .io_request                     (_slots_21_io_request),
    .io_grant                       (issue_slots_21_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_20),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_21_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_84 ? io_dis_uops_1_bits_uopc : _GEN_83 ? io_dis_uops_0_bits_uopc : _GEN_82 ? _slots_23_io_out_uop_uopc : _slots_22_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_84 ? io_dis_uops_1_bits_inst : _GEN_83 ? io_dis_uops_0_bits_inst : _GEN_82 ? _slots_23_io_out_uop_inst : _slots_22_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_84 ? io_dis_uops_1_bits_debug_inst : _GEN_83 ? io_dis_uops_0_bits_debug_inst : _GEN_82 ? _slots_23_io_out_uop_debug_inst : _slots_22_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_84 ? io_dis_uops_1_bits_is_rvc : _GEN_83 ? io_dis_uops_0_bits_is_rvc : _GEN_82 ? _slots_23_io_out_uop_is_rvc : _slots_22_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_84 ? io_dis_uops_1_bits_debug_pc : _GEN_83 ? io_dis_uops_0_bits_debug_pc : _GEN_82 ? _slots_23_io_out_uop_debug_pc : _slots_22_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_84 ? io_dis_uops_1_bits_iq_type : _GEN_83 ? io_dis_uops_0_bits_iq_type : _GEN_82 ? _slots_23_io_out_uop_iq_type : _slots_22_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_84 ? io_dis_uops_1_bits_fu_code : _GEN_83 ? io_dis_uops_0_bits_fu_code : _GEN_82 ? _slots_23_io_out_uop_fu_code : _slots_22_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_84 ? _GEN_7 : _GEN_83 ? _GEN_1 : _GEN_82 ? _slots_23_io_out_uop_iw_state : _slots_22_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_85 & (_GEN_82 ? _slots_23_io_out_uop_iw_p1_poisoned : _slots_22_io_out_uop_iw_p1_poisoned)),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_85 & (_GEN_82 ? _slots_23_io_out_uop_iw_p2_poisoned : _slots_22_io_out_uop_iw_p2_poisoned)),
    .io_in_uop_bits_is_br           (_GEN_84 ? io_dis_uops_1_bits_is_br : _GEN_83 ? io_dis_uops_0_bits_is_br : _GEN_82 ? _slots_23_io_out_uop_is_br : _slots_22_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_84 ? io_dis_uops_1_bits_is_jalr : _GEN_83 ? io_dis_uops_0_bits_is_jalr : _GEN_82 ? _slots_23_io_out_uop_is_jalr : _slots_22_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_84 ? io_dis_uops_1_bits_is_jal : _GEN_83 ? io_dis_uops_0_bits_is_jal : _GEN_82 ? _slots_23_io_out_uop_is_jal : _slots_22_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_84 ? io_dis_uops_1_bits_is_sfb : _GEN_83 ? io_dis_uops_0_bits_is_sfb : _GEN_82 ? _slots_23_io_out_uop_is_sfb : _slots_22_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_84 ? io_dis_uops_1_bits_br_mask : _GEN_83 ? io_dis_uops_0_bits_br_mask : _GEN_82 ? _slots_23_io_out_uop_br_mask : _slots_22_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_84 ? io_dis_uops_1_bits_br_tag : _GEN_83 ? io_dis_uops_0_bits_br_tag : _GEN_82 ? _slots_23_io_out_uop_br_tag : _slots_22_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_84 ? io_dis_uops_1_bits_ftq_idx : _GEN_83 ? io_dis_uops_0_bits_ftq_idx : _GEN_82 ? _slots_23_io_out_uop_ftq_idx : _slots_22_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_84 ? io_dis_uops_1_bits_edge_inst : _GEN_83 ? io_dis_uops_0_bits_edge_inst : _GEN_82 ? _slots_23_io_out_uop_edge_inst : _slots_22_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_84 ? io_dis_uops_1_bits_pc_lob : _GEN_83 ? io_dis_uops_0_bits_pc_lob : _GEN_82 ? _slots_23_io_out_uop_pc_lob : _slots_22_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_84 ? io_dis_uops_1_bits_taken : _GEN_83 ? io_dis_uops_0_bits_taken : _GEN_82 ? _slots_23_io_out_uop_taken : _slots_22_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_84 ? io_dis_uops_1_bits_imm_packed : _GEN_83 ? io_dis_uops_0_bits_imm_packed : _GEN_82 ? _slots_23_io_out_uop_imm_packed : _slots_22_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_84 ? io_dis_uops_1_bits_csr_addr : _GEN_83 ? io_dis_uops_0_bits_csr_addr : _GEN_82 ? _slots_23_io_out_uop_csr_addr : _slots_22_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_84 ? io_dis_uops_1_bits_rob_idx : _GEN_83 ? io_dis_uops_0_bits_rob_idx : _GEN_82 ? _slots_23_io_out_uop_rob_idx : _slots_22_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_84 ? io_dis_uops_1_bits_ldq_idx : _GEN_83 ? io_dis_uops_0_bits_ldq_idx : _GEN_82 ? _slots_23_io_out_uop_ldq_idx : _slots_22_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_84 ? io_dis_uops_1_bits_stq_idx : _GEN_83 ? io_dis_uops_0_bits_stq_idx : _GEN_82 ? _slots_23_io_out_uop_stq_idx : _slots_22_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_84 ? io_dis_uops_1_bits_rxq_idx : _GEN_83 ? io_dis_uops_0_bits_rxq_idx : _GEN_82 ? _slots_23_io_out_uop_rxq_idx : _slots_22_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_84 ? io_dis_uops_1_bits_pdst : _GEN_83 ? io_dis_uops_0_bits_pdst : _GEN_82 ? _slots_23_io_out_uop_pdst : _slots_22_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_84 ? io_dis_uops_1_bits_prs1 : _GEN_83 ? io_dis_uops_0_bits_prs1 : _GEN_82 ? _slots_23_io_out_uop_prs1 : _slots_22_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_84 ? io_dis_uops_1_bits_prs2 : _GEN_83 ? io_dis_uops_0_bits_prs2 : _GEN_82 ? _slots_23_io_out_uop_prs2 : _slots_22_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_84 ? io_dis_uops_1_bits_prs3 : _GEN_83 ? io_dis_uops_0_bits_prs3 : _GEN_82 ? _slots_23_io_out_uop_prs3 : _slots_22_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_85 ? 6'h0 : _GEN_82 ? _slots_23_io_out_uop_ppred : _slots_22_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_84 ? io_dis_uops_1_bits_prs1_busy : _GEN_83 ? io_dis_uops_0_bits_prs1_busy : _GEN_82 ? _slots_23_io_out_uop_prs1_busy : _slots_22_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_84 ? _GEN_10 : _GEN_83 ? _GEN_4 : _GEN_82 ? _slots_23_io_out_uop_prs2_busy : _slots_22_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_85 & (_GEN_82 ? _slots_23_io_out_uop_prs3_busy : _slots_22_io_out_uop_prs3_busy)),
    .io_in_uop_bits_ppred_busy      (~_GEN_85 & (_GEN_82 ? _slots_23_io_out_uop_ppred_busy : _slots_22_io_out_uop_ppred_busy)),
    .io_in_uop_bits_stale_pdst      (_GEN_84 ? io_dis_uops_1_bits_stale_pdst : _GEN_83 ? io_dis_uops_0_bits_stale_pdst : _GEN_82 ? _slots_23_io_out_uop_stale_pdst : _slots_22_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_84 ? io_dis_uops_1_bits_exception : _GEN_83 ? io_dis_uops_0_bits_exception : _GEN_82 ? _slots_23_io_out_uop_exception : _slots_22_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_84 ? io_dis_uops_1_bits_exc_cause : _GEN_83 ? io_dis_uops_0_bits_exc_cause : _GEN_82 ? _slots_23_io_out_uop_exc_cause : _slots_22_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_84 ? io_dis_uops_1_bits_bypassable : _GEN_83 ? io_dis_uops_0_bits_bypassable : _GEN_82 ? _slots_23_io_out_uop_bypassable : _slots_22_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_84 ? io_dis_uops_1_bits_mem_cmd : _GEN_83 ? io_dis_uops_0_bits_mem_cmd : _GEN_82 ? _slots_23_io_out_uop_mem_cmd : _slots_22_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_84 ? io_dis_uops_1_bits_mem_size : _GEN_83 ? io_dis_uops_0_bits_mem_size : _GEN_82 ? _slots_23_io_out_uop_mem_size : _slots_22_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_84 ? io_dis_uops_1_bits_mem_signed : _GEN_83 ? io_dis_uops_0_bits_mem_signed : _GEN_82 ? _slots_23_io_out_uop_mem_signed : _slots_22_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_84 ? io_dis_uops_1_bits_is_fence : _GEN_83 ? io_dis_uops_0_bits_is_fence : _GEN_82 ? _slots_23_io_out_uop_is_fence : _slots_22_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_84 ? io_dis_uops_1_bits_is_fencei : _GEN_83 ? io_dis_uops_0_bits_is_fencei : _GEN_82 ? _slots_23_io_out_uop_is_fencei : _slots_22_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_84 ? io_dis_uops_1_bits_is_amo : _GEN_83 ? io_dis_uops_0_bits_is_amo : _GEN_82 ? _slots_23_io_out_uop_is_amo : _slots_22_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_84 ? io_dis_uops_1_bits_uses_ldq : _GEN_83 ? io_dis_uops_0_bits_uses_ldq : _GEN_82 ? _slots_23_io_out_uop_uses_ldq : _slots_22_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_84 ? io_dis_uops_1_bits_uses_stq : _GEN_83 ? io_dis_uops_0_bits_uses_stq : _GEN_82 ? _slots_23_io_out_uop_uses_stq : _slots_22_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_84 ? io_dis_uops_1_bits_is_sys_pc2epc : _GEN_83 ? io_dis_uops_0_bits_is_sys_pc2epc : _GEN_82 ? _slots_23_io_out_uop_is_sys_pc2epc : _slots_22_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_84 ? io_dis_uops_1_bits_is_unique : _GEN_83 ? io_dis_uops_0_bits_is_unique : _GEN_82 ? _slots_23_io_out_uop_is_unique : _slots_22_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_84 ? io_dis_uops_1_bits_flush_on_commit : _GEN_83 ? io_dis_uops_0_bits_flush_on_commit : _GEN_82 ? _slots_23_io_out_uop_flush_on_commit : _slots_22_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_84 ? io_dis_uops_1_bits_ldst_is_rs1 : _GEN_83 ? io_dis_uops_0_bits_ldst_is_rs1 : _GEN_82 ? _slots_23_io_out_uop_ldst_is_rs1 : _slots_22_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_84 ? io_dis_uops_1_bits_ldst : _GEN_83 ? io_dis_uops_0_bits_ldst : _GEN_82 ? _slots_23_io_out_uop_ldst : _slots_22_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_84 ? io_dis_uops_1_bits_lrs1 : _GEN_83 ? io_dis_uops_0_bits_lrs1 : _GEN_82 ? _slots_23_io_out_uop_lrs1 : _slots_22_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_84 ? io_dis_uops_1_bits_lrs2 : _GEN_83 ? io_dis_uops_0_bits_lrs2 : _GEN_82 ? _slots_23_io_out_uop_lrs2 : _slots_22_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_84 ? io_dis_uops_1_bits_lrs3 : _GEN_83 ? io_dis_uops_0_bits_lrs3 : _GEN_82 ? _slots_23_io_out_uop_lrs3 : _slots_22_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_84 ? io_dis_uops_1_bits_ldst_val : _GEN_83 ? io_dis_uops_0_bits_ldst_val : _GEN_82 ? _slots_23_io_out_uop_ldst_val : _slots_22_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_84 ? io_dis_uops_1_bits_dst_rtype : _GEN_83 ? io_dis_uops_0_bits_dst_rtype : _GEN_82 ? _slots_23_io_out_uop_dst_rtype : _slots_22_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_84 ? io_dis_uops_1_bits_lrs1_rtype : _GEN_83 ? io_dis_uops_0_bits_lrs1_rtype : _GEN_82 ? _slots_23_io_out_uop_lrs1_rtype : _slots_22_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_84 ? _GEN_9 : _GEN_83 ? _GEN_3 : _GEN_82 ? _slots_23_io_out_uop_lrs2_rtype : _slots_22_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_84 ? io_dis_uops_1_bits_frs3_en : _GEN_83 ? io_dis_uops_0_bits_frs3_en : _GEN_82 ? _slots_23_io_out_uop_frs3_en : _slots_22_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_84 ? io_dis_uops_1_bits_fp_val : _GEN_83 ? io_dis_uops_0_bits_fp_val : _GEN_82 ? _slots_23_io_out_uop_fp_val : _slots_22_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_84 ? io_dis_uops_1_bits_fp_single : _GEN_83 ? io_dis_uops_0_bits_fp_single : _GEN_82 ? _slots_23_io_out_uop_fp_single : _slots_22_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_84 ? io_dis_uops_1_bits_xcpt_pf_if : _GEN_83 ? io_dis_uops_0_bits_xcpt_pf_if : _GEN_82 ? _slots_23_io_out_uop_xcpt_pf_if : _slots_22_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_84 ? io_dis_uops_1_bits_xcpt_ae_if : _GEN_83 ? io_dis_uops_0_bits_xcpt_ae_if : _GEN_82 ? _slots_23_io_out_uop_xcpt_ae_if : _slots_22_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_84 ? io_dis_uops_1_bits_xcpt_ma_if : _GEN_83 ? io_dis_uops_0_bits_xcpt_ma_if : _GEN_82 ? _slots_23_io_out_uop_xcpt_ma_if : _slots_22_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_84 ? io_dis_uops_1_bits_bp_debug_if : _GEN_83 ? io_dis_uops_0_bits_bp_debug_if : _GEN_82 ? _slots_23_io_out_uop_bp_debug_if : _slots_22_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_84 ? io_dis_uops_1_bits_bp_xcpt_if : _GEN_83 ? io_dis_uops_0_bits_bp_xcpt_if : _GEN_82 ? _slots_23_io_out_uop_bp_xcpt_if : _slots_22_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_84 ? io_dis_uops_1_bits_debug_fsrc : _GEN_83 ? io_dis_uops_0_bits_debug_fsrc : _GEN_82 ? _slots_23_io_out_uop_debug_fsrc : _slots_22_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_84 ? io_dis_uops_1_bits_debug_tsrc : _GEN_83 ? io_dis_uops_0_bits_debug_tsrc : _GEN_82 ? _slots_23_io_out_uop_debug_tsrc : _slots_22_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_21_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_21_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_21_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_21_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_21_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_21_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_21_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_21_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_21_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_21_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_21_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_21_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_21_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_21_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_21_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_21_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_21_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_21_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_21_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_21_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_21_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_21_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_21_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_21_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_21_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_21_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_21_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_21_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_21_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_21_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_21_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_21_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_21_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_21_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_21_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_21_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_21_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_21_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_21_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_21_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_21_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_21_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_21_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_21_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_21_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_21_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_21_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_21_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_21_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_21_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_21_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_21_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_21_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_21_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_21_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_21_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_21_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_21_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_21_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_21_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_21_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_21_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_21_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_21_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_21_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_21_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_21_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_21_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_21_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_21_io_uop_uopc),
    .io_uop_inst                    (_slots_21_io_uop_inst),
    .io_uop_debug_inst              (_slots_21_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_21_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_21_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_21_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_21_io_uop_fu_code),
    .io_uop_iw_state                (_slots_21_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_21_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_21_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_21_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_21_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_21_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_21_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_21_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_21_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_21_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_21_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_21_io_uop_pc_lob),
    .io_uop_taken                   (_slots_21_io_uop_taken),
    .io_uop_imm_packed              (_slots_21_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_21_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_21_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_21_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_21_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_21_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_21_io_uop_pdst),
    .io_uop_prs1                    (_slots_21_io_uop_prs1),
    .io_uop_prs2                    (_slots_21_io_uop_prs2),
    .io_uop_prs3                    (_slots_21_io_uop_prs3),
    .io_uop_ppred                   (_slots_21_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_21_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_21_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_21_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_21_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_21_io_uop_stale_pdst),
    .io_uop_exception               (_slots_21_io_uop_exception),
    .io_uop_exc_cause               (_slots_21_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_21_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_21_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_21_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_21_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_21_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_21_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_21_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_21_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_21_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_21_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_21_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_21_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_21_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_21_io_uop_ldst),
    .io_uop_lrs1                    (_slots_21_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_21_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_21_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_21_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_21_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_21_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_21_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_21_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_21_io_uop_fp_val),
    .io_uop_fp_single               (_slots_21_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_21_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_21_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_21_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_21_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_21_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_21_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_21_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_22 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_22_io_valid),
    .io_will_be_valid               (_slots_22_io_will_be_valid),
    .io_request                     (_slots_22_io_request),
    .io_grant                       (issue_slots_22_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_21),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_22_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_88 ? io_dis_uops_2_bits_uopc : _GEN_87 ? io_dis_uops_1_bits_uopc : _GEN_86 ? io_dis_uops_0_bits_uopc : _slots_23_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_88 ? io_dis_uops_2_bits_inst : _GEN_87 ? io_dis_uops_1_bits_inst : _GEN_86 ? io_dis_uops_0_bits_inst : _slots_23_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_88 ? io_dis_uops_2_bits_debug_inst : _GEN_87 ? io_dis_uops_1_bits_debug_inst : _GEN_86 ? io_dis_uops_0_bits_debug_inst : _slots_23_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_88 ? io_dis_uops_2_bits_is_rvc : _GEN_87 ? io_dis_uops_1_bits_is_rvc : _GEN_86 ? io_dis_uops_0_bits_is_rvc : _slots_23_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_88 ? io_dis_uops_2_bits_debug_pc : _GEN_87 ? io_dis_uops_1_bits_debug_pc : _GEN_86 ? io_dis_uops_0_bits_debug_pc : _slots_23_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_88 ? io_dis_uops_2_bits_iq_type : _GEN_87 ? io_dis_uops_1_bits_iq_type : _GEN_86 ? io_dis_uops_0_bits_iq_type : _slots_23_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_88 ? io_dis_uops_2_bits_fu_code : _GEN_87 ? io_dis_uops_1_bits_fu_code : _GEN_86 ? io_dis_uops_0_bits_fu_code : _slots_23_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_88 ? (_GEN_12 ? 2'h2 : 2'h1) : _GEN_87 ? _GEN_7 : _GEN_86 ? _GEN_1 : _slots_23_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_89 & _slots_23_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_89 & _slots_23_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_88 ? io_dis_uops_2_bits_is_br : _GEN_87 ? io_dis_uops_1_bits_is_br : _GEN_86 ? io_dis_uops_0_bits_is_br : _slots_23_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_88 ? io_dis_uops_2_bits_is_jalr : _GEN_87 ? io_dis_uops_1_bits_is_jalr : _GEN_86 ? io_dis_uops_0_bits_is_jalr : _slots_23_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_88 ? io_dis_uops_2_bits_is_jal : _GEN_87 ? io_dis_uops_1_bits_is_jal : _GEN_86 ? io_dis_uops_0_bits_is_jal : _slots_23_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_88 ? io_dis_uops_2_bits_is_sfb : _GEN_87 ? io_dis_uops_1_bits_is_sfb : _GEN_86 ? io_dis_uops_0_bits_is_sfb : _slots_23_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_88 ? io_dis_uops_2_bits_br_mask : _GEN_87 ? io_dis_uops_1_bits_br_mask : _GEN_86 ? io_dis_uops_0_bits_br_mask : _slots_23_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_88 ? io_dis_uops_2_bits_br_tag : _GEN_87 ? io_dis_uops_1_bits_br_tag : _GEN_86 ? io_dis_uops_0_bits_br_tag : _slots_23_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_88 ? io_dis_uops_2_bits_ftq_idx : _GEN_87 ? io_dis_uops_1_bits_ftq_idx : _GEN_86 ? io_dis_uops_0_bits_ftq_idx : _slots_23_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_88 ? io_dis_uops_2_bits_edge_inst : _GEN_87 ? io_dis_uops_1_bits_edge_inst : _GEN_86 ? io_dis_uops_0_bits_edge_inst : _slots_23_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_88 ? io_dis_uops_2_bits_pc_lob : _GEN_87 ? io_dis_uops_1_bits_pc_lob : _GEN_86 ? io_dis_uops_0_bits_pc_lob : _slots_23_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_88 ? io_dis_uops_2_bits_taken : _GEN_87 ? io_dis_uops_1_bits_taken : _GEN_86 ? io_dis_uops_0_bits_taken : _slots_23_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_88 ? io_dis_uops_2_bits_imm_packed : _GEN_87 ? io_dis_uops_1_bits_imm_packed : _GEN_86 ? io_dis_uops_0_bits_imm_packed : _slots_23_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_88 ? io_dis_uops_2_bits_csr_addr : _GEN_87 ? io_dis_uops_1_bits_csr_addr : _GEN_86 ? io_dis_uops_0_bits_csr_addr : _slots_23_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_88 ? io_dis_uops_2_bits_rob_idx : _GEN_87 ? io_dis_uops_1_bits_rob_idx : _GEN_86 ? io_dis_uops_0_bits_rob_idx : _slots_23_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_88 ? io_dis_uops_2_bits_ldq_idx : _GEN_87 ? io_dis_uops_1_bits_ldq_idx : _GEN_86 ? io_dis_uops_0_bits_ldq_idx : _slots_23_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_88 ? io_dis_uops_2_bits_stq_idx : _GEN_87 ? io_dis_uops_1_bits_stq_idx : _GEN_86 ? io_dis_uops_0_bits_stq_idx : _slots_23_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_88 ? io_dis_uops_2_bits_rxq_idx : _GEN_87 ? io_dis_uops_1_bits_rxq_idx : _GEN_86 ? io_dis_uops_0_bits_rxq_idx : _slots_23_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_88 ? io_dis_uops_2_bits_pdst : _GEN_87 ? io_dis_uops_1_bits_pdst : _GEN_86 ? io_dis_uops_0_bits_pdst : _slots_23_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_88 ? io_dis_uops_2_bits_prs1 : _GEN_87 ? io_dis_uops_1_bits_prs1 : _GEN_86 ? io_dis_uops_0_bits_prs1 : _slots_23_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_88 ? io_dis_uops_2_bits_prs2 : _GEN_87 ? io_dis_uops_1_bits_prs2 : _GEN_86 ? io_dis_uops_0_bits_prs2 : _slots_23_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_88 ? io_dis_uops_2_bits_prs3 : _GEN_87 ? io_dis_uops_1_bits_prs3 : _GEN_86 ? io_dis_uops_0_bits_prs3 : _slots_23_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_89 ? 6'h0 : _slots_23_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_88 ? io_dis_uops_2_bits_prs1_busy : _GEN_87 ? io_dis_uops_1_bits_prs1_busy : _GEN_86 ? io_dis_uops_0_bits_prs1_busy : _slots_23_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_88 ? _GEN_15 : _GEN_87 ? _GEN_10 : _GEN_86 ? _GEN_4 : _slots_23_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_89 & _slots_23_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (~_GEN_89 & _slots_23_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_88 ? io_dis_uops_2_bits_stale_pdst : _GEN_87 ? io_dis_uops_1_bits_stale_pdst : _GEN_86 ? io_dis_uops_0_bits_stale_pdst : _slots_23_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_88 ? io_dis_uops_2_bits_exception : _GEN_87 ? io_dis_uops_1_bits_exception : _GEN_86 ? io_dis_uops_0_bits_exception : _slots_23_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_88 ? io_dis_uops_2_bits_exc_cause : _GEN_87 ? io_dis_uops_1_bits_exc_cause : _GEN_86 ? io_dis_uops_0_bits_exc_cause : _slots_23_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_88 ? io_dis_uops_2_bits_bypassable : _GEN_87 ? io_dis_uops_1_bits_bypassable : _GEN_86 ? io_dis_uops_0_bits_bypassable : _slots_23_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_88 ? io_dis_uops_2_bits_mem_cmd : _GEN_87 ? io_dis_uops_1_bits_mem_cmd : _GEN_86 ? io_dis_uops_0_bits_mem_cmd : _slots_23_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_88 ? io_dis_uops_2_bits_mem_size : _GEN_87 ? io_dis_uops_1_bits_mem_size : _GEN_86 ? io_dis_uops_0_bits_mem_size : _slots_23_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_88 ? io_dis_uops_2_bits_mem_signed : _GEN_87 ? io_dis_uops_1_bits_mem_signed : _GEN_86 ? io_dis_uops_0_bits_mem_signed : _slots_23_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_88 ? io_dis_uops_2_bits_is_fence : _GEN_87 ? io_dis_uops_1_bits_is_fence : _GEN_86 ? io_dis_uops_0_bits_is_fence : _slots_23_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_88 ? io_dis_uops_2_bits_is_fencei : _GEN_87 ? io_dis_uops_1_bits_is_fencei : _GEN_86 ? io_dis_uops_0_bits_is_fencei : _slots_23_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_88 ? io_dis_uops_2_bits_is_amo : _GEN_87 ? io_dis_uops_1_bits_is_amo : _GEN_86 ? io_dis_uops_0_bits_is_amo : _slots_23_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_88 ? io_dis_uops_2_bits_uses_ldq : _GEN_87 ? io_dis_uops_1_bits_uses_ldq : _GEN_86 ? io_dis_uops_0_bits_uses_ldq : _slots_23_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_88 ? io_dis_uops_2_bits_uses_stq : _GEN_87 ? io_dis_uops_1_bits_uses_stq : _GEN_86 ? io_dis_uops_0_bits_uses_stq : _slots_23_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_88 ? io_dis_uops_2_bits_is_sys_pc2epc : _GEN_87 ? io_dis_uops_1_bits_is_sys_pc2epc : _GEN_86 ? io_dis_uops_0_bits_is_sys_pc2epc : _slots_23_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_88 ? io_dis_uops_2_bits_is_unique : _GEN_87 ? io_dis_uops_1_bits_is_unique : _GEN_86 ? io_dis_uops_0_bits_is_unique : _slots_23_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_88 ? io_dis_uops_2_bits_flush_on_commit : _GEN_87 ? io_dis_uops_1_bits_flush_on_commit : _GEN_86 ? io_dis_uops_0_bits_flush_on_commit : _slots_23_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_88 ? io_dis_uops_2_bits_ldst_is_rs1 : _GEN_87 ? io_dis_uops_1_bits_ldst_is_rs1 : _GEN_86 ? io_dis_uops_0_bits_ldst_is_rs1 : _slots_23_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_88 ? io_dis_uops_2_bits_ldst : _GEN_87 ? io_dis_uops_1_bits_ldst : _GEN_86 ? io_dis_uops_0_bits_ldst : _slots_23_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_88 ? io_dis_uops_2_bits_lrs1 : _GEN_87 ? io_dis_uops_1_bits_lrs1 : _GEN_86 ? io_dis_uops_0_bits_lrs1 : _slots_23_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_88 ? io_dis_uops_2_bits_lrs2 : _GEN_87 ? io_dis_uops_1_bits_lrs2 : _GEN_86 ? io_dis_uops_0_bits_lrs2 : _slots_23_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_88 ? io_dis_uops_2_bits_lrs3 : _GEN_87 ? io_dis_uops_1_bits_lrs3 : _GEN_86 ? io_dis_uops_0_bits_lrs3 : _slots_23_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_88 ? io_dis_uops_2_bits_ldst_val : _GEN_87 ? io_dis_uops_1_bits_ldst_val : _GEN_86 ? io_dis_uops_0_bits_ldst_val : _slots_23_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_88 ? io_dis_uops_2_bits_dst_rtype : _GEN_87 ? io_dis_uops_1_bits_dst_rtype : _GEN_86 ? io_dis_uops_0_bits_dst_rtype : _slots_23_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_88 ? io_dis_uops_2_bits_lrs1_rtype : _GEN_87 ? io_dis_uops_1_bits_lrs1_rtype : _GEN_86 ? io_dis_uops_0_bits_lrs1_rtype : _slots_23_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_88 ? _GEN_14 : _GEN_87 ? _GEN_9 : _GEN_86 ? _GEN_3 : _slots_23_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_88 ? io_dis_uops_2_bits_frs3_en : _GEN_87 ? io_dis_uops_1_bits_frs3_en : _GEN_86 ? io_dis_uops_0_bits_frs3_en : _slots_23_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_88 ? io_dis_uops_2_bits_fp_val : _GEN_87 ? io_dis_uops_1_bits_fp_val : _GEN_86 ? io_dis_uops_0_bits_fp_val : _slots_23_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_88 ? io_dis_uops_2_bits_fp_single : _GEN_87 ? io_dis_uops_1_bits_fp_single : _GEN_86 ? io_dis_uops_0_bits_fp_single : _slots_23_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_88 ? io_dis_uops_2_bits_xcpt_pf_if : _GEN_87 ? io_dis_uops_1_bits_xcpt_pf_if : _GEN_86 ? io_dis_uops_0_bits_xcpt_pf_if : _slots_23_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_88 ? io_dis_uops_2_bits_xcpt_ae_if : _GEN_87 ? io_dis_uops_1_bits_xcpt_ae_if : _GEN_86 ? io_dis_uops_0_bits_xcpt_ae_if : _slots_23_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_88 ? io_dis_uops_2_bits_xcpt_ma_if : _GEN_87 ? io_dis_uops_1_bits_xcpt_ma_if : _GEN_86 ? io_dis_uops_0_bits_xcpt_ma_if : _slots_23_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_88 ? io_dis_uops_2_bits_bp_debug_if : _GEN_87 ? io_dis_uops_1_bits_bp_debug_if : _GEN_86 ? io_dis_uops_0_bits_bp_debug_if : _slots_23_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_88 ? io_dis_uops_2_bits_bp_xcpt_if : _GEN_87 ? io_dis_uops_1_bits_bp_xcpt_if : _GEN_86 ? io_dis_uops_0_bits_bp_xcpt_if : _slots_23_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_88 ? io_dis_uops_2_bits_debug_fsrc : _GEN_87 ? io_dis_uops_1_bits_debug_fsrc : _GEN_86 ? io_dis_uops_0_bits_debug_fsrc : _slots_23_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_88 ? io_dis_uops_2_bits_debug_tsrc : _GEN_87 ? io_dis_uops_1_bits_debug_tsrc : _GEN_86 ? io_dis_uops_0_bits_debug_tsrc : _slots_23_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_22_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_22_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_22_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_22_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_22_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_22_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_22_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_22_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_22_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_22_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_22_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_22_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_22_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_22_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_22_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_22_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_22_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_22_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_22_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_22_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_22_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_22_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_22_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_22_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_22_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_22_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_22_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_22_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_22_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_22_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_22_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_22_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_22_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_22_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_22_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_22_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_22_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_22_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_22_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_22_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_22_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_22_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_22_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_22_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_22_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_22_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_22_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_22_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_22_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_22_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_22_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_22_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_22_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_22_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_22_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_22_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_22_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_22_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_22_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_22_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_22_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_22_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_22_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_22_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_22_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_22_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_22_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_22_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_22_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_22_io_uop_uopc),
    .io_uop_inst                    (_slots_22_io_uop_inst),
    .io_uop_debug_inst              (_slots_22_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_22_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_22_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_22_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_22_io_uop_fu_code),
    .io_uop_iw_state                (_slots_22_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_22_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_22_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_22_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_22_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_22_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_22_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_22_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_22_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_22_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_22_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_22_io_uop_pc_lob),
    .io_uop_taken                   (_slots_22_io_uop_taken),
    .io_uop_imm_packed              (_slots_22_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_22_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_22_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_22_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_22_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_22_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_22_io_uop_pdst),
    .io_uop_prs1                    (_slots_22_io_uop_prs1),
    .io_uop_prs2                    (_slots_22_io_uop_prs2),
    .io_uop_prs3                    (_slots_22_io_uop_prs3),
    .io_uop_ppred                   (_slots_22_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_22_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_22_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_22_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_22_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_22_io_uop_stale_pdst),
    .io_uop_exception               (_slots_22_io_uop_exception),
    .io_uop_exc_cause               (_slots_22_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_22_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_22_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_22_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_22_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_22_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_22_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_22_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_22_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_22_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_22_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_22_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_22_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_22_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_22_io_uop_ldst),
    .io_uop_lrs1                    (_slots_22_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_22_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_22_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_22_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_22_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_22_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_22_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_22_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_22_io_uop_fp_val),
    .io_uop_fp_single               (_slots_22_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_22_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_22_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_22_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_22_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_22_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_22_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_22_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_23 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_23_io_valid),
    .io_will_be_valid               (_slots_23_io_will_be_valid),
    .io_request                     (_slots_23_io_request),
    .io_grant                       (issue_slots_23_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_22),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_23_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_92 ? io_dis_uops_3_bits_uopc : _GEN_91 ? io_dis_uops_2_bits_uopc : _GEN_90 ? io_dis_uops_1_bits_uopc : io_dis_uops_0_bits_uopc),
    .io_in_uop_bits_inst            (_GEN_92 ? io_dis_uops_3_bits_inst : _GEN_91 ? io_dis_uops_2_bits_inst : _GEN_90 ? io_dis_uops_1_bits_inst : io_dis_uops_0_bits_inst),
    .io_in_uop_bits_debug_inst      (_GEN_92 ? io_dis_uops_3_bits_debug_inst : _GEN_91 ? io_dis_uops_2_bits_debug_inst : _GEN_90 ? io_dis_uops_1_bits_debug_inst : io_dis_uops_0_bits_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_92 ? io_dis_uops_3_bits_is_rvc : _GEN_91 ? io_dis_uops_2_bits_is_rvc : _GEN_90 ? io_dis_uops_1_bits_is_rvc : io_dis_uops_0_bits_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_92 ? io_dis_uops_3_bits_debug_pc : _GEN_91 ? io_dis_uops_2_bits_debug_pc : _GEN_90 ? io_dis_uops_1_bits_debug_pc : io_dis_uops_0_bits_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_92 ? io_dis_uops_3_bits_iq_type : _GEN_91 ? io_dis_uops_2_bits_iq_type : _GEN_90 ? io_dis_uops_1_bits_iq_type : io_dis_uops_0_bits_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_92 ? io_dis_uops_3_bits_fu_code : _GEN_91 ? io_dis_uops_2_bits_fu_code : _GEN_90 ? io_dis_uops_1_bits_fu_code : io_dis_uops_0_bits_fu_code),
    .io_in_uop_bits_iw_state        ((_GEN_92 ? _GEN_17 : _GEN_91 ? _GEN_12 : _GEN_90 ? _GEN_6 : _GEN_0) ? 2'h2 : 2'h1),
    .io_in_uop_bits_iw_p1_poisoned  (1'h0),
    .io_in_uop_bits_iw_p2_poisoned  (1'h0),
    .io_in_uop_bits_is_br           (_GEN_92 ? io_dis_uops_3_bits_is_br : _GEN_91 ? io_dis_uops_2_bits_is_br : _GEN_90 ? io_dis_uops_1_bits_is_br : io_dis_uops_0_bits_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_92 ? io_dis_uops_3_bits_is_jalr : _GEN_91 ? io_dis_uops_2_bits_is_jalr : _GEN_90 ? io_dis_uops_1_bits_is_jalr : io_dis_uops_0_bits_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_92 ? io_dis_uops_3_bits_is_jal : _GEN_91 ? io_dis_uops_2_bits_is_jal : _GEN_90 ? io_dis_uops_1_bits_is_jal : io_dis_uops_0_bits_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_92 ? io_dis_uops_3_bits_is_sfb : _GEN_91 ? io_dis_uops_2_bits_is_sfb : _GEN_90 ? io_dis_uops_1_bits_is_sfb : io_dis_uops_0_bits_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_92 ? io_dis_uops_3_bits_br_mask : _GEN_91 ? io_dis_uops_2_bits_br_mask : _GEN_90 ? io_dis_uops_1_bits_br_mask : io_dis_uops_0_bits_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_92 ? io_dis_uops_3_bits_br_tag : _GEN_91 ? io_dis_uops_2_bits_br_tag : _GEN_90 ? io_dis_uops_1_bits_br_tag : io_dis_uops_0_bits_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_92 ? io_dis_uops_3_bits_ftq_idx : _GEN_91 ? io_dis_uops_2_bits_ftq_idx : _GEN_90 ? io_dis_uops_1_bits_ftq_idx : io_dis_uops_0_bits_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_92 ? io_dis_uops_3_bits_edge_inst : _GEN_91 ? io_dis_uops_2_bits_edge_inst : _GEN_90 ? io_dis_uops_1_bits_edge_inst : io_dis_uops_0_bits_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_92 ? io_dis_uops_3_bits_pc_lob : _GEN_91 ? io_dis_uops_2_bits_pc_lob : _GEN_90 ? io_dis_uops_1_bits_pc_lob : io_dis_uops_0_bits_pc_lob),
    .io_in_uop_bits_taken           (_GEN_92 ? io_dis_uops_3_bits_taken : _GEN_91 ? io_dis_uops_2_bits_taken : _GEN_90 ? io_dis_uops_1_bits_taken : io_dis_uops_0_bits_taken),
    .io_in_uop_bits_imm_packed      (_GEN_92 ? io_dis_uops_3_bits_imm_packed : _GEN_91 ? io_dis_uops_2_bits_imm_packed : _GEN_90 ? io_dis_uops_1_bits_imm_packed : io_dis_uops_0_bits_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_92 ? io_dis_uops_3_bits_csr_addr : _GEN_91 ? io_dis_uops_2_bits_csr_addr : _GEN_90 ? io_dis_uops_1_bits_csr_addr : io_dis_uops_0_bits_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_92 ? io_dis_uops_3_bits_rob_idx : _GEN_91 ? io_dis_uops_2_bits_rob_idx : _GEN_90 ? io_dis_uops_1_bits_rob_idx : io_dis_uops_0_bits_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_92 ? io_dis_uops_3_bits_ldq_idx : _GEN_91 ? io_dis_uops_2_bits_ldq_idx : _GEN_90 ? io_dis_uops_1_bits_ldq_idx : io_dis_uops_0_bits_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_92 ? io_dis_uops_3_bits_stq_idx : _GEN_91 ? io_dis_uops_2_bits_stq_idx : _GEN_90 ? io_dis_uops_1_bits_stq_idx : io_dis_uops_0_bits_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_92 ? io_dis_uops_3_bits_rxq_idx : _GEN_91 ? io_dis_uops_2_bits_rxq_idx : _GEN_90 ? io_dis_uops_1_bits_rxq_idx : io_dis_uops_0_bits_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_92 ? io_dis_uops_3_bits_pdst : _GEN_91 ? io_dis_uops_2_bits_pdst : _GEN_90 ? io_dis_uops_1_bits_pdst : io_dis_uops_0_bits_pdst),
    .io_in_uop_bits_prs1            (_GEN_92 ? io_dis_uops_3_bits_prs1 : _GEN_91 ? io_dis_uops_2_bits_prs1 : _GEN_90 ? io_dis_uops_1_bits_prs1 : io_dis_uops_0_bits_prs1),
    .io_in_uop_bits_prs2            (_GEN_92 ? io_dis_uops_3_bits_prs2 : _GEN_91 ? io_dis_uops_2_bits_prs2 : _GEN_90 ? io_dis_uops_1_bits_prs2 : io_dis_uops_0_bits_prs2),
    .io_in_uop_bits_prs3            (_GEN_92 ? io_dis_uops_3_bits_prs3 : _GEN_91 ? io_dis_uops_2_bits_prs3 : _GEN_90 ? io_dis_uops_1_bits_prs3 : io_dis_uops_0_bits_prs3),
    .io_in_uop_bits_ppred           (6'h0),
    .io_in_uop_bits_prs1_busy       (_GEN_92 ? io_dis_uops_3_bits_prs1_busy : _GEN_91 ? io_dis_uops_2_bits_prs1_busy : _GEN_90 ? io_dis_uops_1_bits_prs1_busy : io_dis_uops_0_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_92 ? _GEN_18 & io_dis_uops_3_bits_prs2_busy : _GEN_91 ? _GEN_15 : _GEN_90 ? _GEN_10 : _GEN_4),
    .io_in_uop_bits_prs3_busy       (1'h0),
    .io_in_uop_bits_ppred_busy      (1'h0),
    .io_in_uop_bits_stale_pdst      (_GEN_92 ? io_dis_uops_3_bits_stale_pdst : _GEN_91 ? io_dis_uops_2_bits_stale_pdst : _GEN_90 ? io_dis_uops_1_bits_stale_pdst : io_dis_uops_0_bits_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_92 ? io_dis_uops_3_bits_exception : _GEN_91 ? io_dis_uops_2_bits_exception : _GEN_90 ? io_dis_uops_1_bits_exception : io_dis_uops_0_bits_exception),
    .io_in_uop_bits_exc_cause       (_GEN_92 ? io_dis_uops_3_bits_exc_cause : _GEN_91 ? io_dis_uops_2_bits_exc_cause : _GEN_90 ? io_dis_uops_1_bits_exc_cause : io_dis_uops_0_bits_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_92 ? io_dis_uops_3_bits_bypassable : _GEN_91 ? io_dis_uops_2_bits_bypassable : _GEN_90 ? io_dis_uops_1_bits_bypassable : io_dis_uops_0_bits_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_92 ? io_dis_uops_3_bits_mem_cmd : _GEN_91 ? io_dis_uops_2_bits_mem_cmd : _GEN_90 ? io_dis_uops_1_bits_mem_cmd : io_dis_uops_0_bits_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_92 ? io_dis_uops_3_bits_mem_size : _GEN_91 ? io_dis_uops_2_bits_mem_size : _GEN_90 ? io_dis_uops_1_bits_mem_size : io_dis_uops_0_bits_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_92 ? io_dis_uops_3_bits_mem_signed : _GEN_91 ? io_dis_uops_2_bits_mem_signed : _GEN_90 ? io_dis_uops_1_bits_mem_signed : io_dis_uops_0_bits_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_92 ? io_dis_uops_3_bits_is_fence : _GEN_91 ? io_dis_uops_2_bits_is_fence : _GEN_90 ? io_dis_uops_1_bits_is_fence : io_dis_uops_0_bits_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_92 ? io_dis_uops_3_bits_is_fencei : _GEN_91 ? io_dis_uops_2_bits_is_fencei : _GEN_90 ? io_dis_uops_1_bits_is_fencei : io_dis_uops_0_bits_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_92 ? io_dis_uops_3_bits_is_amo : _GEN_91 ? io_dis_uops_2_bits_is_amo : _GEN_90 ? io_dis_uops_1_bits_is_amo : io_dis_uops_0_bits_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_92 ? io_dis_uops_3_bits_uses_ldq : _GEN_91 ? io_dis_uops_2_bits_uses_ldq : _GEN_90 ? io_dis_uops_1_bits_uses_ldq : io_dis_uops_0_bits_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_92 ? io_dis_uops_3_bits_uses_stq : _GEN_91 ? io_dis_uops_2_bits_uses_stq : _GEN_90 ? io_dis_uops_1_bits_uses_stq : io_dis_uops_0_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_92 ? io_dis_uops_3_bits_is_sys_pc2epc : _GEN_91 ? io_dis_uops_2_bits_is_sys_pc2epc : _GEN_90 ? io_dis_uops_1_bits_is_sys_pc2epc : io_dis_uops_0_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_92 ? io_dis_uops_3_bits_is_unique : _GEN_91 ? io_dis_uops_2_bits_is_unique : _GEN_90 ? io_dis_uops_1_bits_is_unique : io_dis_uops_0_bits_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_92 ? io_dis_uops_3_bits_flush_on_commit : _GEN_91 ? io_dis_uops_2_bits_flush_on_commit : _GEN_90 ? io_dis_uops_1_bits_flush_on_commit : io_dis_uops_0_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_92 ? io_dis_uops_3_bits_ldst_is_rs1 : _GEN_91 ? io_dis_uops_2_bits_ldst_is_rs1 : _GEN_90 ? io_dis_uops_1_bits_ldst_is_rs1 : io_dis_uops_0_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_92 ? io_dis_uops_3_bits_ldst : _GEN_91 ? io_dis_uops_2_bits_ldst : _GEN_90 ? io_dis_uops_1_bits_ldst : io_dis_uops_0_bits_ldst),
    .io_in_uop_bits_lrs1            (_GEN_92 ? io_dis_uops_3_bits_lrs1 : _GEN_91 ? io_dis_uops_2_bits_lrs1 : _GEN_90 ? io_dis_uops_1_bits_lrs1 : io_dis_uops_0_bits_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_92 ? io_dis_uops_3_bits_lrs2 : _GEN_91 ? io_dis_uops_2_bits_lrs2 : _GEN_90 ? io_dis_uops_1_bits_lrs2 : io_dis_uops_0_bits_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_92 ? io_dis_uops_3_bits_lrs3 : _GEN_91 ? io_dis_uops_2_bits_lrs3 : _GEN_90 ? io_dis_uops_1_bits_lrs3 : io_dis_uops_0_bits_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_92 ? io_dis_uops_3_bits_ldst_val : _GEN_91 ? io_dis_uops_2_bits_ldst_val : _GEN_90 ? io_dis_uops_1_bits_ldst_val : io_dis_uops_0_bits_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_92 ? io_dis_uops_3_bits_dst_rtype : _GEN_91 ? io_dis_uops_2_bits_dst_rtype : _GEN_90 ? io_dis_uops_1_bits_dst_rtype : io_dis_uops_0_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_92 ? io_dis_uops_3_bits_lrs1_rtype : _GEN_91 ? io_dis_uops_2_bits_lrs1_rtype : _GEN_90 ? io_dis_uops_1_bits_lrs1_rtype : io_dis_uops_0_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_92 ? (_GEN_18 ? io_dis_uops_3_bits_lrs2_rtype : 2'h2) : _GEN_91 ? _GEN_14 : _GEN_90 ? _GEN_9 : _GEN_3),
    .io_in_uop_bits_frs3_en         (_GEN_92 ? io_dis_uops_3_bits_frs3_en : _GEN_91 ? io_dis_uops_2_bits_frs3_en : _GEN_90 ? io_dis_uops_1_bits_frs3_en : io_dis_uops_0_bits_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_92 ? io_dis_uops_3_bits_fp_val : _GEN_91 ? io_dis_uops_2_bits_fp_val : _GEN_90 ? io_dis_uops_1_bits_fp_val : io_dis_uops_0_bits_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_92 ? io_dis_uops_3_bits_fp_single : _GEN_91 ? io_dis_uops_2_bits_fp_single : _GEN_90 ? io_dis_uops_1_bits_fp_single : io_dis_uops_0_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_92 ? io_dis_uops_3_bits_xcpt_pf_if : _GEN_91 ? io_dis_uops_2_bits_xcpt_pf_if : _GEN_90 ? io_dis_uops_1_bits_xcpt_pf_if : io_dis_uops_0_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_92 ? io_dis_uops_3_bits_xcpt_ae_if : _GEN_91 ? io_dis_uops_2_bits_xcpt_ae_if : _GEN_90 ? io_dis_uops_1_bits_xcpt_ae_if : io_dis_uops_0_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_92 ? io_dis_uops_3_bits_xcpt_ma_if : _GEN_91 ? io_dis_uops_2_bits_xcpt_ma_if : _GEN_90 ? io_dis_uops_1_bits_xcpt_ma_if : io_dis_uops_0_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_92 ? io_dis_uops_3_bits_bp_debug_if : _GEN_91 ? io_dis_uops_2_bits_bp_debug_if : _GEN_90 ? io_dis_uops_1_bits_bp_debug_if : io_dis_uops_0_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_92 ? io_dis_uops_3_bits_bp_xcpt_if : _GEN_91 ? io_dis_uops_2_bits_bp_xcpt_if : _GEN_90 ? io_dis_uops_1_bits_bp_xcpt_if : io_dis_uops_0_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_92 ? io_dis_uops_3_bits_debug_fsrc : _GEN_91 ? io_dis_uops_2_bits_debug_fsrc : _GEN_90 ? io_dis_uops_1_bits_debug_fsrc : io_dis_uops_0_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_92 ? io_dis_uops_3_bits_debug_tsrc : _GEN_91 ? io_dis_uops_2_bits_debug_tsrc : _GEN_90 ? io_dis_uops_1_bits_debug_tsrc : io_dis_uops_0_bits_debug_tsrc),
    .io_out_uop_uopc                (_slots_23_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_23_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_23_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_23_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_23_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_23_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_23_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_23_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_23_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_23_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_23_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_23_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_23_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_23_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_23_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_23_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_23_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_23_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_23_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_23_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_23_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_23_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_23_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_23_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_23_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_23_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_23_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_23_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_23_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_23_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_23_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_23_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_23_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_23_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_23_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_23_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_23_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_23_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_23_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_23_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_23_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_23_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_23_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_23_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_23_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_23_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_23_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_23_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_23_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_23_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_23_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_23_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_23_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_23_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_23_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_23_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_23_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_23_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_23_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_23_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_23_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_23_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_23_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_23_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_23_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_23_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_23_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_23_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_23_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_23_io_uop_uopc),
    .io_uop_inst                    (_slots_23_io_uop_inst),
    .io_uop_debug_inst              (_slots_23_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_23_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_23_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_23_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_23_io_uop_fu_code),
    .io_uop_iw_state                (_slots_23_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_23_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_23_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_23_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_23_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_23_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_23_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_23_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_23_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_23_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_23_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_23_io_uop_pc_lob),
    .io_uop_taken                   (_slots_23_io_uop_taken),
    .io_uop_imm_packed              (_slots_23_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_23_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_23_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_23_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_23_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_23_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_23_io_uop_pdst),
    .io_uop_prs1                    (_slots_23_io_uop_prs1),
    .io_uop_prs2                    (_slots_23_io_uop_prs2),
    .io_uop_prs3                    (_slots_23_io_uop_prs3),
    .io_uop_ppred                   (_slots_23_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_23_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_23_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_23_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_23_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_23_io_uop_stale_pdst),
    .io_uop_exception               (_slots_23_io_uop_exception),
    .io_uop_exc_cause               (_slots_23_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_23_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_23_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_23_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_23_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_23_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_23_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_23_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_23_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_23_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_23_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_23_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_23_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_23_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_23_io_uop_ldst),
    .io_uop_lrs1                    (_slots_23_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_23_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_23_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_23_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_23_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_23_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_23_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_23_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_23_io_uop_fp_val),
    .io_uop_fp_single               (_slots_23_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_23_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_23_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_23_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_23_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_23_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_23_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_23_io_uop_debug_tsrc)
  );
  assign io_dis_uops_0_ready = io_dis_uops_0_ready_REG;
  assign io_dis_uops_1_ready = io_dis_uops_1_ready_REG;
  assign io_dis_uops_2_ready = io_dis_uops_2_ready_REG;
  assign io_dis_uops_3_ready = io_dis_uops_3_ready_REG;
  assign io_iss_valids_0 = _GEN_225 | _GEN_222 | _GEN_216 | _GEN_210 | _GEN_204 | _GEN_198 | _GEN_192 | _GEN_186 | _GEN_180 | _GEN_174 | _GEN_168 | _GEN_162 | _GEN_156 | _GEN_150 | _GEN_144 | _GEN_138 | _GEN_132 | _GEN_126 | _GEN_120 | _GEN_114 | _GEN_108 | _GEN_102 | _GEN_96 | _GEN_93;
  assign io_iss_valids_1 = _GEN_226 | _GEN_224 | _GEN_219 | _GEN_213 | _GEN_207 | _GEN_201 | _GEN_195 | _GEN_189 | _GEN_183 | _GEN_177 | _GEN_171 | _GEN_165 | _GEN_159 | _GEN_153 | _GEN_147 | _GEN_141 | _GEN_135 | _GEN_129 | _GEN_123 | _GEN_117 | _GEN_111 | _GEN_105 | _GEN_99 | _GEN_94;
  assign io_iss_uops_0_uopc = _GEN_225 ? _slots_23_io_uop_uopc : _GEN_222 ? _slots_22_io_uop_uopc : _GEN_216 ? _slots_21_io_uop_uopc : _GEN_210 ? _slots_20_io_uop_uopc : _GEN_204 ? _slots_19_io_uop_uopc : _GEN_198 ? _slots_18_io_uop_uopc : _GEN_192 ? _slots_17_io_uop_uopc : _GEN_186 ? _slots_16_io_uop_uopc : _GEN_180 ? _slots_15_io_uop_uopc : _GEN_174 ? _slots_14_io_uop_uopc : _GEN_168 ? _slots_13_io_uop_uopc : _GEN_162 ? _slots_12_io_uop_uopc : _GEN_156 ? _slots_11_io_uop_uopc : _GEN_150 ? _slots_10_io_uop_uopc : _GEN_144 ? _slots_9_io_uop_uopc : _GEN_138 ? _slots_8_io_uop_uopc : _GEN_132 ? _slots_7_io_uop_uopc : _GEN_126 ? _slots_6_io_uop_uopc : _GEN_120 ? _slots_5_io_uop_uopc : _GEN_114 ? _slots_4_io_uop_uopc : _GEN_108 ? _slots_3_io_uop_uopc : _GEN_102 ? _slots_2_io_uop_uopc : _GEN_96 ? _slots_1_io_uop_uopc : _GEN_93 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_0_inst = _GEN_225 ? _slots_23_io_uop_inst : _GEN_222 ? _slots_22_io_uop_inst : _GEN_216 ? _slots_21_io_uop_inst : _GEN_210 ? _slots_20_io_uop_inst : _GEN_204 ? _slots_19_io_uop_inst : _GEN_198 ? _slots_18_io_uop_inst : _GEN_192 ? _slots_17_io_uop_inst : _GEN_186 ? _slots_16_io_uop_inst : _GEN_180 ? _slots_15_io_uop_inst : _GEN_174 ? _slots_14_io_uop_inst : _GEN_168 ? _slots_13_io_uop_inst : _GEN_162 ? _slots_12_io_uop_inst : _GEN_156 ? _slots_11_io_uop_inst : _GEN_150 ? _slots_10_io_uop_inst : _GEN_144 ? _slots_9_io_uop_inst : _GEN_138 ? _slots_8_io_uop_inst : _GEN_132 ? _slots_7_io_uop_inst : _GEN_126 ? _slots_6_io_uop_inst : _GEN_120 ? _slots_5_io_uop_inst : _GEN_114 ? _slots_4_io_uop_inst : _GEN_108 ? _slots_3_io_uop_inst : _GEN_102 ? _slots_2_io_uop_inst : _GEN_96 ? _slots_1_io_uop_inst : _GEN_93 ? _slots_0_io_uop_inst : 32'h0;
  assign io_iss_uops_0_debug_inst = _GEN_225 ? _slots_23_io_uop_debug_inst : _GEN_222 ? _slots_22_io_uop_debug_inst : _GEN_216 ? _slots_21_io_uop_debug_inst : _GEN_210 ? _slots_20_io_uop_debug_inst : _GEN_204 ? _slots_19_io_uop_debug_inst : _GEN_198 ? _slots_18_io_uop_debug_inst : _GEN_192 ? _slots_17_io_uop_debug_inst : _GEN_186 ? _slots_16_io_uop_debug_inst : _GEN_180 ? _slots_15_io_uop_debug_inst : _GEN_174 ? _slots_14_io_uop_debug_inst : _GEN_168 ? _slots_13_io_uop_debug_inst : _GEN_162 ? _slots_12_io_uop_debug_inst : _GEN_156 ? _slots_11_io_uop_debug_inst : _GEN_150 ? _slots_10_io_uop_debug_inst : _GEN_144 ? _slots_9_io_uop_debug_inst : _GEN_138 ? _slots_8_io_uop_debug_inst : _GEN_132 ? _slots_7_io_uop_debug_inst : _GEN_126 ? _slots_6_io_uop_debug_inst : _GEN_120 ? _slots_5_io_uop_debug_inst : _GEN_114 ? _slots_4_io_uop_debug_inst : _GEN_108 ? _slots_3_io_uop_debug_inst : _GEN_102 ? _slots_2_io_uop_debug_inst : _GEN_96 ? _slots_1_io_uop_debug_inst : _GEN_93 ? _slots_0_io_uop_debug_inst : 32'h0;
  assign io_iss_uops_0_is_rvc = _GEN_225 ? _slots_23_io_uop_is_rvc : _GEN_222 ? _slots_22_io_uop_is_rvc : _GEN_216 ? _slots_21_io_uop_is_rvc : _GEN_210 ? _slots_20_io_uop_is_rvc : _GEN_204 ? _slots_19_io_uop_is_rvc : _GEN_198 ? _slots_18_io_uop_is_rvc : _GEN_192 ? _slots_17_io_uop_is_rvc : _GEN_186 ? _slots_16_io_uop_is_rvc : _GEN_180 ? _slots_15_io_uop_is_rvc : _GEN_174 ? _slots_14_io_uop_is_rvc : _GEN_168 ? _slots_13_io_uop_is_rvc : _GEN_162 ? _slots_12_io_uop_is_rvc : _GEN_156 ? _slots_11_io_uop_is_rvc : _GEN_150 ? _slots_10_io_uop_is_rvc : _GEN_144 ? _slots_9_io_uop_is_rvc : _GEN_138 ? _slots_8_io_uop_is_rvc : _GEN_132 ? _slots_7_io_uop_is_rvc : _GEN_126 ? _slots_6_io_uop_is_rvc : _GEN_120 ? _slots_5_io_uop_is_rvc : _GEN_114 ? _slots_4_io_uop_is_rvc : _GEN_108 ? _slots_3_io_uop_is_rvc : _GEN_102 ? _slots_2_io_uop_is_rvc : _GEN_96 ? _slots_1_io_uop_is_rvc : _GEN_93 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_0_debug_pc = _GEN_225 ? _slots_23_io_uop_debug_pc : _GEN_222 ? _slots_22_io_uop_debug_pc : _GEN_216 ? _slots_21_io_uop_debug_pc : _GEN_210 ? _slots_20_io_uop_debug_pc : _GEN_204 ? _slots_19_io_uop_debug_pc : _GEN_198 ? _slots_18_io_uop_debug_pc : _GEN_192 ? _slots_17_io_uop_debug_pc : _GEN_186 ? _slots_16_io_uop_debug_pc : _GEN_180 ? _slots_15_io_uop_debug_pc : _GEN_174 ? _slots_14_io_uop_debug_pc : _GEN_168 ? _slots_13_io_uop_debug_pc : _GEN_162 ? _slots_12_io_uop_debug_pc : _GEN_156 ? _slots_11_io_uop_debug_pc : _GEN_150 ? _slots_10_io_uop_debug_pc : _GEN_144 ? _slots_9_io_uop_debug_pc : _GEN_138 ? _slots_8_io_uop_debug_pc : _GEN_132 ? _slots_7_io_uop_debug_pc : _GEN_126 ? _slots_6_io_uop_debug_pc : _GEN_120 ? _slots_5_io_uop_debug_pc : _GEN_114 ? _slots_4_io_uop_debug_pc : _GEN_108 ? _slots_3_io_uop_debug_pc : _GEN_102 ? _slots_2_io_uop_debug_pc : _GEN_96 ? _slots_1_io_uop_debug_pc : _GEN_93 ? _slots_0_io_uop_debug_pc : 40'h0;
  assign io_iss_uops_0_iq_type = _GEN_225 ? _slots_23_io_uop_iq_type : _GEN_222 ? _slots_22_io_uop_iq_type : _GEN_216 ? _slots_21_io_uop_iq_type : _GEN_210 ? _slots_20_io_uop_iq_type : _GEN_204 ? _slots_19_io_uop_iq_type : _GEN_198 ? _slots_18_io_uop_iq_type : _GEN_192 ? _slots_17_io_uop_iq_type : _GEN_186 ? _slots_16_io_uop_iq_type : _GEN_180 ? _slots_15_io_uop_iq_type : _GEN_174 ? _slots_14_io_uop_iq_type : _GEN_168 ? _slots_13_io_uop_iq_type : _GEN_162 ? _slots_12_io_uop_iq_type : _GEN_156 ? _slots_11_io_uop_iq_type : _GEN_150 ? _slots_10_io_uop_iq_type : _GEN_144 ? _slots_9_io_uop_iq_type : _GEN_138 ? _slots_8_io_uop_iq_type : _GEN_132 ? _slots_7_io_uop_iq_type : _GEN_126 ? _slots_6_io_uop_iq_type : _GEN_120 ? _slots_5_io_uop_iq_type : _GEN_114 ? _slots_4_io_uop_iq_type : _GEN_108 ? _slots_3_io_uop_iq_type : _GEN_102 ? _slots_2_io_uop_iq_type : _GEN_96 ? _slots_1_io_uop_iq_type : _GEN_93 ? _slots_0_io_uop_iq_type : 3'h0;
  assign io_iss_uops_0_fu_code = _GEN_225 ? _slots_23_io_uop_fu_code : _GEN_222 ? _slots_22_io_uop_fu_code : _GEN_216 ? _slots_21_io_uop_fu_code : _GEN_210 ? _slots_20_io_uop_fu_code : _GEN_204 ? _slots_19_io_uop_fu_code : _GEN_198 ? _slots_18_io_uop_fu_code : _GEN_192 ? _slots_17_io_uop_fu_code : _GEN_186 ? _slots_16_io_uop_fu_code : _GEN_180 ? _slots_15_io_uop_fu_code : _GEN_174 ? _slots_14_io_uop_fu_code : _GEN_168 ? _slots_13_io_uop_fu_code : _GEN_162 ? _slots_12_io_uop_fu_code : _GEN_156 ? _slots_11_io_uop_fu_code : _GEN_150 ? _slots_10_io_uop_fu_code : _GEN_144 ? _slots_9_io_uop_fu_code : _GEN_138 ? _slots_8_io_uop_fu_code : _GEN_132 ? _slots_7_io_uop_fu_code : _GEN_126 ? _slots_6_io_uop_fu_code : _GEN_120 ? _slots_5_io_uop_fu_code : _GEN_114 ? _slots_4_io_uop_fu_code : _GEN_108 ? _slots_3_io_uop_fu_code : _GEN_102 ? _slots_2_io_uop_fu_code : _GEN_96 ? _slots_1_io_uop_fu_code : _GEN_93 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_0_iw_state = _GEN_225 ? _slots_23_io_uop_iw_state : _GEN_222 ? _slots_22_io_uop_iw_state : _GEN_216 ? _slots_21_io_uop_iw_state : _GEN_210 ? _slots_20_io_uop_iw_state : _GEN_204 ? _slots_19_io_uop_iw_state : _GEN_198 ? _slots_18_io_uop_iw_state : _GEN_192 ? _slots_17_io_uop_iw_state : _GEN_186 ? _slots_16_io_uop_iw_state : _GEN_180 ? _slots_15_io_uop_iw_state : _GEN_174 ? _slots_14_io_uop_iw_state : _GEN_168 ? _slots_13_io_uop_iw_state : _GEN_162 ? _slots_12_io_uop_iw_state : _GEN_156 ? _slots_11_io_uop_iw_state : _GEN_150 ? _slots_10_io_uop_iw_state : _GEN_144 ? _slots_9_io_uop_iw_state : _GEN_138 ? _slots_8_io_uop_iw_state : _GEN_132 ? _slots_7_io_uop_iw_state : _GEN_126 ? _slots_6_io_uop_iw_state : _GEN_120 ? _slots_5_io_uop_iw_state : _GEN_114 ? _slots_4_io_uop_iw_state : _GEN_108 ? _slots_3_io_uop_iw_state : _GEN_102 ? _slots_2_io_uop_iw_state : _GEN_96 ? _slots_1_io_uop_iw_state : _GEN_93 ? _slots_0_io_uop_iw_state : 2'h0;
  assign io_iss_uops_0_iw_p1_poisoned = _GEN_225 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_222 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_216 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_210 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_204 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_198 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_192 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_186 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_180 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_174 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_168 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_162 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_156 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_150 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_144 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_138 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_132 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_126 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_120 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_114 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_108 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_102 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_96 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_93 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_0_iw_p2_poisoned = _GEN_225 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_222 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_216 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_210 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_204 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_198 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_192 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_186 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_180 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_174 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_168 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_162 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_156 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_150 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_144 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_138 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_132 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_126 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_120 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_114 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_108 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_102 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_96 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_93 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_0_is_br = _GEN_225 ? _slots_23_io_uop_is_br : _GEN_222 ? _slots_22_io_uop_is_br : _GEN_216 ? _slots_21_io_uop_is_br : _GEN_210 ? _slots_20_io_uop_is_br : _GEN_204 ? _slots_19_io_uop_is_br : _GEN_198 ? _slots_18_io_uop_is_br : _GEN_192 ? _slots_17_io_uop_is_br : _GEN_186 ? _slots_16_io_uop_is_br : _GEN_180 ? _slots_15_io_uop_is_br : _GEN_174 ? _slots_14_io_uop_is_br : _GEN_168 ? _slots_13_io_uop_is_br : _GEN_162 ? _slots_12_io_uop_is_br : _GEN_156 ? _slots_11_io_uop_is_br : _GEN_150 ? _slots_10_io_uop_is_br : _GEN_144 ? _slots_9_io_uop_is_br : _GEN_138 ? _slots_8_io_uop_is_br : _GEN_132 ? _slots_7_io_uop_is_br : _GEN_126 ? _slots_6_io_uop_is_br : _GEN_120 ? _slots_5_io_uop_is_br : _GEN_114 ? _slots_4_io_uop_is_br : _GEN_108 ? _slots_3_io_uop_is_br : _GEN_102 ? _slots_2_io_uop_is_br : _GEN_96 ? _slots_1_io_uop_is_br : _GEN_93 & _slots_0_io_uop_is_br;
  assign io_iss_uops_0_is_jalr = _GEN_225 ? _slots_23_io_uop_is_jalr : _GEN_222 ? _slots_22_io_uop_is_jalr : _GEN_216 ? _slots_21_io_uop_is_jalr : _GEN_210 ? _slots_20_io_uop_is_jalr : _GEN_204 ? _slots_19_io_uop_is_jalr : _GEN_198 ? _slots_18_io_uop_is_jalr : _GEN_192 ? _slots_17_io_uop_is_jalr : _GEN_186 ? _slots_16_io_uop_is_jalr : _GEN_180 ? _slots_15_io_uop_is_jalr : _GEN_174 ? _slots_14_io_uop_is_jalr : _GEN_168 ? _slots_13_io_uop_is_jalr : _GEN_162 ? _slots_12_io_uop_is_jalr : _GEN_156 ? _slots_11_io_uop_is_jalr : _GEN_150 ? _slots_10_io_uop_is_jalr : _GEN_144 ? _slots_9_io_uop_is_jalr : _GEN_138 ? _slots_8_io_uop_is_jalr : _GEN_132 ? _slots_7_io_uop_is_jalr : _GEN_126 ? _slots_6_io_uop_is_jalr : _GEN_120 ? _slots_5_io_uop_is_jalr : _GEN_114 ? _slots_4_io_uop_is_jalr : _GEN_108 ? _slots_3_io_uop_is_jalr : _GEN_102 ? _slots_2_io_uop_is_jalr : _GEN_96 ? _slots_1_io_uop_is_jalr : _GEN_93 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_0_is_jal = _GEN_225 ? _slots_23_io_uop_is_jal : _GEN_222 ? _slots_22_io_uop_is_jal : _GEN_216 ? _slots_21_io_uop_is_jal : _GEN_210 ? _slots_20_io_uop_is_jal : _GEN_204 ? _slots_19_io_uop_is_jal : _GEN_198 ? _slots_18_io_uop_is_jal : _GEN_192 ? _slots_17_io_uop_is_jal : _GEN_186 ? _slots_16_io_uop_is_jal : _GEN_180 ? _slots_15_io_uop_is_jal : _GEN_174 ? _slots_14_io_uop_is_jal : _GEN_168 ? _slots_13_io_uop_is_jal : _GEN_162 ? _slots_12_io_uop_is_jal : _GEN_156 ? _slots_11_io_uop_is_jal : _GEN_150 ? _slots_10_io_uop_is_jal : _GEN_144 ? _slots_9_io_uop_is_jal : _GEN_138 ? _slots_8_io_uop_is_jal : _GEN_132 ? _slots_7_io_uop_is_jal : _GEN_126 ? _slots_6_io_uop_is_jal : _GEN_120 ? _slots_5_io_uop_is_jal : _GEN_114 ? _slots_4_io_uop_is_jal : _GEN_108 ? _slots_3_io_uop_is_jal : _GEN_102 ? _slots_2_io_uop_is_jal : _GEN_96 ? _slots_1_io_uop_is_jal : _GEN_93 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_0_is_sfb = _GEN_225 ? _slots_23_io_uop_is_sfb : _GEN_222 ? _slots_22_io_uop_is_sfb : _GEN_216 ? _slots_21_io_uop_is_sfb : _GEN_210 ? _slots_20_io_uop_is_sfb : _GEN_204 ? _slots_19_io_uop_is_sfb : _GEN_198 ? _slots_18_io_uop_is_sfb : _GEN_192 ? _slots_17_io_uop_is_sfb : _GEN_186 ? _slots_16_io_uop_is_sfb : _GEN_180 ? _slots_15_io_uop_is_sfb : _GEN_174 ? _slots_14_io_uop_is_sfb : _GEN_168 ? _slots_13_io_uop_is_sfb : _GEN_162 ? _slots_12_io_uop_is_sfb : _GEN_156 ? _slots_11_io_uop_is_sfb : _GEN_150 ? _slots_10_io_uop_is_sfb : _GEN_144 ? _slots_9_io_uop_is_sfb : _GEN_138 ? _slots_8_io_uop_is_sfb : _GEN_132 ? _slots_7_io_uop_is_sfb : _GEN_126 ? _slots_6_io_uop_is_sfb : _GEN_120 ? _slots_5_io_uop_is_sfb : _GEN_114 ? _slots_4_io_uop_is_sfb : _GEN_108 ? _slots_3_io_uop_is_sfb : _GEN_102 ? _slots_2_io_uop_is_sfb : _GEN_96 ? _slots_1_io_uop_is_sfb : _GEN_93 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_0_br_mask = _GEN_225 ? _slots_23_io_uop_br_mask : _GEN_222 ? _slots_22_io_uop_br_mask : _GEN_216 ? _slots_21_io_uop_br_mask : _GEN_210 ? _slots_20_io_uop_br_mask : _GEN_204 ? _slots_19_io_uop_br_mask : _GEN_198 ? _slots_18_io_uop_br_mask : _GEN_192 ? _slots_17_io_uop_br_mask : _GEN_186 ? _slots_16_io_uop_br_mask : _GEN_180 ? _slots_15_io_uop_br_mask : _GEN_174 ? _slots_14_io_uop_br_mask : _GEN_168 ? _slots_13_io_uop_br_mask : _GEN_162 ? _slots_12_io_uop_br_mask : _GEN_156 ? _slots_11_io_uop_br_mask : _GEN_150 ? _slots_10_io_uop_br_mask : _GEN_144 ? _slots_9_io_uop_br_mask : _GEN_138 ? _slots_8_io_uop_br_mask : _GEN_132 ? _slots_7_io_uop_br_mask : _GEN_126 ? _slots_6_io_uop_br_mask : _GEN_120 ? _slots_5_io_uop_br_mask : _GEN_114 ? _slots_4_io_uop_br_mask : _GEN_108 ? _slots_3_io_uop_br_mask : _GEN_102 ? _slots_2_io_uop_br_mask : _GEN_96 ? _slots_1_io_uop_br_mask : _GEN_93 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_0_br_tag = _GEN_225 ? _slots_23_io_uop_br_tag : _GEN_222 ? _slots_22_io_uop_br_tag : _GEN_216 ? _slots_21_io_uop_br_tag : _GEN_210 ? _slots_20_io_uop_br_tag : _GEN_204 ? _slots_19_io_uop_br_tag : _GEN_198 ? _slots_18_io_uop_br_tag : _GEN_192 ? _slots_17_io_uop_br_tag : _GEN_186 ? _slots_16_io_uop_br_tag : _GEN_180 ? _slots_15_io_uop_br_tag : _GEN_174 ? _slots_14_io_uop_br_tag : _GEN_168 ? _slots_13_io_uop_br_tag : _GEN_162 ? _slots_12_io_uop_br_tag : _GEN_156 ? _slots_11_io_uop_br_tag : _GEN_150 ? _slots_10_io_uop_br_tag : _GEN_144 ? _slots_9_io_uop_br_tag : _GEN_138 ? _slots_8_io_uop_br_tag : _GEN_132 ? _slots_7_io_uop_br_tag : _GEN_126 ? _slots_6_io_uop_br_tag : _GEN_120 ? _slots_5_io_uop_br_tag : _GEN_114 ? _slots_4_io_uop_br_tag : _GEN_108 ? _slots_3_io_uop_br_tag : _GEN_102 ? _slots_2_io_uop_br_tag : _GEN_96 ? _slots_1_io_uop_br_tag : _GEN_93 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_0_ftq_idx = _GEN_225 ? _slots_23_io_uop_ftq_idx : _GEN_222 ? _slots_22_io_uop_ftq_idx : _GEN_216 ? _slots_21_io_uop_ftq_idx : _GEN_210 ? _slots_20_io_uop_ftq_idx : _GEN_204 ? _slots_19_io_uop_ftq_idx : _GEN_198 ? _slots_18_io_uop_ftq_idx : _GEN_192 ? _slots_17_io_uop_ftq_idx : _GEN_186 ? _slots_16_io_uop_ftq_idx : _GEN_180 ? _slots_15_io_uop_ftq_idx : _GEN_174 ? _slots_14_io_uop_ftq_idx : _GEN_168 ? _slots_13_io_uop_ftq_idx : _GEN_162 ? _slots_12_io_uop_ftq_idx : _GEN_156 ? _slots_11_io_uop_ftq_idx : _GEN_150 ? _slots_10_io_uop_ftq_idx : _GEN_144 ? _slots_9_io_uop_ftq_idx : _GEN_138 ? _slots_8_io_uop_ftq_idx : _GEN_132 ? _slots_7_io_uop_ftq_idx : _GEN_126 ? _slots_6_io_uop_ftq_idx : _GEN_120 ? _slots_5_io_uop_ftq_idx : _GEN_114 ? _slots_4_io_uop_ftq_idx : _GEN_108 ? _slots_3_io_uop_ftq_idx : _GEN_102 ? _slots_2_io_uop_ftq_idx : _GEN_96 ? _slots_1_io_uop_ftq_idx : _GEN_93 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_0_edge_inst = _GEN_225 ? _slots_23_io_uop_edge_inst : _GEN_222 ? _slots_22_io_uop_edge_inst : _GEN_216 ? _slots_21_io_uop_edge_inst : _GEN_210 ? _slots_20_io_uop_edge_inst : _GEN_204 ? _slots_19_io_uop_edge_inst : _GEN_198 ? _slots_18_io_uop_edge_inst : _GEN_192 ? _slots_17_io_uop_edge_inst : _GEN_186 ? _slots_16_io_uop_edge_inst : _GEN_180 ? _slots_15_io_uop_edge_inst : _GEN_174 ? _slots_14_io_uop_edge_inst : _GEN_168 ? _slots_13_io_uop_edge_inst : _GEN_162 ? _slots_12_io_uop_edge_inst : _GEN_156 ? _slots_11_io_uop_edge_inst : _GEN_150 ? _slots_10_io_uop_edge_inst : _GEN_144 ? _slots_9_io_uop_edge_inst : _GEN_138 ? _slots_8_io_uop_edge_inst : _GEN_132 ? _slots_7_io_uop_edge_inst : _GEN_126 ? _slots_6_io_uop_edge_inst : _GEN_120 ? _slots_5_io_uop_edge_inst : _GEN_114 ? _slots_4_io_uop_edge_inst : _GEN_108 ? _slots_3_io_uop_edge_inst : _GEN_102 ? _slots_2_io_uop_edge_inst : _GEN_96 ? _slots_1_io_uop_edge_inst : _GEN_93 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_0_pc_lob = _GEN_225 ? _slots_23_io_uop_pc_lob : _GEN_222 ? _slots_22_io_uop_pc_lob : _GEN_216 ? _slots_21_io_uop_pc_lob : _GEN_210 ? _slots_20_io_uop_pc_lob : _GEN_204 ? _slots_19_io_uop_pc_lob : _GEN_198 ? _slots_18_io_uop_pc_lob : _GEN_192 ? _slots_17_io_uop_pc_lob : _GEN_186 ? _slots_16_io_uop_pc_lob : _GEN_180 ? _slots_15_io_uop_pc_lob : _GEN_174 ? _slots_14_io_uop_pc_lob : _GEN_168 ? _slots_13_io_uop_pc_lob : _GEN_162 ? _slots_12_io_uop_pc_lob : _GEN_156 ? _slots_11_io_uop_pc_lob : _GEN_150 ? _slots_10_io_uop_pc_lob : _GEN_144 ? _slots_9_io_uop_pc_lob : _GEN_138 ? _slots_8_io_uop_pc_lob : _GEN_132 ? _slots_7_io_uop_pc_lob : _GEN_126 ? _slots_6_io_uop_pc_lob : _GEN_120 ? _slots_5_io_uop_pc_lob : _GEN_114 ? _slots_4_io_uop_pc_lob : _GEN_108 ? _slots_3_io_uop_pc_lob : _GEN_102 ? _slots_2_io_uop_pc_lob : _GEN_96 ? _slots_1_io_uop_pc_lob : _GEN_93 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_0_taken = _GEN_225 ? _slots_23_io_uop_taken : _GEN_222 ? _slots_22_io_uop_taken : _GEN_216 ? _slots_21_io_uop_taken : _GEN_210 ? _slots_20_io_uop_taken : _GEN_204 ? _slots_19_io_uop_taken : _GEN_198 ? _slots_18_io_uop_taken : _GEN_192 ? _slots_17_io_uop_taken : _GEN_186 ? _slots_16_io_uop_taken : _GEN_180 ? _slots_15_io_uop_taken : _GEN_174 ? _slots_14_io_uop_taken : _GEN_168 ? _slots_13_io_uop_taken : _GEN_162 ? _slots_12_io_uop_taken : _GEN_156 ? _slots_11_io_uop_taken : _GEN_150 ? _slots_10_io_uop_taken : _GEN_144 ? _slots_9_io_uop_taken : _GEN_138 ? _slots_8_io_uop_taken : _GEN_132 ? _slots_7_io_uop_taken : _GEN_126 ? _slots_6_io_uop_taken : _GEN_120 ? _slots_5_io_uop_taken : _GEN_114 ? _slots_4_io_uop_taken : _GEN_108 ? _slots_3_io_uop_taken : _GEN_102 ? _slots_2_io_uop_taken : _GEN_96 ? _slots_1_io_uop_taken : _GEN_93 & _slots_0_io_uop_taken;
  assign io_iss_uops_0_imm_packed = _GEN_225 ? _slots_23_io_uop_imm_packed : _GEN_222 ? _slots_22_io_uop_imm_packed : _GEN_216 ? _slots_21_io_uop_imm_packed : _GEN_210 ? _slots_20_io_uop_imm_packed : _GEN_204 ? _slots_19_io_uop_imm_packed : _GEN_198 ? _slots_18_io_uop_imm_packed : _GEN_192 ? _slots_17_io_uop_imm_packed : _GEN_186 ? _slots_16_io_uop_imm_packed : _GEN_180 ? _slots_15_io_uop_imm_packed : _GEN_174 ? _slots_14_io_uop_imm_packed : _GEN_168 ? _slots_13_io_uop_imm_packed : _GEN_162 ? _slots_12_io_uop_imm_packed : _GEN_156 ? _slots_11_io_uop_imm_packed : _GEN_150 ? _slots_10_io_uop_imm_packed : _GEN_144 ? _slots_9_io_uop_imm_packed : _GEN_138 ? _slots_8_io_uop_imm_packed : _GEN_132 ? _slots_7_io_uop_imm_packed : _GEN_126 ? _slots_6_io_uop_imm_packed : _GEN_120 ? _slots_5_io_uop_imm_packed : _GEN_114 ? _slots_4_io_uop_imm_packed : _GEN_108 ? _slots_3_io_uop_imm_packed : _GEN_102 ? _slots_2_io_uop_imm_packed : _GEN_96 ? _slots_1_io_uop_imm_packed : _GEN_93 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_0_csr_addr = _GEN_225 ? _slots_23_io_uop_csr_addr : _GEN_222 ? _slots_22_io_uop_csr_addr : _GEN_216 ? _slots_21_io_uop_csr_addr : _GEN_210 ? _slots_20_io_uop_csr_addr : _GEN_204 ? _slots_19_io_uop_csr_addr : _GEN_198 ? _slots_18_io_uop_csr_addr : _GEN_192 ? _slots_17_io_uop_csr_addr : _GEN_186 ? _slots_16_io_uop_csr_addr : _GEN_180 ? _slots_15_io_uop_csr_addr : _GEN_174 ? _slots_14_io_uop_csr_addr : _GEN_168 ? _slots_13_io_uop_csr_addr : _GEN_162 ? _slots_12_io_uop_csr_addr : _GEN_156 ? _slots_11_io_uop_csr_addr : _GEN_150 ? _slots_10_io_uop_csr_addr : _GEN_144 ? _slots_9_io_uop_csr_addr : _GEN_138 ? _slots_8_io_uop_csr_addr : _GEN_132 ? _slots_7_io_uop_csr_addr : _GEN_126 ? _slots_6_io_uop_csr_addr : _GEN_120 ? _slots_5_io_uop_csr_addr : _GEN_114 ? _slots_4_io_uop_csr_addr : _GEN_108 ? _slots_3_io_uop_csr_addr : _GEN_102 ? _slots_2_io_uop_csr_addr : _GEN_96 ? _slots_1_io_uop_csr_addr : _GEN_93 ? _slots_0_io_uop_csr_addr : 12'h0;
  assign io_iss_uops_0_rob_idx = _GEN_225 ? _slots_23_io_uop_rob_idx : _GEN_222 ? _slots_22_io_uop_rob_idx : _GEN_216 ? _slots_21_io_uop_rob_idx : _GEN_210 ? _slots_20_io_uop_rob_idx : _GEN_204 ? _slots_19_io_uop_rob_idx : _GEN_198 ? _slots_18_io_uop_rob_idx : _GEN_192 ? _slots_17_io_uop_rob_idx : _GEN_186 ? _slots_16_io_uop_rob_idx : _GEN_180 ? _slots_15_io_uop_rob_idx : _GEN_174 ? _slots_14_io_uop_rob_idx : _GEN_168 ? _slots_13_io_uop_rob_idx : _GEN_162 ? _slots_12_io_uop_rob_idx : _GEN_156 ? _slots_11_io_uop_rob_idx : _GEN_150 ? _slots_10_io_uop_rob_idx : _GEN_144 ? _slots_9_io_uop_rob_idx : _GEN_138 ? _slots_8_io_uop_rob_idx : _GEN_132 ? _slots_7_io_uop_rob_idx : _GEN_126 ? _slots_6_io_uop_rob_idx : _GEN_120 ? _slots_5_io_uop_rob_idx : _GEN_114 ? _slots_4_io_uop_rob_idx : _GEN_108 ? _slots_3_io_uop_rob_idx : _GEN_102 ? _slots_2_io_uop_rob_idx : _GEN_96 ? _slots_1_io_uop_rob_idx : _GEN_93 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_0_ldq_idx = _GEN_225 ? _slots_23_io_uop_ldq_idx : _GEN_222 ? _slots_22_io_uop_ldq_idx : _GEN_216 ? _slots_21_io_uop_ldq_idx : _GEN_210 ? _slots_20_io_uop_ldq_idx : _GEN_204 ? _slots_19_io_uop_ldq_idx : _GEN_198 ? _slots_18_io_uop_ldq_idx : _GEN_192 ? _slots_17_io_uop_ldq_idx : _GEN_186 ? _slots_16_io_uop_ldq_idx : _GEN_180 ? _slots_15_io_uop_ldq_idx : _GEN_174 ? _slots_14_io_uop_ldq_idx : _GEN_168 ? _slots_13_io_uop_ldq_idx : _GEN_162 ? _slots_12_io_uop_ldq_idx : _GEN_156 ? _slots_11_io_uop_ldq_idx : _GEN_150 ? _slots_10_io_uop_ldq_idx : _GEN_144 ? _slots_9_io_uop_ldq_idx : _GEN_138 ? _slots_8_io_uop_ldq_idx : _GEN_132 ? _slots_7_io_uop_ldq_idx : _GEN_126 ? _slots_6_io_uop_ldq_idx : _GEN_120 ? _slots_5_io_uop_ldq_idx : _GEN_114 ? _slots_4_io_uop_ldq_idx : _GEN_108 ? _slots_3_io_uop_ldq_idx : _GEN_102 ? _slots_2_io_uop_ldq_idx : _GEN_96 ? _slots_1_io_uop_ldq_idx : _GEN_93 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_0_stq_idx = _GEN_225 ? _slots_23_io_uop_stq_idx : _GEN_222 ? _slots_22_io_uop_stq_idx : _GEN_216 ? _slots_21_io_uop_stq_idx : _GEN_210 ? _slots_20_io_uop_stq_idx : _GEN_204 ? _slots_19_io_uop_stq_idx : _GEN_198 ? _slots_18_io_uop_stq_idx : _GEN_192 ? _slots_17_io_uop_stq_idx : _GEN_186 ? _slots_16_io_uop_stq_idx : _GEN_180 ? _slots_15_io_uop_stq_idx : _GEN_174 ? _slots_14_io_uop_stq_idx : _GEN_168 ? _slots_13_io_uop_stq_idx : _GEN_162 ? _slots_12_io_uop_stq_idx : _GEN_156 ? _slots_11_io_uop_stq_idx : _GEN_150 ? _slots_10_io_uop_stq_idx : _GEN_144 ? _slots_9_io_uop_stq_idx : _GEN_138 ? _slots_8_io_uop_stq_idx : _GEN_132 ? _slots_7_io_uop_stq_idx : _GEN_126 ? _slots_6_io_uop_stq_idx : _GEN_120 ? _slots_5_io_uop_stq_idx : _GEN_114 ? _slots_4_io_uop_stq_idx : _GEN_108 ? _slots_3_io_uop_stq_idx : _GEN_102 ? _slots_2_io_uop_stq_idx : _GEN_96 ? _slots_1_io_uop_stq_idx : _GEN_93 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_0_rxq_idx = _GEN_225 ? _slots_23_io_uop_rxq_idx : _GEN_222 ? _slots_22_io_uop_rxq_idx : _GEN_216 ? _slots_21_io_uop_rxq_idx : _GEN_210 ? _slots_20_io_uop_rxq_idx : _GEN_204 ? _slots_19_io_uop_rxq_idx : _GEN_198 ? _slots_18_io_uop_rxq_idx : _GEN_192 ? _slots_17_io_uop_rxq_idx : _GEN_186 ? _slots_16_io_uop_rxq_idx : _GEN_180 ? _slots_15_io_uop_rxq_idx : _GEN_174 ? _slots_14_io_uop_rxq_idx : _GEN_168 ? _slots_13_io_uop_rxq_idx : _GEN_162 ? _slots_12_io_uop_rxq_idx : _GEN_156 ? _slots_11_io_uop_rxq_idx : _GEN_150 ? _slots_10_io_uop_rxq_idx : _GEN_144 ? _slots_9_io_uop_rxq_idx : _GEN_138 ? _slots_8_io_uop_rxq_idx : _GEN_132 ? _slots_7_io_uop_rxq_idx : _GEN_126 ? _slots_6_io_uop_rxq_idx : _GEN_120 ? _slots_5_io_uop_rxq_idx : _GEN_114 ? _slots_4_io_uop_rxq_idx : _GEN_108 ? _slots_3_io_uop_rxq_idx : _GEN_102 ? _slots_2_io_uop_rxq_idx : _GEN_96 ? _slots_1_io_uop_rxq_idx : _GEN_93 ? _slots_0_io_uop_rxq_idx : 2'h0;
  assign io_iss_uops_0_pdst = _GEN_225 ? _slots_23_io_uop_pdst : _GEN_222 ? _slots_22_io_uop_pdst : _GEN_216 ? _slots_21_io_uop_pdst : _GEN_210 ? _slots_20_io_uop_pdst : _GEN_204 ? _slots_19_io_uop_pdst : _GEN_198 ? _slots_18_io_uop_pdst : _GEN_192 ? _slots_17_io_uop_pdst : _GEN_186 ? _slots_16_io_uop_pdst : _GEN_180 ? _slots_15_io_uop_pdst : _GEN_174 ? _slots_14_io_uop_pdst : _GEN_168 ? _slots_13_io_uop_pdst : _GEN_162 ? _slots_12_io_uop_pdst : _GEN_156 ? _slots_11_io_uop_pdst : _GEN_150 ? _slots_10_io_uop_pdst : _GEN_144 ? _slots_9_io_uop_pdst : _GEN_138 ? _slots_8_io_uop_pdst : _GEN_132 ? _slots_7_io_uop_pdst : _GEN_126 ? _slots_6_io_uop_pdst : _GEN_120 ? _slots_5_io_uop_pdst : _GEN_114 ? _slots_4_io_uop_pdst : _GEN_108 ? _slots_3_io_uop_pdst : _GEN_102 ? _slots_2_io_uop_pdst : _GEN_96 ? _slots_1_io_uop_pdst : _GEN_93 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_0_prs1 = _GEN_225 ? _slots_23_io_uop_prs1 : _GEN_222 ? _slots_22_io_uop_prs1 : _GEN_216 ? _slots_21_io_uop_prs1 : _GEN_210 ? _slots_20_io_uop_prs1 : _GEN_204 ? _slots_19_io_uop_prs1 : _GEN_198 ? _slots_18_io_uop_prs1 : _GEN_192 ? _slots_17_io_uop_prs1 : _GEN_186 ? _slots_16_io_uop_prs1 : _GEN_180 ? _slots_15_io_uop_prs1 : _GEN_174 ? _slots_14_io_uop_prs1 : _GEN_168 ? _slots_13_io_uop_prs1 : _GEN_162 ? _slots_12_io_uop_prs1 : _GEN_156 ? _slots_11_io_uop_prs1 : _GEN_150 ? _slots_10_io_uop_prs1 : _GEN_144 ? _slots_9_io_uop_prs1 : _GEN_138 ? _slots_8_io_uop_prs1 : _GEN_132 ? _slots_7_io_uop_prs1 : _GEN_126 ? _slots_6_io_uop_prs1 : _GEN_120 ? _slots_5_io_uop_prs1 : _GEN_114 ? _slots_4_io_uop_prs1 : _GEN_108 ? _slots_3_io_uop_prs1 : _GEN_102 ? _slots_2_io_uop_prs1 : _GEN_96 ? _slots_1_io_uop_prs1 : _GEN_93 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_0_prs2 = _GEN_225 ? _slots_23_io_uop_prs2 : _GEN_222 ? _slots_22_io_uop_prs2 : _GEN_216 ? _slots_21_io_uop_prs2 : _GEN_210 ? _slots_20_io_uop_prs2 : _GEN_204 ? _slots_19_io_uop_prs2 : _GEN_198 ? _slots_18_io_uop_prs2 : _GEN_192 ? _slots_17_io_uop_prs2 : _GEN_186 ? _slots_16_io_uop_prs2 : _GEN_180 ? _slots_15_io_uop_prs2 : _GEN_174 ? _slots_14_io_uop_prs2 : _GEN_168 ? _slots_13_io_uop_prs2 : _GEN_162 ? _slots_12_io_uop_prs2 : _GEN_156 ? _slots_11_io_uop_prs2 : _GEN_150 ? _slots_10_io_uop_prs2 : _GEN_144 ? _slots_9_io_uop_prs2 : _GEN_138 ? _slots_8_io_uop_prs2 : _GEN_132 ? _slots_7_io_uop_prs2 : _GEN_126 ? _slots_6_io_uop_prs2 : _GEN_120 ? _slots_5_io_uop_prs2 : _GEN_114 ? _slots_4_io_uop_prs2 : _GEN_108 ? _slots_3_io_uop_prs2 : _GEN_102 ? _slots_2_io_uop_prs2 : _GEN_96 ? _slots_1_io_uop_prs2 : _GEN_93 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_0_prs3 = _GEN_225 ? _slots_23_io_uop_prs3 : _GEN_222 ? _slots_22_io_uop_prs3 : _GEN_216 ? _slots_21_io_uop_prs3 : _GEN_210 ? _slots_20_io_uop_prs3 : _GEN_204 ? _slots_19_io_uop_prs3 : _GEN_198 ? _slots_18_io_uop_prs3 : _GEN_192 ? _slots_17_io_uop_prs3 : _GEN_186 ? _slots_16_io_uop_prs3 : _GEN_180 ? _slots_15_io_uop_prs3 : _GEN_174 ? _slots_14_io_uop_prs3 : _GEN_168 ? _slots_13_io_uop_prs3 : _GEN_162 ? _slots_12_io_uop_prs3 : _GEN_156 ? _slots_11_io_uop_prs3 : _GEN_150 ? _slots_10_io_uop_prs3 : _GEN_144 ? _slots_9_io_uop_prs3 : _GEN_138 ? _slots_8_io_uop_prs3 : _GEN_132 ? _slots_7_io_uop_prs3 : _GEN_126 ? _slots_6_io_uop_prs3 : _GEN_120 ? _slots_5_io_uop_prs3 : _GEN_114 ? _slots_4_io_uop_prs3 : _GEN_108 ? _slots_3_io_uop_prs3 : _GEN_102 ? _slots_2_io_uop_prs3 : _GEN_96 ? _slots_1_io_uop_prs3 : _GEN_93 ? _slots_0_io_uop_prs3 : 7'h0;
  assign io_iss_uops_0_ppred = _GEN_225 ? _slots_23_io_uop_ppred : _GEN_222 ? _slots_22_io_uop_ppred : _GEN_216 ? _slots_21_io_uop_ppred : _GEN_210 ? _slots_20_io_uop_ppred : _GEN_204 ? _slots_19_io_uop_ppred : _GEN_198 ? _slots_18_io_uop_ppred : _GEN_192 ? _slots_17_io_uop_ppred : _GEN_186 ? _slots_16_io_uop_ppred : _GEN_180 ? _slots_15_io_uop_ppred : _GEN_174 ? _slots_14_io_uop_ppred : _GEN_168 ? _slots_13_io_uop_ppred : _GEN_162 ? _slots_12_io_uop_ppred : _GEN_156 ? _slots_11_io_uop_ppred : _GEN_150 ? _slots_10_io_uop_ppred : _GEN_144 ? _slots_9_io_uop_ppred : _GEN_138 ? _slots_8_io_uop_ppred : _GEN_132 ? _slots_7_io_uop_ppred : _GEN_126 ? _slots_6_io_uop_ppred : _GEN_120 ? _slots_5_io_uop_ppred : _GEN_114 ? _slots_4_io_uop_ppred : _GEN_108 ? _slots_3_io_uop_ppred : _GEN_102 ? _slots_2_io_uop_ppred : _GEN_96 ? _slots_1_io_uop_ppred : _GEN_93 ? _slots_0_io_uop_ppred : 6'h0;
  assign io_iss_uops_0_prs1_busy = _GEN_225 ? _slots_23_io_uop_prs1_busy : _GEN_222 ? _slots_22_io_uop_prs1_busy : _GEN_216 ? _slots_21_io_uop_prs1_busy : _GEN_210 ? _slots_20_io_uop_prs1_busy : _GEN_204 ? _slots_19_io_uop_prs1_busy : _GEN_198 ? _slots_18_io_uop_prs1_busy : _GEN_192 ? _slots_17_io_uop_prs1_busy : _GEN_186 ? _slots_16_io_uop_prs1_busy : _GEN_180 ? _slots_15_io_uop_prs1_busy : _GEN_174 ? _slots_14_io_uop_prs1_busy : _GEN_168 ? _slots_13_io_uop_prs1_busy : _GEN_162 ? _slots_12_io_uop_prs1_busy : _GEN_156 ? _slots_11_io_uop_prs1_busy : _GEN_150 ? _slots_10_io_uop_prs1_busy : _GEN_144 ? _slots_9_io_uop_prs1_busy : _GEN_138 ? _slots_8_io_uop_prs1_busy : _GEN_132 ? _slots_7_io_uop_prs1_busy : _GEN_126 ? _slots_6_io_uop_prs1_busy : _GEN_120 ? _slots_5_io_uop_prs1_busy : _GEN_114 ? _slots_4_io_uop_prs1_busy : _GEN_108 ? _slots_3_io_uop_prs1_busy : _GEN_102 ? _slots_2_io_uop_prs1_busy : _GEN_96 ? _slots_1_io_uop_prs1_busy : _GEN_93 & _slots_0_io_uop_prs1_busy;
  assign io_iss_uops_0_prs2_busy = _GEN_225 ? _slots_23_io_uop_prs2_busy : _GEN_222 ? _slots_22_io_uop_prs2_busy : _GEN_216 ? _slots_21_io_uop_prs2_busy : _GEN_210 ? _slots_20_io_uop_prs2_busy : _GEN_204 ? _slots_19_io_uop_prs2_busy : _GEN_198 ? _slots_18_io_uop_prs2_busy : _GEN_192 ? _slots_17_io_uop_prs2_busy : _GEN_186 ? _slots_16_io_uop_prs2_busy : _GEN_180 ? _slots_15_io_uop_prs2_busy : _GEN_174 ? _slots_14_io_uop_prs2_busy : _GEN_168 ? _slots_13_io_uop_prs2_busy : _GEN_162 ? _slots_12_io_uop_prs2_busy : _GEN_156 ? _slots_11_io_uop_prs2_busy : _GEN_150 ? _slots_10_io_uop_prs2_busy : _GEN_144 ? _slots_9_io_uop_prs2_busy : _GEN_138 ? _slots_8_io_uop_prs2_busy : _GEN_132 ? _slots_7_io_uop_prs2_busy : _GEN_126 ? _slots_6_io_uop_prs2_busy : _GEN_120 ? _slots_5_io_uop_prs2_busy : _GEN_114 ? _slots_4_io_uop_prs2_busy : _GEN_108 ? _slots_3_io_uop_prs2_busy : _GEN_102 ? _slots_2_io_uop_prs2_busy : _GEN_96 ? _slots_1_io_uop_prs2_busy : _GEN_93 & _slots_0_io_uop_prs2_busy;
  assign io_iss_uops_0_prs3_busy = _GEN_225 ? _slots_23_io_uop_prs3_busy : _GEN_222 ? _slots_22_io_uop_prs3_busy : _GEN_216 ? _slots_21_io_uop_prs3_busy : _GEN_210 ? _slots_20_io_uop_prs3_busy : _GEN_204 ? _slots_19_io_uop_prs3_busy : _GEN_198 ? _slots_18_io_uop_prs3_busy : _GEN_192 ? _slots_17_io_uop_prs3_busy : _GEN_186 ? _slots_16_io_uop_prs3_busy : _GEN_180 ? _slots_15_io_uop_prs3_busy : _GEN_174 ? _slots_14_io_uop_prs3_busy : _GEN_168 ? _slots_13_io_uop_prs3_busy : _GEN_162 ? _slots_12_io_uop_prs3_busy : _GEN_156 ? _slots_11_io_uop_prs3_busy : _GEN_150 ? _slots_10_io_uop_prs3_busy : _GEN_144 ? _slots_9_io_uop_prs3_busy : _GEN_138 ? _slots_8_io_uop_prs3_busy : _GEN_132 ? _slots_7_io_uop_prs3_busy : _GEN_126 ? _slots_6_io_uop_prs3_busy : _GEN_120 ? _slots_5_io_uop_prs3_busy : _GEN_114 ? _slots_4_io_uop_prs3_busy : _GEN_108 ? _slots_3_io_uop_prs3_busy : _GEN_102 ? _slots_2_io_uop_prs3_busy : _GEN_96 ? _slots_1_io_uop_prs3_busy : _GEN_93 & _slots_0_io_uop_prs3_busy;
  assign io_iss_uops_0_ppred_busy = _GEN_225 ? _slots_23_io_uop_ppred_busy : _GEN_222 ? _slots_22_io_uop_ppred_busy : _GEN_216 ? _slots_21_io_uop_ppred_busy : _GEN_210 ? _slots_20_io_uop_ppred_busy : _GEN_204 ? _slots_19_io_uop_ppred_busy : _GEN_198 ? _slots_18_io_uop_ppred_busy : _GEN_192 ? _slots_17_io_uop_ppred_busy : _GEN_186 ? _slots_16_io_uop_ppred_busy : _GEN_180 ? _slots_15_io_uop_ppred_busy : _GEN_174 ? _slots_14_io_uop_ppred_busy : _GEN_168 ? _slots_13_io_uop_ppred_busy : _GEN_162 ? _slots_12_io_uop_ppred_busy : _GEN_156 ? _slots_11_io_uop_ppred_busy : _GEN_150 ? _slots_10_io_uop_ppred_busy : _GEN_144 ? _slots_9_io_uop_ppred_busy : _GEN_138 ? _slots_8_io_uop_ppred_busy : _GEN_132 ? _slots_7_io_uop_ppred_busy : _GEN_126 ? _slots_6_io_uop_ppred_busy : _GEN_120 ? _slots_5_io_uop_ppred_busy : _GEN_114 ? _slots_4_io_uop_ppred_busy : _GEN_108 ? _slots_3_io_uop_ppred_busy : _GEN_102 ? _slots_2_io_uop_ppred_busy : _GEN_96 ? _slots_1_io_uop_ppred_busy : _GEN_93 & _slots_0_io_uop_ppred_busy;
  assign io_iss_uops_0_stale_pdst = _GEN_225 ? _slots_23_io_uop_stale_pdst : _GEN_222 ? _slots_22_io_uop_stale_pdst : _GEN_216 ? _slots_21_io_uop_stale_pdst : _GEN_210 ? _slots_20_io_uop_stale_pdst : _GEN_204 ? _slots_19_io_uop_stale_pdst : _GEN_198 ? _slots_18_io_uop_stale_pdst : _GEN_192 ? _slots_17_io_uop_stale_pdst : _GEN_186 ? _slots_16_io_uop_stale_pdst : _GEN_180 ? _slots_15_io_uop_stale_pdst : _GEN_174 ? _slots_14_io_uop_stale_pdst : _GEN_168 ? _slots_13_io_uop_stale_pdst : _GEN_162 ? _slots_12_io_uop_stale_pdst : _GEN_156 ? _slots_11_io_uop_stale_pdst : _GEN_150 ? _slots_10_io_uop_stale_pdst : _GEN_144 ? _slots_9_io_uop_stale_pdst : _GEN_138 ? _slots_8_io_uop_stale_pdst : _GEN_132 ? _slots_7_io_uop_stale_pdst : _GEN_126 ? _slots_6_io_uop_stale_pdst : _GEN_120 ? _slots_5_io_uop_stale_pdst : _GEN_114 ? _slots_4_io_uop_stale_pdst : _GEN_108 ? _slots_3_io_uop_stale_pdst : _GEN_102 ? _slots_2_io_uop_stale_pdst : _GEN_96 ? _slots_1_io_uop_stale_pdst : _GEN_93 ? _slots_0_io_uop_stale_pdst : 7'h0;
  assign io_iss_uops_0_exception = _GEN_225 ? _slots_23_io_uop_exception : _GEN_222 ? _slots_22_io_uop_exception : _GEN_216 ? _slots_21_io_uop_exception : _GEN_210 ? _slots_20_io_uop_exception : _GEN_204 ? _slots_19_io_uop_exception : _GEN_198 ? _slots_18_io_uop_exception : _GEN_192 ? _slots_17_io_uop_exception : _GEN_186 ? _slots_16_io_uop_exception : _GEN_180 ? _slots_15_io_uop_exception : _GEN_174 ? _slots_14_io_uop_exception : _GEN_168 ? _slots_13_io_uop_exception : _GEN_162 ? _slots_12_io_uop_exception : _GEN_156 ? _slots_11_io_uop_exception : _GEN_150 ? _slots_10_io_uop_exception : _GEN_144 ? _slots_9_io_uop_exception : _GEN_138 ? _slots_8_io_uop_exception : _GEN_132 ? _slots_7_io_uop_exception : _GEN_126 ? _slots_6_io_uop_exception : _GEN_120 ? _slots_5_io_uop_exception : _GEN_114 ? _slots_4_io_uop_exception : _GEN_108 ? _slots_3_io_uop_exception : _GEN_102 ? _slots_2_io_uop_exception : _GEN_96 ? _slots_1_io_uop_exception : _GEN_93 & _slots_0_io_uop_exception;
  assign io_iss_uops_0_exc_cause = _GEN_225 ? _slots_23_io_uop_exc_cause : _GEN_222 ? _slots_22_io_uop_exc_cause : _GEN_216 ? _slots_21_io_uop_exc_cause : _GEN_210 ? _slots_20_io_uop_exc_cause : _GEN_204 ? _slots_19_io_uop_exc_cause : _GEN_198 ? _slots_18_io_uop_exc_cause : _GEN_192 ? _slots_17_io_uop_exc_cause : _GEN_186 ? _slots_16_io_uop_exc_cause : _GEN_180 ? _slots_15_io_uop_exc_cause : _GEN_174 ? _slots_14_io_uop_exc_cause : _GEN_168 ? _slots_13_io_uop_exc_cause : _GEN_162 ? _slots_12_io_uop_exc_cause : _GEN_156 ? _slots_11_io_uop_exc_cause : _GEN_150 ? _slots_10_io_uop_exc_cause : _GEN_144 ? _slots_9_io_uop_exc_cause : _GEN_138 ? _slots_8_io_uop_exc_cause : _GEN_132 ? _slots_7_io_uop_exc_cause : _GEN_126 ? _slots_6_io_uop_exc_cause : _GEN_120 ? _slots_5_io_uop_exc_cause : _GEN_114 ? _slots_4_io_uop_exc_cause : _GEN_108 ? _slots_3_io_uop_exc_cause : _GEN_102 ? _slots_2_io_uop_exc_cause : _GEN_96 ? _slots_1_io_uop_exc_cause : _GEN_93 ? _slots_0_io_uop_exc_cause : 64'h0;
  assign io_iss_uops_0_bypassable = _GEN_225 ? _slots_23_io_uop_bypassable : _GEN_222 ? _slots_22_io_uop_bypassable : _GEN_216 ? _slots_21_io_uop_bypassable : _GEN_210 ? _slots_20_io_uop_bypassable : _GEN_204 ? _slots_19_io_uop_bypassable : _GEN_198 ? _slots_18_io_uop_bypassable : _GEN_192 ? _slots_17_io_uop_bypassable : _GEN_186 ? _slots_16_io_uop_bypassable : _GEN_180 ? _slots_15_io_uop_bypassable : _GEN_174 ? _slots_14_io_uop_bypassable : _GEN_168 ? _slots_13_io_uop_bypassable : _GEN_162 ? _slots_12_io_uop_bypassable : _GEN_156 ? _slots_11_io_uop_bypassable : _GEN_150 ? _slots_10_io_uop_bypassable : _GEN_144 ? _slots_9_io_uop_bypassable : _GEN_138 ? _slots_8_io_uop_bypassable : _GEN_132 ? _slots_7_io_uop_bypassable : _GEN_126 ? _slots_6_io_uop_bypassable : _GEN_120 ? _slots_5_io_uop_bypassable : _GEN_114 ? _slots_4_io_uop_bypassable : _GEN_108 ? _slots_3_io_uop_bypassable : _GEN_102 ? _slots_2_io_uop_bypassable : _GEN_96 ? _slots_1_io_uop_bypassable : _GEN_93 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_0_mem_cmd = _GEN_225 ? _slots_23_io_uop_mem_cmd : _GEN_222 ? _slots_22_io_uop_mem_cmd : _GEN_216 ? _slots_21_io_uop_mem_cmd : _GEN_210 ? _slots_20_io_uop_mem_cmd : _GEN_204 ? _slots_19_io_uop_mem_cmd : _GEN_198 ? _slots_18_io_uop_mem_cmd : _GEN_192 ? _slots_17_io_uop_mem_cmd : _GEN_186 ? _slots_16_io_uop_mem_cmd : _GEN_180 ? _slots_15_io_uop_mem_cmd : _GEN_174 ? _slots_14_io_uop_mem_cmd : _GEN_168 ? _slots_13_io_uop_mem_cmd : _GEN_162 ? _slots_12_io_uop_mem_cmd : _GEN_156 ? _slots_11_io_uop_mem_cmd : _GEN_150 ? _slots_10_io_uop_mem_cmd : _GEN_144 ? _slots_9_io_uop_mem_cmd : _GEN_138 ? _slots_8_io_uop_mem_cmd : _GEN_132 ? _slots_7_io_uop_mem_cmd : _GEN_126 ? _slots_6_io_uop_mem_cmd : _GEN_120 ? _slots_5_io_uop_mem_cmd : _GEN_114 ? _slots_4_io_uop_mem_cmd : _GEN_108 ? _slots_3_io_uop_mem_cmd : _GEN_102 ? _slots_2_io_uop_mem_cmd : _GEN_96 ? _slots_1_io_uop_mem_cmd : _GEN_93 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_0_mem_size = _GEN_225 ? _slots_23_io_uop_mem_size : _GEN_222 ? _slots_22_io_uop_mem_size : _GEN_216 ? _slots_21_io_uop_mem_size : _GEN_210 ? _slots_20_io_uop_mem_size : _GEN_204 ? _slots_19_io_uop_mem_size : _GEN_198 ? _slots_18_io_uop_mem_size : _GEN_192 ? _slots_17_io_uop_mem_size : _GEN_186 ? _slots_16_io_uop_mem_size : _GEN_180 ? _slots_15_io_uop_mem_size : _GEN_174 ? _slots_14_io_uop_mem_size : _GEN_168 ? _slots_13_io_uop_mem_size : _GEN_162 ? _slots_12_io_uop_mem_size : _GEN_156 ? _slots_11_io_uop_mem_size : _GEN_150 ? _slots_10_io_uop_mem_size : _GEN_144 ? _slots_9_io_uop_mem_size : _GEN_138 ? _slots_8_io_uop_mem_size : _GEN_132 ? _slots_7_io_uop_mem_size : _GEN_126 ? _slots_6_io_uop_mem_size : _GEN_120 ? _slots_5_io_uop_mem_size : _GEN_114 ? _slots_4_io_uop_mem_size : _GEN_108 ? _slots_3_io_uop_mem_size : _GEN_102 ? _slots_2_io_uop_mem_size : _GEN_96 ? _slots_1_io_uop_mem_size : _GEN_93 ? _slots_0_io_uop_mem_size : 2'h0;
  assign io_iss_uops_0_mem_signed = _GEN_225 ? _slots_23_io_uop_mem_signed : _GEN_222 ? _slots_22_io_uop_mem_signed : _GEN_216 ? _slots_21_io_uop_mem_signed : _GEN_210 ? _slots_20_io_uop_mem_signed : _GEN_204 ? _slots_19_io_uop_mem_signed : _GEN_198 ? _slots_18_io_uop_mem_signed : _GEN_192 ? _slots_17_io_uop_mem_signed : _GEN_186 ? _slots_16_io_uop_mem_signed : _GEN_180 ? _slots_15_io_uop_mem_signed : _GEN_174 ? _slots_14_io_uop_mem_signed : _GEN_168 ? _slots_13_io_uop_mem_signed : _GEN_162 ? _slots_12_io_uop_mem_signed : _GEN_156 ? _slots_11_io_uop_mem_signed : _GEN_150 ? _slots_10_io_uop_mem_signed : _GEN_144 ? _slots_9_io_uop_mem_signed : _GEN_138 ? _slots_8_io_uop_mem_signed : _GEN_132 ? _slots_7_io_uop_mem_signed : _GEN_126 ? _slots_6_io_uop_mem_signed : _GEN_120 ? _slots_5_io_uop_mem_signed : _GEN_114 ? _slots_4_io_uop_mem_signed : _GEN_108 ? _slots_3_io_uop_mem_signed : _GEN_102 ? _slots_2_io_uop_mem_signed : _GEN_96 ? _slots_1_io_uop_mem_signed : _GEN_93 & _slots_0_io_uop_mem_signed;
  assign io_iss_uops_0_is_fence = _GEN_225 ? _slots_23_io_uop_is_fence : _GEN_222 ? _slots_22_io_uop_is_fence : _GEN_216 ? _slots_21_io_uop_is_fence : _GEN_210 ? _slots_20_io_uop_is_fence : _GEN_204 ? _slots_19_io_uop_is_fence : _GEN_198 ? _slots_18_io_uop_is_fence : _GEN_192 ? _slots_17_io_uop_is_fence : _GEN_186 ? _slots_16_io_uop_is_fence : _GEN_180 ? _slots_15_io_uop_is_fence : _GEN_174 ? _slots_14_io_uop_is_fence : _GEN_168 ? _slots_13_io_uop_is_fence : _GEN_162 ? _slots_12_io_uop_is_fence : _GEN_156 ? _slots_11_io_uop_is_fence : _GEN_150 ? _slots_10_io_uop_is_fence : _GEN_144 ? _slots_9_io_uop_is_fence : _GEN_138 ? _slots_8_io_uop_is_fence : _GEN_132 ? _slots_7_io_uop_is_fence : _GEN_126 ? _slots_6_io_uop_is_fence : _GEN_120 ? _slots_5_io_uop_is_fence : _GEN_114 ? _slots_4_io_uop_is_fence : _GEN_108 ? _slots_3_io_uop_is_fence : _GEN_102 ? _slots_2_io_uop_is_fence : _GEN_96 ? _slots_1_io_uop_is_fence : _GEN_93 & _slots_0_io_uop_is_fence;
  assign io_iss_uops_0_is_fencei = _GEN_225 ? _slots_23_io_uop_is_fencei : _GEN_222 ? _slots_22_io_uop_is_fencei : _GEN_216 ? _slots_21_io_uop_is_fencei : _GEN_210 ? _slots_20_io_uop_is_fencei : _GEN_204 ? _slots_19_io_uop_is_fencei : _GEN_198 ? _slots_18_io_uop_is_fencei : _GEN_192 ? _slots_17_io_uop_is_fencei : _GEN_186 ? _slots_16_io_uop_is_fencei : _GEN_180 ? _slots_15_io_uop_is_fencei : _GEN_174 ? _slots_14_io_uop_is_fencei : _GEN_168 ? _slots_13_io_uop_is_fencei : _GEN_162 ? _slots_12_io_uop_is_fencei : _GEN_156 ? _slots_11_io_uop_is_fencei : _GEN_150 ? _slots_10_io_uop_is_fencei : _GEN_144 ? _slots_9_io_uop_is_fencei : _GEN_138 ? _slots_8_io_uop_is_fencei : _GEN_132 ? _slots_7_io_uop_is_fencei : _GEN_126 ? _slots_6_io_uop_is_fencei : _GEN_120 ? _slots_5_io_uop_is_fencei : _GEN_114 ? _slots_4_io_uop_is_fencei : _GEN_108 ? _slots_3_io_uop_is_fencei : _GEN_102 ? _slots_2_io_uop_is_fencei : _GEN_96 ? _slots_1_io_uop_is_fencei : _GEN_93 & _slots_0_io_uop_is_fencei;
  assign io_iss_uops_0_is_amo = _GEN_225 ? _slots_23_io_uop_is_amo : _GEN_222 ? _slots_22_io_uop_is_amo : _GEN_216 ? _slots_21_io_uop_is_amo : _GEN_210 ? _slots_20_io_uop_is_amo : _GEN_204 ? _slots_19_io_uop_is_amo : _GEN_198 ? _slots_18_io_uop_is_amo : _GEN_192 ? _slots_17_io_uop_is_amo : _GEN_186 ? _slots_16_io_uop_is_amo : _GEN_180 ? _slots_15_io_uop_is_amo : _GEN_174 ? _slots_14_io_uop_is_amo : _GEN_168 ? _slots_13_io_uop_is_amo : _GEN_162 ? _slots_12_io_uop_is_amo : _GEN_156 ? _slots_11_io_uop_is_amo : _GEN_150 ? _slots_10_io_uop_is_amo : _GEN_144 ? _slots_9_io_uop_is_amo : _GEN_138 ? _slots_8_io_uop_is_amo : _GEN_132 ? _slots_7_io_uop_is_amo : _GEN_126 ? _slots_6_io_uop_is_amo : _GEN_120 ? _slots_5_io_uop_is_amo : _GEN_114 ? _slots_4_io_uop_is_amo : _GEN_108 ? _slots_3_io_uop_is_amo : _GEN_102 ? _slots_2_io_uop_is_amo : _GEN_96 ? _slots_1_io_uop_is_amo : _GEN_93 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_0_uses_ldq = _GEN_225 ? _slots_23_io_uop_uses_ldq : _GEN_222 ? _slots_22_io_uop_uses_ldq : _GEN_216 ? _slots_21_io_uop_uses_ldq : _GEN_210 ? _slots_20_io_uop_uses_ldq : _GEN_204 ? _slots_19_io_uop_uses_ldq : _GEN_198 ? _slots_18_io_uop_uses_ldq : _GEN_192 ? _slots_17_io_uop_uses_ldq : _GEN_186 ? _slots_16_io_uop_uses_ldq : _GEN_180 ? _slots_15_io_uop_uses_ldq : _GEN_174 ? _slots_14_io_uop_uses_ldq : _GEN_168 ? _slots_13_io_uop_uses_ldq : _GEN_162 ? _slots_12_io_uop_uses_ldq : _GEN_156 ? _slots_11_io_uop_uses_ldq : _GEN_150 ? _slots_10_io_uop_uses_ldq : _GEN_144 ? _slots_9_io_uop_uses_ldq : _GEN_138 ? _slots_8_io_uop_uses_ldq : _GEN_132 ? _slots_7_io_uop_uses_ldq : _GEN_126 ? _slots_6_io_uop_uses_ldq : _GEN_120 ? _slots_5_io_uop_uses_ldq : _GEN_114 ? _slots_4_io_uop_uses_ldq : _GEN_108 ? _slots_3_io_uop_uses_ldq : _GEN_102 ? _slots_2_io_uop_uses_ldq : _GEN_96 ? _slots_1_io_uop_uses_ldq : _GEN_93 & _slots_0_io_uop_uses_ldq;
  assign io_iss_uops_0_uses_stq = _GEN_225 ? _slots_23_io_uop_uses_stq : _GEN_222 ? _slots_22_io_uop_uses_stq : _GEN_216 ? _slots_21_io_uop_uses_stq : _GEN_210 ? _slots_20_io_uop_uses_stq : _GEN_204 ? _slots_19_io_uop_uses_stq : _GEN_198 ? _slots_18_io_uop_uses_stq : _GEN_192 ? _slots_17_io_uop_uses_stq : _GEN_186 ? _slots_16_io_uop_uses_stq : _GEN_180 ? _slots_15_io_uop_uses_stq : _GEN_174 ? _slots_14_io_uop_uses_stq : _GEN_168 ? _slots_13_io_uop_uses_stq : _GEN_162 ? _slots_12_io_uop_uses_stq : _GEN_156 ? _slots_11_io_uop_uses_stq : _GEN_150 ? _slots_10_io_uop_uses_stq : _GEN_144 ? _slots_9_io_uop_uses_stq : _GEN_138 ? _slots_8_io_uop_uses_stq : _GEN_132 ? _slots_7_io_uop_uses_stq : _GEN_126 ? _slots_6_io_uop_uses_stq : _GEN_120 ? _slots_5_io_uop_uses_stq : _GEN_114 ? _slots_4_io_uop_uses_stq : _GEN_108 ? _slots_3_io_uop_uses_stq : _GEN_102 ? _slots_2_io_uop_uses_stq : _GEN_96 ? _slots_1_io_uop_uses_stq : _GEN_93 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_0_is_sys_pc2epc = _GEN_225 ? _slots_23_io_uop_is_sys_pc2epc : _GEN_222 ? _slots_22_io_uop_is_sys_pc2epc : _GEN_216 ? _slots_21_io_uop_is_sys_pc2epc : _GEN_210 ? _slots_20_io_uop_is_sys_pc2epc : _GEN_204 ? _slots_19_io_uop_is_sys_pc2epc : _GEN_198 ? _slots_18_io_uop_is_sys_pc2epc : _GEN_192 ? _slots_17_io_uop_is_sys_pc2epc : _GEN_186 ? _slots_16_io_uop_is_sys_pc2epc : _GEN_180 ? _slots_15_io_uop_is_sys_pc2epc : _GEN_174 ? _slots_14_io_uop_is_sys_pc2epc : _GEN_168 ? _slots_13_io_uop_is_sys_pc2epc : _GEN_162 ? _slots_12_io_uop_is_sys_pc2epc : _GEN_156 ? _slots_11_io_uop_is_sys_pc2epc : _GEN_150 ? _slots_10_io_uop_is_sys_pc2epc : _GEN_144 ? _slots_9_io_uop_is_sys_pc2epc : _GEN_138 ? _slots_8_io_uop_is_sys_pc2epc : _GEN_132 ? _slots_7_io_uop_is_sys_pc2epc : _GEN_126 ? _slots_6_io_uop_is_sys_pc2epc : _GEN_120 ? _slots_5_io_uop_is_sys_pc2epc : _GEN_114 ? _slots_4_io_uop_is_sys_pc2epc : _GEN_108 ? _slots_3_io_uop_is_sys_pc2epc : _GEN_102 ? _slots_2_io_uop_is_sys_pc2epc : _GEN_96 ? _slots_1_io_uop_is_sys_pc2epc : _GEN_93 & _slots_0_io_uop_is_sys_pc2epc;
  assign io_iss_uops_0_is_unique = _GEN_225 ? _slots_23_io_uop_is_unique : _GEN_222 ? _slots_22_io_uop_is_unique : _GEN_216 ? _slots_21_io_uop_is_unique : _GEN_210 ? _slots_20_io_uop_is_unique : _GEN_204 ? _slots_19_io_uop_is_unique : _GEN_198 ? _slots_18_io_uop_is_unique : _GEN_192 ? _slots_17_io_uop_is_unique : _GEN_186 ? _slots_16_io_uop_is_unique : _GEN_180 ? _slots_15_io_uop_is_unique : _GEN_174 ? _slots_14_io_uop_is_unique : _GEN_168 ? _slots_13_io_uop_is_unique : _GEN_162 ? _slots_12_io_uop_is_unique : _GEN_156 ? _slots_11_io_uop_is_unique : _GEN_150 ? _slots_10_io_uop_is_unique : _GEN_144 ? _slots_9_io_uop_is_unique : _GEN_138 ? _slots_8_io_uop_is_unique : _GEN_132 ? _slots_7_io_uop_is_unique : _GEN_126 ? _slots_6_io_uop_is_unique : _GEN_120 ? _slots_5_io_uop_is_unique : _GEN_114 ? _slots_4_io_uop_is_unique : _GEN_108 ? _slots_3_io_uop_is_unique : _GEN_102 ? _slots_2_io_uop_is_unique : _GEN_96 ? _slots_1_io_uop_is_unique : _GEN_93 & _slots_0_io_uop_is_unique;
  assign io_iss_uops_0_flush_on_commit = _GEN_225 ? _slots_23_io_uop_flush_on_commit : _GEN_222 ? _slots_22_io_uop_flush_on_commit : _GEN_216 ? _slots_21_io_uop_flush_on_commit : _GEN_210 ? _slots_20_io_uop_flush_on_commit : _GEN_204 ? _slots_19_io_uop_flush_on_commit : _GEN_198 ? _slots_18_io_uop_flush_on_commit : _GEN_192 ? _slots_17_io_uop_flush_on_commit : _GEN_186 ? _slots_16_io_uop_flush_on_commit : _GEN_180 ? _slots_15_io_uop_flush_on_commit : _GEN_174 ? _slots_14_io_uop_flush_on_commit : _GEN_168 ? _slots_13_io_uop_flush_on_commit : _GEN_162 ? _slots_12_io_uop_flush_on_commit : _GEN_156 ? _slots_11_io_uop_flush_on_commit : _GEN_150 ? _slots_10_io_uop_flush_on_commit : _GEN_144 ? _slots_9_io_uop_flush_on_commit : _GEN_138 ? _slots_8_io_uop_flush_on_commit : _GEN_132 ? _slots_7_io_uop_flush_on_commit : _GEN_126 ? _slots_6_io_uop_flush_on_commit : _GEN_120 ? _slots_5_io_uop_flush_on_commit : _GEN_114 ? _slots_4_io_uop_flush_on_commit : _GEN_108 ? _slots_3_io_uop_flush_on_commit : _GEN_102 ? _slots_2_io_uop_flush_on_commit : _GEN_96 ? _slots_1_io_uop_flush_on_commit : _GEN_93 & _slots_0_io_uop_flush_on_commit;
  assign io_iss_uops_0_ldst_is_rs1 = _GEN_225 ? _slots_23_io_uop_ldst_is_rs1 : _GEN_222 ? _slots_22_io_uop_ldst_is_rs1 : _GEN_216 ? _slots_21_io_uop_ldst_is_rs1 : _GEN_210 ? _slots_20_io_uop_ldst_is_rs1 : _GEN_204 ? _slots_19_io_uop_ldst_is_rs1 : _GEN_198 ? _slots_18_io_uop_ldst_is_rs1 : _GEN_192 ? _slots_17_io_uop_ldst_is_rs1 : _GEN_186 ? _slots_16_io_uop_ldst_is_rs1 : _GEN_180 ? _slots_15_io_uop_ldst_is_rs1 : _GEN_174 ? _slots_14_io_uop_ldst_is_rs1 : _GEN_168 ? _slots_13_io_uop_ldst_is_rs1 : _GEN_162 ? _slots_12_io_uop_ldst_is_rs1 : _GEN_156 ? _slots_11_io_uop_ldst_is_rs1 : _GEN_150 ? _slots_10_io_uop_ldst_is_rs1 : _GEN_144 ? _slots_9_io_uop_ldst_is_rs1 : _GEN_138 ? _slots_8_io_uop_ldst_is_rs1 : _GEN_132 ? _slots_7_io_uop_ldst_is_rs1 : _GEN_126 ? _slots_6_io_uop_ldst_is_rs1 : _GEN_120 ? _slots_5_io_uop_ldst_is_rs1 : _GEN_114 ? _slots_4_io_uop_ldst_is_rs1 : _GEN_108 ? _slots_3_io_uop_ldst_is_rs1 : _GEN_102 ? _slots_2_io_uop_ldst_is_rs1 : _GEN_96 ? _slots_1_io_uop_ldst_is_rs1 : _GEN_93 & _slots_0_io_uop_ldst_is_rs1;
  assign io_iss_uops_0_ldst = _GEN_225 ? _slots_23_io_uop_ldst : _GEN_222 ? _slots_22_io_uop_ldst : _GEN_216 ? _slots_21_io_uop_ldst : _GEN_210 ? _slots_20_io_uop_ldst : _GEN_204 ? _slots_19_io_uop_ldst : _GEN_198 ? _slots_18_io_uop_ldst : _GEN_192 ? _slots_17_io_uop_ldst : _GEN_186 ? _slots_16_io_uop_ldst : _GEN_180 ? _slots_15_io_uop_ldst : _GEN_174 ? _slots_14_io_uop_ldst : _GEN_168 ? _slots_13_io_uop_ldst : _GEN_162 ? _slots_12_io_uop_ldst : _GEN_156 ? _slots_11_io_uop_ldst : _GEN_150 ? _slots_10_io_uop_ldst : _GEN_144 ? _slots_9_io_uop_ldst : _GEN_138 ? _slots_8_io_uop_ldst : _GEN_132 ? _slots_7_io_uop_ldst : _GEN_126 ? _slots_6_io_uop_ldst : _GEN_120 ? _slots_5_io_uop_ldst : _GEN_114 ? _slots_4_io_uop_ldst : _GEN_108 ? _slots_3_io_uop_ldst : _GEN_102 ? _slots_2_io_uop_ldst : _GEN_96 ? _slots_1_io_uop_ldst : _GEN_93 ? _slots_0_io_uop_ldst : 6'h0;
  assign io_iss_uops_0_lrs1 = _GEN_225 ? _slots_23_io_uop_lrs1 : _GEN_222 ? _slots_22_io_uop_lrs1 : _GEN_216 ? _slots_21_io_uop_lrs1 : _GEN_210 ? _slots_20_io_uop_lrs1 : _GEN_204 ? _slots_19_io_uop_lrs1 : _GEN_198 ? _slots_18_io_uop_lrs1 : _GEN_192 ? _slots_17_io_uop_lrs1 : _GEN_186 ? _slots_16_io_uop_lrs1 : _GEN_180 ? _slots_15_io_uop_lrs1 : _GEN_174 ? _slots_14_io_uop_lrs1 : _GEN_168 ? _slots_13_io_uop_lrs1 : _GEN_162 ? _slots_12_io_uop_lrs1 : _GEN_156 ? _slots_11_io_uop_lrs1 : _GEN_150 ? _slots_10_io_uop_lrs1 : _GEN_144 ? _slots_9_io_uop_lrs1 : _GEN_138 ? _slots_8_io_uop_lrs1 : _GEN_132 ? _slots_7_io_uop_lrs1 : _GEN_126 ? _slots_6_io_uop_lrs1 : _GEN_120 ? _slots_5_io_uop_lrs1 : _GEN_114 ? _slots_4_io_uop_lrs1 : _GEN_108 ? _slots_3_io_uop_lrs1 : _GEN_102 ? _slots_2_io_uop_lrs1 : _GEN_96 ? _slots_1_io_uop_lrs1 : _GEN_93 ? _slots_0_io_uop_lrs1 : 6'h0;
  assign io_iss_uops_0_lrs2 = _GEN_225 ? _slots_23_io_uop_lrs2 : _GEN_222 ? _slots_22_io_uop_lrs2 : _GEN_216 ? _slots_21_io_uop_lrs2 : _GEN_210 ? _slots_20_io_uop_lrs2 : _GEN_204 ? _slots_19_io_uop_lrs2 : _GEN_198 ? _slots_18_io_uop_lrs2 : _GEN_192 ? _slots_17_io_uop_lrs2 : _GEN_186 ? _slots_16_io_uop_lrs2 : _GEN_180 ? _slots_15_io_uop_lrs2 : _GEN_174 ? _slots_14_io_uop_lrs2 : _GEN_168 ? _slots_13_io_uop_lrs2 : _GEN_162 ? _slots_12_io_uop_lrs2 : _GEN_156 ? _slots_11_io_uop_lrs2 : _GEN_150 ? _slots_10_io_uop_lrs2 : _GEN_144 ? _slots_9_io_uop_lrs2 : _GEN_138 ? _slots_8_io_uop_lrs2 : _GEN_132 ? _slots_7_io_uop_lrs2 : _GEN_126 ? _slots_6_io_uop_lrs2 : _GEN_120 ? _slots_5_io_uop_lrs2 : _GEN_114 ? _slots_4_io_uop_lrs2 : _GEN_108 ? _slots_3_io_uop_lrs2 : _GEN_102 ? _slots_2_io_uop_lrs2 : _GEN_96 ? _slots_1_io_uop_lrs2 : _GEN_93 ? _slots_0_io_uop_lrs2 : 6'h0;
  assign io_iss_uops_0_lrs3 = _GEN_225 ? _slots_23_io_uop_lrs3 : _GEN_222 ? _slots_22_io_uop_lrs3 : _GEN_216 ? _slots_21_io_uop_lrs3 : _GEN_210 ? _slots_20_io_uop_lrs3 : _GEN_204 ? _slots_19_io_uop_lrs3 : _GEN_198 ? _slots_18_io_uop_lrs3 : _GEN_192 ? _slots_17_io_uop_lrs3 : _GEN_186 ? _slots_16_io_uop_lrs3 : _GEN_180 ? _slots_15_io_uop_lrs3 : _GEN_174 ? _slots_14_io_uop_lrs3 : _GEN_168 ? _slots_13_io_uop_lrs3 : _GEN_162 ? _slots_12_io_uop_lrs3 : _GEN_156 ? _slots_11_io_uop_lrs3 : _GEN_150 ? _slots_10_io_uop_lrs3 : _GEN_144 ? _slots_9_io_uop_lrs3 : _GEN_138 ? _slots_8_io_uop_lrs3 : _GEN_132 ? _slots_7_io_uop_lrs3 : _GEN_126 ? _slots_6_io_uop_lrs3 : _GEN_120 ? _slots_5_io_uop_lrs3 : _GEN_114 ? _slots_4_io_uop_lrs3 : _GEN_108 ? _slots_3_io_uop_lrs3 : _GEN_102 ? _slots_2_io_uop_lrs3 : _GEN_96 ? _slots_1_io_uop_lrs3 : _GEN_93 ? _slots_0_io_uop_lrs3 : 6'h0;
  assign io_iss_uops_0_ldst_val = _GEN_225 ? _slots_23_io_uop_ldst_val : _GEN_222 ? _slots_22_io_uop_ldst_val : _GEN_216 ? _slots_21_io_uop_ldst_val : _GEN_210 ? _slots_20_io_uop_ldst_val : _GEN_204 ? _slots_19_io_uop_ldst_val : _GEN_198 ? _slots_18_io_uop_ldst_val : _GEN_192 ? _slots_17_io_uop_ldst_val : _GEN_186 ? _slots_16_io_uop_ldst_val : _GEN_180 ? _slots_15_io_uop_ldst_val : _GEN_174 ? _slots_14_io_uop_ldst_val : _GEN_168 ? _slots_13_io_uop_ldst_val : _GEN_162 ? _slots_12_io_uop_ldst_val : _GEN_156 ? _slots_11_io_uop_ldst_val : _GEN_150 ? _slots_10_io_uop_ldst_val : _GEN_144 ? _slots_9_io_uop_ldst_val : _GEN_138 ? _slots_8_io_uop_ldst_val : _GEN_132 ? _slots_7_io_uop_ldst_val : _GEN_126 ? _slots_6_io_uop_ldst_val : _GEN_120 ? _slots_5_io_uop_ldst_val : _GEN_114 ? _slots_4_io_uop_ldst_val : _GEN_108 ? _slots_3_io_uop_ldst_val : _GEN_102 ? _slots_2_io_uop_ldst_val : _GEN_96 ? _slots_1_io_uop_ldst_val : _GEN_93 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_0_dst_rtype = _GEN_225 ? _slots_23_io_uop_dst_rtype : _GEN_222 ? _slots_22_io_uop_dst_rtype : _GEN_216 ? _slots_21_io_uop_dst_rtype : _GEN_210 ? _slots_20_io_uop_dst_rtype : _GEN_204 ? _slots_19_io_uop_dst_rtype : _GEN_198 ? _slots_18_io_uop_dst_rtype : _GEN_192 ? _slots_17_io_uop_dst_rtype : _GEN_186 ? _slots_16_io_uop_dst_rtype : _GEN_180 ? _slots_15_io_uop_dst_rtype : _GEN_174 ? _slots_14_io_uop_dst_rtype : _GEN_168 ? _slots_13_io_uop_dst_rtype : _GEN_162 ? _slots_12_io_uop_dst_rtype : _GEN_156 ? _slots_11_io_uop_dst_rtype : _GEN_150 ? _slots_10_io_uop_dst_rtype : _GEN_144 ? _slots_9_io_uop_dst_rtype : _GEN_138 ? _slots_8_io_uop_dst_rtype : _GEN_132 ? _slots_7_io_uop_dst_rtype : _GEN_126 ? _slots_6_io_uop_dst_rtype : _GEN_120 ? _slots_5_io_uop_dst_rtype : _GEN_114 ? _slots_4_io_uop_dst_rtype : _GEN_108 ? _slots_3_io_uop_dst_rtype : _GEN_102 ? _slots_2_io_uop_dst_rtype : _GEN_96 ? _slots_1_io_uop_dst_rtype : _GEN_93 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_0_lrs1_rtype = _GEN_225 ? _slots_23_io_uop_lrs1_rtype : _GEN_222 ? _slots_22_io_uop_lrs1_rtype : _GEN_216 ? _slots_21_io_uop_lrs1_rtype : _GEN_210 ? _slots_20_io_uop_lrs1_rtype : _GEN_204 ? _slots_19_io_uop_lrs1_rtype : _GEN_198 ? _slots_18_io_uop_lrs1_rtype : _GEN_192 ? _slots_17_io_uop_lrs1_rtype : _GEN_186 ? _slots_16_io_uop_lrs1_rtype : _GEN_180 ? _slots_15_io_uop_lrs1_rtype : _GEN_174 ? _slots_14_io_uop_lrs1_rtype : _GEN_168 ? _slots_13_io_uop_lrs1_rtype : _GEN_162 ? _slots_12_io_uop_lrs1_rtype : _GEN_156 ? _slots_11_io_uop_lrs1_rtype : _GEN_150 ? _slots_10_io_uop_lrs1_rtype : _GEN_144 ? _slots_9_io_uop_lrs1_rtype : _GEN_138 ? _slots_8_io_uop_lrs1_rtype : _GEN_132 ? _slots_7_io_uop_lrs1_rtype : _GEN_126 ? _slots_6_io_uop_lrs1_rtype : _GEN_120 ? _slots_5_io_uop_lrs1_rtype : _GEN_114 ? _slots_4_io_uop_lrs1_rtype : _GEN_108 ? _slots_3_io_uop_lrs1_rtype : _GEN_102 ? _slots_2_io_uop_lrs1_rtype : _GEN_96 ? _slots_1_io_uop_lrs1_rtype : _GEN_93 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_0_lrs2_rtype = _GEN_225 ? _slots_23_io_uop_lrs2_rtype : _GEN_222 ? _slots_22_io_uop_lrs2_rtype : _GEN_216 ? _slots_21_io_uop_lrs2_rtype : _GEN_210 ? _slots_20_io_uop_lrs2_rtype : _GEN_204 ? _slots_19_io_uop_lrs2_rtype : _GEN_198 ? _slots_18_io_uop_lrs2_rtype : _GEN_192 ? _slots_17_io_uop_lrs2_rtype : _GEN_186 ? _slots_16_io_uop_lrs2_rtype : _GEN_180 ? _slots_15_io_uop_lrs2_rtype : _GEN_174 ? _slots_14_io_uop_lrs2_rtype : _GEN_168 ? _slots_13_io_uop_lrs2_rtype : _GEN_162 ? _slots_12_io_uop_lrs2_rtype : _GEN_156 ? _slots_11_io_uop_lrs2_rtype : _GEN_150 ? _slots_10_io_uop_lrs2_rtype : _GEN_144 ? _slots_9_io_uop_lrs2_rtype : _GEN_138 ? _slots_8_io_uop_lrs2_rtype : _GEN_132 ? _slots_7_io_uop_lrs2_rtype : _GEN_126 ? _slots_6_io_uop_lrs2_rtype : _GEN_120 ? _slots_5_io_uop_lrs2_rtype : _GEN_114 ? _slots_4_io_uop_lrs2_rtype : _GEN_108 ? _slots_3_io_uop_lrs2_rtype : _GEN_102 ? _slots_2_io_uop_lrs2_rtype : _GEN_96 ? _slots_1_io_uop_lrs2_rtype : _GEN_93 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_0_frs3_en = _GEN_225 ? _slots_23_io_uop_frs3_en : _GEN_222 ? _slots_22_io_uop_frs3_en : _GEN_216 ? _slots_21_io_uop_frs3_en : _GEN_210 ? _slots_20_io_uop_frs3_en : _GEN_204 ? _slots_19_io_uop_frs3_en : _GEN_198 ? _slots_18_io_uop_frs3_en : _GEN_192 ? _slots_17_io_uop_frs3_en : _GEN_186 ? _slots_16_io_uop_frs3_en : _GEN_180 ? _slots_15_io_uop_frs3_en : _GEN_174 ? _slots_14_io_uop_frs3_en : _GEN_168 ? _slots_13_io_uop_frs3_en : _GEN_162 ? _slots_12_io_uop_frs3_en : _GEN_156 ? _slots_11_io_uop_frs3_en : _GEN_150 ? _slots_10_io_uop_frs3_en : _GEN_144 ? _slots_9_io_uop_frs3_en : _GEN_138 ? _slots_8_io_uop_frs3_en : _GEN_132 ? _slots_7_io_uop_frs3_en : _GEN_126 ? _slots_6_io_uop_frs3_en : _GEN_120 ? _slots_5_io_uop_frs3_en : _GEN_114 ? _slots_4_io_uop_frs3_en : _GEN_108 ? _slots_3_io_uop_frs3_en : _GEN_102 ? _slots_2_io_uop_frs3_en : _GEN_96 ? _slots_1_io_uop_frs3_en : _GEN_93 & _slots_0_io_uop_frs3_en;
  assign io_iss_uops_0_fp_val = _GEN_225 ? _slots_23_io_uop_fp_val : _GEN_222 ? _slots_22_io_uop_fp_val : _GEN_216 ? _slots_21_io_uop_fp_val : _GEN_210 ? _slots_20_io_uop_fp_val : _GEN_204 ? _slots_19_io_uop_fp_val : _GEN_198 ? _slots_18_io_uop_fp_val : _GEN_192 ? _slots_17_io_uop_fp_val : _GEN_186 ? _slots_16_io_uop_fp_val : _GEN_180 ? _slots_15_io_uop_fp_val : _GEN_174 ? _slots_14_io_uop_fp_val : _GEN_168 ? _slots_13_io_uop_fp_val : _GEN_162 ? _slots_12_io_uop_fp_val : _GEN_156 ? _slots_11_io_uop_fp_val : _GEN_150 ? _slots_10_io_uop_fp_val : _GEN_144 ? _slots_9_io_uop_fp_val : _GEN_138 ? _slots_8_io_uop_fp_val : _GEN_132 ? _slots_7_io_uop_fp_val : _GEN_126 ? _slots_6_io_uop_fp_val : _GEN_120 ? _slots_5_io_uop_fp_val : _GEN_114 ? _slots_4_io_uop_fp_val : _GEN_108 ? _slots_3_io_uop_fp_val : _GEN_102 ? _slots_2_io_uop_fp_val : _GEN_96 ? _slots_1_io_uop_fp_val : _GEN_93 & _slots_0_io_uop_fp_val;
  assign io_iss_uops_0_fp_single = _GEN_225 ? _slots_23_io_uop_fp_single : _GEN_222 ? _slots_22_io_uop_fp_single : _GEN_216 ? _slots_21_io_uop_fp_single : _GEN_210 ? _slots_20_io_uop_fp_single : _GEN_204 ? _slots_19_io_uop_fp_single : _GEN_198 ? _slots_18_io_uop_fp_single : _GEN_192 ? _slots_17_io_uop_fp_single : _GEN_186 ? _slots_16_io_uop_fp_single : _GEN_180 ? _slots_15_io_uop_fp_single : _GEN_174 ? _slots_14_io_uop_fp_single : _GEN_168 ? _slots_13_io_uop_fp_single : _GEN_162 ? _slots_12_io_uop_fp_single : _GEN_156 ? _slots_11_io_uop_fp_single : _GEN_150 ? _slots_10_io_uop_fp_single : _GEN_144 ? _slots_9_io_uop_fp_single : _GEN_138 ? _slots_8_io_uop_fp_single : _GEN_132 ? _slots_7_io_uop_fp_single : _GEN_126 ? _slots_6_io_uop_fp_single : _GEN_120 ? _slots_5_io_uop_fp_single : _GEN_114 ? _slots_4_io_uop_fp_single : _GEN_108 ? _slots_3_io_uop_fp_single : _GEN_102 ? _slots_2_io_uop_fp_single : _GEN_96 ? _slots_1_io_uop_fp_single : _GEN_93 & _slots_0_io_uop_fp_single;
  assign io_iss_uops_0_xcpt_pf_if = _GEN_225 ? _slots_23_io_uop_xcpt_pf_if : _GEN_222 ? _slots_22_io_uop_xcpt_pf_if : _GEN_216 ? _slots_21_io_uop_xcpt_pf_if : _GEN_210 ? _slots_20_io_uop_xcpt_pf_if : _GEN_204 ? _slots_19_io_uop_xcpt_pf_if : _GEN_198 ? _slots_18_io_uop_xcpt_pf_if : _GEN_192 ? _slots_17_io_uop_xcpt_pf_if : _GEN_186 ? _slots_16_io_uop_xcpt_pf_if : _GEN_180 ? _slots_15_io_uop_xcpt_pf_if : _GEN_174 ? _slots_14_io_uop_xcpt_pf_if : _GEN_168 ? _slots_13_io_uop_xcpt_pf_if : _GEN_162 ? _slots_12_io_uop_xcpt_pf_if : _GEN_156 ? _slots_11_io_uop_xcpt_pf_if : _GEN_150 ? _slots_10_io_uop_xcpt_pf_if : _GEN_144 ? _slots_9_io_uop_xcpt_pf_if : _GEN_138 ? _slots_8_io_uop_xcpt_pf_if : _GEN_132 ? _slots_7_io_uop_xcpt_pf_if : _GEN_126 ? _slots_6_io_uop_xcpt_pf_if : _GEN_120 ? _slots_5_io_uop_xcpt_pf_if : _GEN_114 ? _slots_4_io_uop_xcpt_pf_if : _GEN_108 ? _slots_3_io_uop_xcpt_pf_if : _GEN_102 ? _slots_2_io_uop_xcpt_pf_if : _GEN_96 ? _slots_1_io_uop_xcpt_pf_if : _GEN_93 & _slots_0_io_uop_xcpt_pf_if;
  assign io_iss_uops_0_xcpt_ae_if = _GEN_225 ? _slots_23_io_uop_xcpt_ae_if : _GEN_222 ? _slots_22_io_uop_xcpt_ae_if : _GEN_216 ? _slots_21_io_uop_xcpt_ae_if : _GEN_210 ? _slots_20_io_uop_xcpt_ae_if : _GEN_204 ? _slots_19_io_uop_xcpt_ae_if : _GEN_198 ? _slots_18_io_uop_xcpt_ae_if : _GEN_192 ? _slots_17_io_uop_xcpt_ae_if : _GEN_186 ? _slots_16_io_uop_xcpt_ae_if : _GEN_180 ? _slots_15_io_uop_xcpt_ae_if : _GEN_174 ? _slots_14_io_uop_xcpt_ae_if : _GEN_168 ? _slots_13_io_uop_xcpt_ae_if : _GEN_162 ? _slots_12_io_uop_xcpt_ae_if : _GEN_156 ? _slots_11_io_uop_xcpt_ae_if : _GEN_150 ? _slots_10_io_uop_xcpt_ae_if : _GEN_144 ? _slots_9_io_uop_xcpt_ae_if : _GEN_138 ? _slots_8_io_uop_xcpt_ae_if : _GEN_132 ? _slots_7_io_uop_xcpt_ae_if : _GEN_126 ? _slots_6_io_uop_xcpt_ae_if : _GEN_120 ? _slots_5_io_uop_xcpt_ae_if : _GEN_114 ? _slots_4_io_uop_xcpt_ae_if : _GEN_108 ? _slots_3_io_uop_xcpt_ae_if : _GEN_102 ? _slots_2_io_uop_xcpt_ae_if : _GEN_96 ? _slots_1_io_uop_xcpt_ae_if : _GEN_93 & _slots_0_io_uop_xcpt_ae_if;
  assign io_iss_uops_0_xcpt_ma_if = _GEN_225 ? _slots_23_io_uop_xcpt_ma_if : _GEN_222 ? _slots_22_io_uop_xcpt_ma_if : _GEN_216 ? _slots_21_io_uop_xcpt_ma_if : _GEN_210 ? _slots_20_io_uop_xcpt_ma_if : _GEN_204 ? _slots_19_io_uop_xcpt_ma_if : _GEN_198 ? _slots_18_io_uop_xcpt_ma_if : _GEN_192 ? _slots_17_io_uop_xcpt_ma_if : _GEN_186 ? _slots_16_io_uop_xcpt_ma_if : _GEN_180 ? _slots_15_io_uop_xcpt_ma_if : _GEN_174 ? _slots_14_io_uop_xcpt_ma_if : _GEN_168 ? _slots_13_io_uop_xcpt_ma_if : _GEN_162 ? _slots_12_io_uop_xcpt_ma_if : _GEN_156 ? _slots_11_io_uop_xcpt_ma_if : _GEN_150 ? _slots_10_io_uop_xcpt_ma_if : _GEN_144 ? _slots_9_io_uop_xcpt_ma_if : _GEN_138 ? _slots_8_io_uop_xcpt_ma_if : _GEN_132 ? _slots_7_io_uop_xcpt_ma_if : _GEN_126 ? _slots_6_io_uop_xcpt_ma_if : _GEN_120 ? _slots_5_io_uop_xcpt_ma_if : _GEN_114 ? _slots_4_io_uop_xcpt_ma_if : _GEN_108 ? _slots_3_io_uop_xcpt_ma_if : _GEN_102 ? _slots_2_io_uop_xcpt_ma_if : _GEN_96 ? _slots_1_io_uop_xcpt_ma_if : _GEN_93 & _slots_0_io_uop_xcpt_ma_if;
  assign io_iss_uops_0_bp_debug_if = _GEN_225 ? _slots_23_io_uop_bp_debug_if : _GEN_222 ? _slots_22_io_uop_bp_debug_if : _GEN_216 ? _slots_21_io_uop_bp_debug_if : _GEN_210 ? _slots_20_io_uop_bp_debug_if : _GEN_204 ? _slots_19_io_uop_bp_debug_if : _GEN_198 ? _slots_18_io_uop_bp_debug_if : _GEN_192 ? _slots_17_io_uop_bp_debug_if : _GEN_186 ? _slots_16_io_uop_bp_debug_if : _GEN_180 ? _slots_15_io_uop_bp_debug_if : _GEN_174 ? _slots_14_io_uop_bp_debug_if : _GEN_168 ? _slots_13_io_uop_bp_debug_if : _GEN_162 ? _slots_12_io_uop_bp_debug_if : _GEN_156 ? _slots_11_io_uop_bp_debug_if : _GEN_150 ? _slots_10_io_uop_bp_debug_if : _GEN_144 ? _slots_9_io_uop_bp_debug_if : _GEN_138 ? _slots_8_io_uop_bp_debug_if : _GEN_132 ? _slots_7_io_uop_bp_debug_if : _GEN_126 ? _slots_6_io_uop_bp_debug_if : _GEN_120 ? _slots_5_io_uop_bp_debug_if : _GEN_114 ? _slots_4_io_uop_bp_debug_if : _GEN_108 ? _slots_3_io_uop_bp_debug_if : _GEN_102 ? _slots_2_io_uop_bp_debug_if : _GEN_96 ? _slots_1_io_uop_bp_debug_if : _GEN_93 & _slots_0_io_uop_bp_debug_if;
  assign io_iss_uops_0_bp_xcpt_if = _GEN_225 ? _slots_23_io_uop_bp_xcpt_if : _GEN_222 ? _slots_22_io_uop_bp_xcpt_if : _GEN_216 ? _slots_21_io_uop_bp_xcpt_if : _GEN_210 ? _slots_20_io_uop_bp_xcpt_if : _GEN_204 ? _slots_19_io_uop_bp_xcpt_if : _GEN_198 ? _slots_18_io_uop_bp_xcpt_if : _GEN_192 ? _slots_17_io_uop_bp_xcpt_if : _GEN_186 ? _slots_16_io_uop_bp_xcpt_if : _GEN_180 ? _slots_15_io_uop_bp_xcpt_if : _GEN_174 ? _slots_14_io_uop_bp_xcpt_if : _GEN_168 ? _slots_13_io_uop_bp_xcpt_if : _GEN_162 ? _slots_12_io_uop_bp_xcpt_if : _GEN_156 ? _slots_11_io_uop_bp_xcpt_if : _GEN_150 ? _slots_10_io_uop_bp_xcpt_if : _GEN_144 ? _slots_9_io_uop_bp_xcpt_if : _GEN_138 ? _slots_8_io_uop_bp_xcpt_if : _GEN_132 ? _slots_7_io_uop_bp_xcpt_if : _GEN_126 ? _slots_6_io_uop_bp_xcpt_if : _GEN_120 ? _slots_5_io_uop_bp_xcpt_if : _GEN_114 ? _slots_4_io_uop_bp_xcpt_if : _GEN_108 ? _slots_3_io_uop_bp_xcpt_if : _GEN_102 ? _slots_2_io_uop_bp_xcpt_if : _GEN_96 ? _slots_1_io_uop_bp_xcpt_if : _GEN_93 & _slots_0_io_uop_bp_xcpt_if;
  assign io_iss_uops_0_debug_fsrc = _GEN_225 ? _slots_23_io_uop_debug_fsrc : _GEN_222 ? _slots_22_io_uop_debug_fsrc : _GEN_216 ? _slots_21_io_uop_debug_fsrc : _GEN_210 ? _slots_20_io_uop_debug_fsrc : _GEN_204 ? _slots_19_io_uop_debug_fsrc : _GEN_198 ? _slots_18_io_uop_debug_fsrc : _GEN_192 ? _slots_17_io_uop_debug_fsrc : _GEN_186 ? _slots_16_io_uop_debug_fsrc : _GEN_180 ? _slots_15_io_uop_debug_fsrc : _GEN_174 ? _slots_14_io_uop_debug_fsrc : _GEN_168 ? _slots_13_io_uop_debug_fsrc : _GEN_162 ? _slots_12_io_uop_debug_fsrc : _GEN_156 ? _slots_11_io_uop_debug_fsrc : _GEN_150 ? _slots_10_io_uop_debug_fsrc : _GEN_144 ? _slots_9_io_uop_debug_fsrc : _GEN_138 ? _slots_8_io_uop_debug_fsrc : _GEN_132 ? _slots_7_io_uop_debug_fsrc : _GEN_126 ? _slots_6_io_uop_debug_fsrc : _GEN_120 ? _slots_5_io_uop_debug_fsrc : _GEN_114 ? _slots_4_io_uop_debug_fsrc : _GEN_108 ? _slots_3_io_uop_debug_fsrc : _GEN_102 ? _slots_2_io_uop_debug_fsrc : _GEN_96 ? _slots_1_io_uop_debug_fsrc : _GEN_93 ? _slots_0_io_uop_debug_fsrc : 2'h0;
  assign io_iss_uops_0_debug_tsrc = _GEN_225 ? _slots_23_io_uop_debug_tsrc : _GEN_222 ? _slots_22_io_uop_debug_tsrc : _GEN_216 ? _slots_21_io_uop_debug_tsrc : _GEN_210 ? _slots_20_io_uop_debug_tsrc : _GEN_204 ? _slots_19_io_uop_debug_tsrc : _GEN_198 ? _slots_18_io_uop_debug_tsrc : _GEN_192 ? _slots_17_io_uop_debug_tsrc : _GEN_186 ? _slots_16_io_uop_debug_tsrc : _GEN_180 ? _slots_15_io_uop_debug_tsrc : _GEN_174 ? _slots_14_io_uop_debug_tsrc : _GEN_168 ? _slots_13_io_uop_debug_tsrc : _GEN_162 ? _slots_12_io_uop_debug_tsrc : _GEN_156 ? _slots_11_io_uop_debug_tsrc : _GEN_150 ? _slots_10_io_uop_debug_tsrc : _GEN_144 ? _slots_9_io_uop_debug_tsrc : _GEN_138 ? _slots_8_io_uop_debug_tsrc : _GEN_132 ? _slots_7_io_uop_debug_tsrc : _GEN_126 ? _slots_6_io_uop_debug_tsrc : _GEN_120 ? _slots_5_io_uop_debug_tsrc : _GEN_114 ? _slots_4_io_uop_debug_tsrc : _GEN_108 ? _slots_3_io_uop_debug_tsrc : _GEN_102 ? _slots_2_io_uop_debug_tsrc : _GEN_96 ? _slots_1_io_uop_debug_tsrc : _GEN_93 ? _slots_0_io_uop_debug_tsrc : 2'h0;
  assign io_iss_uops_1_uopc = _GEN_226 ? _slots_23_io_uop_uopc : _GEN_224 ? _slots_22_io_uop_uopc : _GEN_219 ? _slots_21_io_uop_uopc : _GEN_213 ? _slots_20_io_uop_uopc : _GEN_207 ? _slots_19_io_uop_uopc : _GEN_201 ? _slots_18_io_uop_uopc : _GEN_195 ? _slots_17_io_uop_uopc : _GEN_189 ? _slots_16_io_uop_uopc : _GEN_183 ? _slots_15_io_uop_uopc : _GEN_177 ? _slots_14_io_uop_uopc : _GEN_171 ? _slots_13_io_uop_uopc : _GEN_165 ? _slots_12_io_uop_uopc : _GEN_159 ? _slots_11_io_uop_uopc : _GEN_153 ? _slots_10_io_uop_uopc : _GEN_147 ? _slots_9_io_uop_uopc : _GEN_141 ? _slots_8_io_uop_uopc : _GEN_135 ? _slots_7_io_uop_uopc : _GEN_129 ? _slots_6_io_uop_uopc : _GEN_123 ? _slots_5_io_uop_uopc : _GEN_117 ? _slots_4_io_uop_uopc : _GEN_111 ? _slots_3_io_uop_uopc : _GEN_105 ? _slots_2_io_uop_uopc : _GEN_99 ? _slots_1_io_uop_uopc : _GEN_94 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_1_inst = _GEN_226 ? _slots_23_io_uop_inst : _GEN_224 ? _slots_22_io_uop_inst : _GEN_219 ? _slots_21_io_uop_inst : _GEN_213 ? _slots_20_io_uop_inst : _GEN_207 ? _slots_19_io_uop_inst : _GEN_201 ? _slots_18_io_uop_inst : _GEN_195 ? _slots_17_io_uop_inst : _GEN_189 ? _slots_16_io_uop_inst : _GEN_183 ? _slots_15_io_uop_inst : _GEN_177 ? _slots_14_io_uop_inst : _GEN_171 ? _slots_13_io_uop_inst : _GEN_165 ? _slots_12_io_uop_inst : _GEN_159 ? _slots_11_io_uop_inst : _GEN_153 ? _slots_10_io_uop_inst : _GEN_147 ? _slots_9_io_uop_inst : _GEN_141 ? _slots_8_io_uop_inst : _GEN_135 ? _slots_7_io_uop_inst : _GEN_129 ? _slots_6_io_uop_inst : _GEN_123 ? _slots_5_io_uop_inst : _GEN_117 ? _slots_4_io_uop_inst : _GEN_111 ? _slots_3_io_uop_inst : _GEN_105 ? _slots_2_io_uop_inst : _GEN_99 ? _slots_1_io_uop_inst : _GEN_94 ? _slots_0_io_uop_inst : 32'h0;
  assign io_iss_uops_1_debug_inst = _GEN_226 ? _slots_23_io_uop_debug_inst : _GEN_224 ? _slots_22_io_uop_debug_inst : _GEN_219 ? _slots_21_io_uop_debug_inst : _GEN_213 ? _slots_20_io_uop_debug_inst : _GEN_207 ? _slots_19_io_uop_debug_inst : _GEN_201 ? _slots_18_io_uop_debug_inst : _GEN_195 ? _slots_17_io_uop_debug_inst : _GEN_189 ? _slots_16_io_uop_debug_inst : _GEN_183 ? _slots_15_io_uop_debug_inst : _GEN_177 ? _slots_14_io_uop_debug_inst : _GEN_171 ? _slots_13_io_uop_debug_inst : _GEN_165 ? _slots_12_io_uop_debug_inst : _GEN_159 ? _slots_11_io_uop_debug_inst : _GEN_153 ? _slots_10_io_uop_debug_inst : _GEN_147 ? _slots_9_io_uop_debug_inst : _GEN_141 ? _slots_8_io_uop_debug_inst : _GEN_135 ? _slots_7_io_uop_debug_inst : _GEN_129 ? _slots_6_io_uop_debug_inst : _GEN_123 ? _slots_5_io_uop_debug_inst : _GEN_117 ? _slots_4_io_uop_debug_inst : _GEN_111 ? _slots_3_io_uop_debug_inst : _GEN_105 ? _slots_2_io_uop_debug_inst : _GEN_99 ? _slots_1_io_uop_debug_inst : _GEN_94 ? _slots_0_io_uop_debug_inst : 32'h0;
  assign io_iss_uops_1_is_rvc = _GEN_226 ? _slots_23_io_uop_is_rvc : _GEN_224 ? _slots_22_io_uop_is_rvc : _GEN_219 ? _slots_21_io_uop_is_rvc : _GEN_213 ? _slots_20_io_uop_is_rvc : _GEN_207 ? _slots_19_io_uop_is_rvc : _GEN_201 ? _slots_18_io_uop_is_rvc : _GEN_195 ? _slots_17_io_uop_is_rvc : _GEN_189 ? _slots_16_io_uop_is_rvc : _GEN_183 ? _slots_15_io_uop_is_rvc : _GEN_177 ? _slots_14_io_uop_is_rvc : _GEN_171 ? _slots_13_io_uop_is_rvc : _GEN_165 ? _slots_12_io_uop_is_rvc : _GEN_159 ? _slots_11_io_uop_is_rvc : _GEN_153 ? _slots_10_io_uop_is_rvc : _GEN_147 ? _slots_9_io_uop_is_rvc : _GEN_141 ? _slots_8_io_uop_is_rvc : _GEN_135 ? _slots_7_io_uop_is_rvc : _GEN_129 ? _slots_6_io_uop_is_rvc : _GEN_123 ? _slots_5_io_uop_is_rvc : _GEN_117 ? _slots_4_io_uop_is_rvc : _GEN_111 ? _slots_3_io_uop_is_rvc : _GEN_105 ? _slots_2_io_uop_is_rvc : _GEN_99 ? _slots_1_io_uop_is_rvc : _GEN_94 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_1_debug_pc = _GEN_226 ? _slots_23_io_uop_debug_pc : _GEN_224 ? _slots_22_io_uop_debug_pc : _GEN_219 ? _slots_21_io_uop_debug_pc : _GEN_213 ? _slots_20_io_uop_debug_pc : _GEN_207 ? _slots_19_io_uop_debug_pc : _GEN_201 ? _slots_18_io_uop_debug_pc : _GEN_195 ? _slots_17_io_uop_debug_pc : _GEN_189 ? _slots_16_io_uop_debug_pc : _GEN_183 ? _slots_15_io_uop_debug_pc : _GEN_177 ? _slots_14_io_uop_debug_pc : _GEN_171 ? _slots_13_io_uop_debug_pc : _GEN_165 ? _slots_12_io_uop_debug_pc : _GEN_159 ? _slots_11_io_uop_debug_pc : _GEN_153 ? _slots_10_io_uop_debug_pc : _GEN_147 ? _slots_9_io_uop_debug_pc : _GEN_141 ? _slots_8_io_uop_debug_pc : _GEN_135 ? _slots_7_io_uop_debug_pc : _GEN_129 ? _slots_6_io_uop_debug_pc : _GEN_123 ? _slots_5_io_uop_debug_pc : _GEN_117 ? _slots_4_io_uop_debug_pc : _GEN_111 ? _slots_3_io_uop_debug_pc : _GEN_105 ? _slots_2_io_uop_debug_pc : _GEN_99 ? _slots_1_io_uop_debug_pc : _GEN_94 ? _slots_0_io_uop_debug_pc : 40'h0;
  assign io_iss_uops_1_iq_type = _GEN_226 ? _slots_23_io_uop_iq_type : _GEN_224 ? _slots_22_io_uop_iq_type : _GEN_219 ? _slots_21_io_uop_iq_type : _GEN_213 ? _slots_20_io_uop_iq_type : _GEN_207 ? _slots_19_io_uop_iq_type : _GEN_201 ? _slots_18_io_uop_iq_type : _GEN_195 ? _slots_17_io_uop_iq_type : _GEN_189 ? _slots_16_io_uop_iq_type : _GEN_183 ? _slots_15_io_uop_iq_type : _GEN_177 ? _slots_14_io_uop_iq_type : _GEN_171 ? _slots_13_io_uop_iq_type : _GEN_165 ? _slots_12_io_uop_iq_type : _GEN_159 ? _slots_11_io_uop_iq_type : _GEN_153 ? _slots_10_io_uop_iq_type : _GEN_147 ? _slots_9_io_uop_iq_type : _GEN_141 ? _slots_8_io_uop_iq_type : _GEN_135 ? _slots_7_io_uop_iq_type : _GEN_129 ? _slots_6_io_uop_iq_type : _GEN_123 ? _slots_5_io_uop_iq_type : _GEN_117 ? _slots_4_io_uop_iq_type : _GEN_111 ? _slots_3_io_uop_iq_type : _GEN_105 ? _slots_2_io_uop_iq_type : _GEN_99 ? _slots_1_io_uop_iq_type : _GEN_94 ? _slots_0_io_uop_iq_type : 3'h0;
  assign io_iss_uops_1_fu_code = _GEN_226 ? _slots_23_io_uop_fu_code : _GEN_224 ? _slots_22_io_uop_fu_code : _GEN_219 ? _slots_21_io_uop_fu_code : _GEN_213 ? _slots_20_io_uop_fu_code : _GEN_207 ? _slots_19_io_uop_fu_code : _GEN_201 ? _slots_18_io_uop_fu_code : _GEN_195 ? _slots_17_io_uop_fu_code : _GEN_189 ? _slots_16_io_uop_fu_code : _GEN_183 ? _slots_15_io_uop_fu_code : _GEN_177 ? _slots_14_io_uop_fu_code : _GEN_171 ? _slots_13_io_uop_fu_code : _GEN_165 ? _slots_12_io_uop_fu_code : _GEN_159 ? _slots_11_io_uop_fu_code : _GEN_153 ? _slots_10_io_uop_fu_code : _GEN_147 ? _slots_9_io_uop_fu_code : _GEN_141 ? _slots_8_io_uop_fu_code : _GEN_135 ? _slots_7_io_uop_fu_code : _GEN_129 ? _slots_6_io_uop_fu_code : _GEN_123 ? _slots_5_io_uop_fu_code : _GEN_117 ? _slots_4_io_uop_fu_code : _GEN_111 ? _slots_3_io_uop_fu_code : _GEN_105 ? _slots_2_io_uop_fu_code : _GEN_99 ? _slots_1_io_uop_fu_code : _GEN_94 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_1_iw_state = _GEN_226 ? _slots_23_io_uop_iw_state : _GEN_224 ? _slots_22_io_uop_iw_state : _GEN_219 ? _slots_21_io_uop_iw_state : _GEN_213 ? _slots_20_io_uop_iw_state : _GEN_207 ? _slots_19_io_uop_iw_state : _GEN_201 ? _slots_18_io_uop_iw_state : _GEN_195 ? _slots_17_io_uop_iw_state : _GEN_189 ? _slots_16_io_uop_iw_state : _GEN_183 ? _slots_15_io_uop_iw_state : _GEN_177 ? _slots_14_io_uop_iw_state : _GEN_171 ? _slots_13_io_uop_iw_state : _GEN_165 ? _slots_12_io_uop_iw_state : _GEN_159 ? _slots_11_io_uop_iw_state : _GEN_153 ? _slots_10_io_uop_iw_state : _GEN_147 ? _slots_9_io_uop_iw_state : _GEN_141 ? _slots_8_io_uop_iw_state : _GEN_135 ? _slots_7_io_uop_iw_state : _GEN_129 ? _slots_6_io_uop_iw_state : _GEN_123 ? _slots_5_io_uop_iw_state : _GEN_117 ? _slots_4_io_uop_iw_state : _GEN_111 ? _slots_3_io_uop_iw_state : _GEN_105 ? _slots_2_io_uop_iw_state : _GEN_99 ? _slots_1_io_uop_iw_state : _GEN_94 ? _slots_0_io_uop_iw_state : 2'h0;
  assign io_iss_uops_1_iw_p1_poisoned = _GEN_226 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_224 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_219 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_213 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_207 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_201 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_195 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_189 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_183 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_177 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_171 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_165 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_159 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_153 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_147 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_141 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_135 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_129 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_123 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_117 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_111 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_105 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_99 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_94 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_1_iw_p2_poisoned = _GEN_226 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_224 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_219 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_213 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_207 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_201 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_195 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_189 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_183 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_177 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_171 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_165 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_159 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_153 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_147 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_141 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_135 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_129 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_123 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_117 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_111 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_105 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_99 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_94 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_1_is_br = _GEN_226 ? _slots_23_io_uop_is_br : _GEN_224 ? _slots_22_io_uop_is_br : _GEN_219 ? _slots_21_io_uop_is_br : _GEN_213 ? _slots_20_io_uop_is_br : _GEN_207 ? _slots_19_io_uop_is_br : _GEN_201 ? _slots_18_io_uop_is_br : _GEN_195 ? _slots_17_io_uop_is_br : _GEN_189 ? _slots_16_io_uop_is_br : _GEN_183 ? _slots_15_io_uop_is_br : _GEN_177 ? _slots_14_io_uop_is_br : _GEN_171 ? _slots_13_io_uop_is_br : _GEN_165 ? _slots_12_io_uop_is_br : _GEN_159 ? _slots_11_io_uop_is_br : _GEN_153 ? _slots_10_io_uop_is_br : _GEN_147 ? _slots_9_io_uop_is_br : _GEN_141 ? _slots_8_io_uop_is_br : _GEN_135 ? _slots_7_io_uop_is_br : _GEN_129 ? _slots_6_io_uop_is_br : _GEN_123 ? _slots_5_io_uop_is_br : _GEN_117 ? _slots_4_io_uop_is_br : _GEN_111 ? _slots_3_io_uop_is_br : _GEN_105 ? _slots_2_io_uop_is_br : _GEN_99 ? _slots_1_io_uop_is_br : _GEN_94 & _slots_0_io_uop_is_br;
  assign io_iss_uops_1_is_jalr = _GEN_226 ? _slots_23_io_uop_is_jalr : _GEN_224 ? _slots_22_io_uop_is_jalr : _GEN_219 ? _slots_21_io_uop_is_jalr : _GEN_213 ? _slots_20_io_uop_is_jalr : _GEN_207 ? _slots_19_io_uop_is_jalr : _GEN_201 ? _slots_18_io_uop_is_jalr : _GEN_195 ? _slots_17_io_uop_is_jalr : _GEN_189 ? _slots_16_io_uop_is_jalr : _GEN_183 ? _slots_15_io_uop_is_jalr : _GEN_177 ? _slots_14_io_uop_is_jalr : _GEN_171 ? _slots_13_io_uop_is_jalr : _GEN_165 ? _slots_12_io_uop_is_jalr : _GEN_159 ? _slots_11_io_uop_is_jalr : _GEN_153 ? _slots_10_io_uop_is_jalr : _GEN_147 ? _slots_9_io_uop_is_jalr : _GEN_141 ? _slots_8_io_uop_is_jalr : _GEN_135 ? _slots_7_io_uop_is_jalr : _GEN_129 ? _slots_6_io_uop_is_jalr : _GEN_123 ? _slots_5_io_uop_is_jalr : _GEN_117 ? _slots_4_io_uop_is_jalr : _GEN_111 ? _slots_3_io_uop_is_jalr : _GEN_105 ? _slots_2_io_uop_is_jalr : _GEN_99 ? _slots_1_io_uop_is_jalr : _GEN_94 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_1_is_jal = _GEN_226 ? _slots_23_io_uop_is_jal : _GEN_224 ? _slots_22_io_uop_is_jal : _GEN_219 ? _slots_21_io_uop_is_jal : _GEN_213 ? _slots_20_io_uop_is_jal : _GEN_207 ? _slots_19_io_uop_is_jal : _GEN_201 ? _slots_18_io_uop_is_jal : _GEN_195 ? _slots_17_io_uop_is_jal : _GEN_189 ? _slots_16_io_uop_is_jal : _GEN_183 ? _slots_15_io_uop_is_jal : _GEN_177 ? _slots_14_io_uop_is_jal : _GEN_171 ? _slots_13_io_uop_is_jal : _GEN_165 ? _slots_12_io_uop_is_jal : _GEN_159 ? _slots_11_io_uop_is_jal : _GEN_153 ? _slots_10_io_uop_is_jal : _GEN_147 ? _slots_9_io_uop_is_jal : _GEN_141 ? _slots_8_io_uop_is_jal : _GEN_135 ? _slots_7_io_uop_is_jal : _GEN_129 ? _slots_6_io_uop_is_jal : _GEN_123 ? _slots_5_io_uop_is_jal : _GEN_117 ? _slots_4_io_uop_is_jal : _GEN_111 ? _slots_3_io_uop_is_jal : _GEN_105 ? _slots_2_io_uop_is_jal : _GEN_99 ? _slots_1_io_uop_is_jal : _GEN_94 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_1_is_sfb = _GEN_226 ? _slots_23_io_uop_is_sfb : _GEN_224 ? _slots_22_io_uop_is_sfb : _GEN_219 ? _slots_21_io_uop_is_sfb : _GEN_213 ? _slots_20_io_uop_is_sfb : _GEN_207 ? _slots_19_io_uop_is_sfb : _GEN_201 ? _slots_18_io_uop_is_sfb : _GEN_195 ? _slots_17_io_uop_is_sfb : _GEN_189 ? _slots_16_io_uop_is_sfb : _GEN_183 ? _slots_15_io_uop_is_sfb : _GEN_177 ? _slots_14_io_uop_is_sfb : _GEN_171 ? _slots_13_io_uop_is_sfb : _GEN_165 ? _slots_12_io_uop_is_sfb : _GEN_159 ? _slots_11_io_uop_is_sfb : _GEN_153 ? _slots_10_io_uop_is_sfb : _GEN_147 ? _slots_9_io_uop_is_sfb : _GEN_141 ? _slots_8_io_uop_is_sfb : _GEN_135 ? _slots_7_io_uop_is_sfb : _GEN_129 ? _slots_6_io_uop_is_sfb : _GEN_123 ? _slots_5_io_uop_is_sfb : _GEN_117 ? _slots_4_io_uop_is_sfb : _GEN_111 ? _slots_3_io_uop_is_sfb : _GEN_105 ? _slots_2_io_uop_is_sfb : _GEN_99 ? _slots_1_io_uop_is_sfb : _GEN_94 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_1_br_mask = _GEN_226 ? _slots_23_io_uop_br_mask : _GEN_224 ? _slots_22_io_uop_br_mask : _GEN_219 ? _slots_21_io_uop_br_mask : _GEN_213 ? _slots_20_io_uop_br_mask : _GEN_207 ? _slots_19_io_uop_br_mask : _GEN_201 ? _slots_18_io_uop_br_mask : _GEN_195 ? _slots_17_io_uop_br_mask : _GEN_189 ? _slots_16_io_uop_br_mask : _GEN_183 ? _slots_15_io_uop_br_mask : _GEN_177 ? _slots_14_io_uop_br_mask : _GEN_171 ? _slots_13_io_uop_br_mask : _GEN_165 ? _slots_12_io_uop_br_mask : _GEN_159 ? _slots_11_io_uop_br_mask : _GEN_153 ? _slots_10_io_uop_br_mask : _GEN_147 ? _slots_9_io_uop_br_mask : _GEN_141 ? _slots_8_io_uop_br_mask : _GEN_135 ? _slots_7_io_uop_br_mask : _GEN_129 ? _slots_6_io_uop_br_mask : _GEN_123 ? _slots_5_io_uop_br_mask : _GEN_117 ? _slots_4_io_uop_br_mask : _GEN_111 ? _slots_3_io_uop_br_mask : _GEN_105 ? _slots_2_io_uop_br_mask : _GEN_99 ? _slots_1_io_uop_br_mask : _GEN_94 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_1_br_tag = _GEN_226 ? _slots_23_io_uop_br_tag : _GEN_224 ? _slots_22_io_uop_br_tag : _GEN_219 ? _slots_21_io_uop_br_tag : _GEN_213 ? _slots_20_io_uop_br_tag : _GEN_207 ? _slots_19_io_uop_br_tag : _GEN_201 ? _slots_18_io_uop_br_tag : _GEN_195 ? _slots_17_io_uop_br_tag : _GEN_189 ? _slots_16_io_uop_br_tag : _GEN_183 ? _slots_15_io_uop_br_tag : _GEN_177 ? _slots_14_io_uop_br_tag : _GEN_171 ? _slots_13_io_uop_br_tag : _GEN_165 ? _slots_12_io_uop_br_tag : _GEN_159 ? _slots_11_io_uop_br_tag : _GEN_153 ? _slots_10_io_uop_br_tag : _GEN_147 ? _slots_9_io_uop_br_tag : _GEN_141 ? _slots_8_io_uop_br_tag : _GEN_135 ? _slots_7_io_uop_br_tag : _GEN_129 ? _slots_6_io_uop_br_tag : _GEN_123 ? _slots_5_io_uop_br_tag : _GEN_117 ? _slots_4_io_uop_br_tag : _GEN_111 ? _slots_3_io_uop_br_tag : _GEN_105 ? _slots_2_io_uop_br_tag : _GEN_99 ? _slots_1_io_uop_br_tag : _GEN_94 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_1_ftq_idx = _GEN_226 ? _slots_23_io_uop_ftq_idx : _GEN_224 ? _slots_22_io_uop_ftq_idx : _GEN_219 ? _slots_21_io_uop_ftq_idx : _GEN_213 ? _slots_20_io_uop_ftq_idx : _GEN_207 ? _slots_19_io_uop_ftq_idx : _GEN_201 ? _slots_18_io_uop_ftq_idx : _GEN_195 ? _slots_17_io_uop_ftq_idx : _GEN_189 ? _slots_16_io_uop_ftq_idx : _GEN_183 ? _slots_15_io_uop_ftq_idx : _GEN_177 ? _slots_14_io_uop_ftq_idx : _GEN_171 ? _slots_13_io_uop_ftq_idx : _GEN_165 ? _slots_12_io_uop_ftq_idx : _GEN_159 ? _slots_11_io_uop_ftq_idx : _GEN_153 ? _slots_10_io_uop_ftq_idx : _GEN_147 ? _slots_9_io_uop_ftq_idx : _GEN_141 ? _slots_8_io_uop_ftq_idx : _GEN_135 ? _slots_7_io_uop_ftq_idx : _GEN_129 ? _slots_6_io_uop_ftq_idx : _GEN_123 ? _slots_5_io_uop_ftq_idx : _GEN_117 ? _slots_4_io_uop_ftq_idx : _GEN_111 ? _slots_3_io_uop_ftq_idx : _GEN_105 ? _slots_2_io_uop_ftq_idx : _GEN_99 ? _slots_1_io_uop_ftq_idx : _GEN_94 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_1_edge_inst = _GEN_226 ? _slots_23_io_uop_edge_inst : _GEN_224 ? _slots_22_io_uop_edge_inst : _GEN_219 ? _slots_21_io_uop_edge_inst : _GEN_213 ? _slots_20_io_uop_edge_inst : _GEN_207 ? _slots_19_io_uop_edge_inst : _GEN_201 ? _slots_18_io_uop_edge_inst : _GEN_195 ? _slots_17_io_uop_edge_inst : _GEN_189 ? _slots_16_io_uop_edge_inst : _GEN_183 ? _slots_15_io_uop_edge_inst : _GEN_177 ? _slots_14_io_uop_edge_inst : _GEN_171 ? _slots_13_io_uop_edge_inst : _GEN_165 ? _slots_12_io_uop_edge_inst : _GEN_159 ? _slots_11_io_uop_edge_inst : _GEN_153 ? _slots_10_io_uop_edge_inst : _GEN_147 ? _slots_9_io_uop_edge_inst : _GEN_141 ? _slots_8_io_uop_edge_inst : _GEN_135 ? _slots_7_io_uop_edge_inst : _GEN_129 ? _slots_6_io_uop_edge_inst : _GEN_123 ? _slots_5_io_uop_edge_inst : _GEN_117 ? _slots_4_io_uop_edge_inst : _GEN_111 ? _slots_3_io_uop_edge_inst : _GEN_105 ? _slots_2_io_uop_edge_inst : _GEN_99 ? _slots_1_io_uop_edge_inst : _GEN_94 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_1_pc_lob = _GEN_226 ? _slots_23_io_uop_pc_lob : _GEN_224 ? _slots_22_io_uop_pc_lob : _GEN_219 ? _slots_21_io_uop_pc_lob : _GEN_213 ? _slots_20_io_uop_pc_lob : _GEN_207 ? _slots_19_io_uop_pc_lob : _GEN_201 ? _slots_18_io_uop_pc_lob : _GEN_195 ? _slots_17_io_uop_pc_lob : _GEN_189 ? _slots_16_io_uop_pc_lob : _GEN_183 ? _slots_15_io_uop_pc_lob : _GEN_177 ? _slots_14_io_uop_pc_lob : _GEN_171 ? _slots_13_io_uop_pc_lob : _GEN_165 ? _slots_12_io_uop_pc_lob : _GEN_159 ? _slots_11_io_uop_pc_lob : _GEN_153 ? _slots_10_io_uop_pc_lob : _GEN_147 ? _slots_9_io_uop_pc_lob : _GEN_141 ? _slots_8_io_uop_pc_lob : _GEN_135 ? _slots_7_io_uop_pc_lob : _GEN_129 ? _slots_6_io_uop_pc_lob : _GEN_123 ? _slots_5_io_uop_pc_lob : _GEN_117 ? _slots_4_io_uop_pc_lob : _GEN_111 ? _slots_3_io_uop_pc_lob : _GEN_105 ? _slots_2_io_uop_pc_lob : _GEN_99 ? _slots_1_io_uop_pc_lob : _GEN_94 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_1_taken = _GEN_226 ? _slots_23_io_uop_taken : _GEN_224 ? _slots_22_io_uop_taken : _GEN_219 ? _slots_21_io_uop_taken : _GEN_213 ? _slots_20_io_uop_taken : _GEN_207 ? _slots_19_io_uop_taken : _GEN_201 ? _slots_18_io_uop_taken : _GEN_195 ? _slots_17_io_uop_taken : _GEN_189 ? _slots_16_io_uop_taken : _GEN_183 ? _slots_15_io_uop_taken : _GEN_177 ? _slots_14_io_uop_taken : _GEN_171 ? _slots_13_io_uop_taken : _GEN_165 ? _slots_12_io_uop_taken : _GEN_159 ? _slots_11_io_uop_taken : _GEN_153 ? _slots_10_io_uop_taken : _GEN_147 ? _slots_9_io_uop_taken : _GEN_141 ? _slots_8_io_uop_taken : _GEN_135 ? _slots_7_io_uop_taken : _GEN_129 ? _slots_6_io_uop_taken : _GEN_123 ? _slots_5_io_uop_taken : _GEN_117 ? _slots_4_io_uop_taken : _GEN_111 ? _slots_3_io_uop_taken : _GEN_105 ? _slots_2_io_uop_taken : _GEN_99 ? _slots_1_io_uop_taken : _GEN_94 & _slots_0_io_uop_taken;
  assign io_iss_uops_1_imm_packed = _GEN_226 ? _slots_23_io_uop_imm_packed : _GEN_224 ? _slots_22_io_uop_imm_packed : _GEN_219 ? _slots_21_io_uop_imm_packed : _GEN_213 ? _slots_20_io_uop_imm_packed : _GEN_207 ? _slots_19_io_uop_imm_packed : _GEN_201 ? _slots_18_io_uop_imm_packed : _GEN_195 ? _slots_17_io_uop_imm_packed : _GEN_189 ? _slots_16_io_uop_imm_packed : _GEN_183 ? _slots_15_io_uop_imm_packed : _GEN_177 ? _slots_14_io_uop_imm_packed : _GEN_171 ? _slots_13_io_uop_imm_packed : _GEN_165 ? _slots_12_io_uop_imm_packed : _GEN_159 ? _slots_11_io_uop_imm_packed : _GEN_153 ? _slots_10_io_uop_imm_packed : _GEN_147 ? _slots_9_io_uop_imm_packed : _GEN_141 ? _slots_8_io_uop_imm_packed : _GEN_135 ? _slots_7_io_uop_imm_packed : _GEN_129 ? _slots_6_io_uop_imm_packed : _GEN_123 ? _slots_5_io_uop_imm_packed : _GEN_117 ? _slots_4_io_uop_imm_packed : _GEN_111 ? _slots_3_io_uop_imm_packed : _GEN_105 ? _slots_2_io_uop_imm_packed : _GEN_99 ? _slots_1_io_uop_imm_packed : _GEN_94 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_1_csr_addr = _GEN_226 ? _slots_23_io_uop_csr_addr : _GEN_224 ? _slots_22_io_uop_csr_addr : _GEN_219 ? _slots_21_io_uop_csr_addr : _GEN_213 ? _slots_20_io_uop_csr_addr : _GEN_207 ? _slots_19_io_uop_csr_addr : _GEN_201 ? _slots_18_io_uop_csr_addr : _GEN_195 ? _slots_17_io_uop_csr_addr : _GEN_189 ? _slots_16_io_uop_csr_addr : _GEN_183 ? _slots_15_io_uop_csr_addr : _GEN_177 ? _slots_14_io_uop_csr_addr : _GEN_171 ? _slots_13_io_uop_csr_addr : _GEN_165 ? _slots_12_io_uop_csr_addr : _GEN_159 ? _slots_11_io_uop_csr_addr : _GEN_153 ? _slots_10_io_uop_csr_addr : _GEN_147 ? _slots_9_io_uop_csr_addr : _GEN_141 ? _slots_8_io_uop_csr_addr : _GEN_135 ? _slots_7_io_uop_csr_addr : _GEN_129 ? _slots_6_io_uop_csr_addr : _GEN_123 ? _slots_5_io_uop_csr_addr : _GEN_117 ? _slots_4_io_uop_csr_addr : _GEN_111 ? _slots_3_io_uop_csr_addr : _GEN_105 ? _slots_2_io_uop_csr_addr : _GEN_99 ? _slots_1_io_uop_csr_addr : _GEN_94 ? _slots_0_io_uop_csr_addr : 12'h0;
  assign io_iss_uops_1_rob_idx = _GEN_226 ? _slots_23_io_uop_rob_idx : _GEN_224 ? _slots_22_io_uop_rob_idx : _GEN_219 ? _slots_21_io_uop_rob_idx : _GEN_213 ? _slots_20_io_uop_rob_idx : _GEN_207 ? _slots_19_io_uop_rob_idx : _GEN_201 ? _slots_18_io_uop_rob_idx : _GEN_195 ? _slots_17_io_uop_rob_idx : _GEN_189 ? _slots_16_io_uop_rob_idx : _GEN_183 ? _slots_15_io_uop_rob_idx : _GEN_177 ? _slots_14_io_uop_rob_idx : _GEN_171 ? _slots_13_io_uop_rob_idx : _GEN_165 ? _slots_12_io_uop_rob_idx : _GEN_159 ? _slots_11_io_uop_rob_idx : _GEN_153 ? _slots_10_io_uop_rob_idx : _GEN_147 ? _slots_9_io_uop_rob_idx : _GEN_141 ? _slots_8_io_uop_rob_idx : _GEN_135 ? _slots_7_io_uop_rob_idx : _GEN_129 ? _slots_6_io_uop_rob_idx : _GEN_123 ? _slots_5_io_uop_rob_idx : _GEN_117 ? _slots_4_io_uop_rob_idx : _GEN_111 ? _slots_3_io_uop_rob_idx : _GEN_105 ? _slots_2_io_uop_rob_idx : _GEN_99 ? _slots_1_io_uop_rob_idx : _GEN_94 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_1_ldq_idx = _GEN_226 ? _slots_23_io_uop_ldq_idx : _GEN_224 ? _slots_22_io_uop_ldq_idx : _GEN_219 ? _slots_21_io_uop_ldq_idx : _GEN_213 ? _slots_20_io_uop_ldq_idx : _GEN_207 ? _slots_19_io_uop_ldq_idx : _GEN_201 ? _slots_18_io_uop_ldq_idx : _GEN_195 ? _slots_17_io_uop_ldq_idx : _GEN_189 ? _slots_16_io_uop_ldq_idx : _GEN_183 ? _slots_15_io_uop_ldq_idx : _GEN_177 ? _slots_14_io_uop_ldq_idx : _GEN_171 ? _slots_13_io_uop_ldq_idx : _GEN_165 ? _slots_12_io_uop_ldq_idx : _GEN_159 ? _slots_11_io_uop_ldq_idx : _GEN_153 ? _slots_10_io_uop_ldq_idx : _GEN_147 ? _slots_9_io_uop_ldq_idx : _GEN_141 ? _slots_8_io_uop_ldq_idx : _GEN_135 ? _slots_7_io_uop_ldq_idx : _GEN_129 ? _slots_6_io_uop_ldq_idx : _GEN_123 ? _slots_5_io_uop_ldq_idx : _GEN_117 ? _slots_4_io_uop_ldq_idx : _GEN_111 ? _slots_3_io_uop_ldq_idx : _GEN_105 ? _slots_2_io_uop_ldq_idx : _GEN_99 ? _slots_1_io_uop_ldq_idx : _GEN_94 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_1_stq_idx = _GEN_226 ? _slots_23_io_uop_stq_idx : _GEN_224 ? _slots_22_io_uop_stq_idx : _GEN_219 ? _slots_21_io_uop_stq_idx : _GEN_213 ? _slots_20_io_uop_stq_idx : _GEN_207 ? _slots_19_io_uop_stq_idx : _GEN_201 ? _slots_18_io_uop_stq_idx : _GEN_195 ? _slots_17_io_uop_stq_idx : _GEN_189 ? _slots_16_io_uop_stq_idx : _GEN_183 ? _slots_15_io_uop_stq_idx : _GEN_177 ? _slots_14_io_uop_stq_idx : _GEN_171 ? _slots_13_io_uop_stq_idx : _GEN_165 ? _slots_12_io_uop_stq_idx : _GEN_159 ? _slots_11_io_uop_stq_idx : _GEN_153 ? _slots_10_io_uop_stq_idx : _GEN_147 ? _slots_9_io_uop_stq_idx : _GEN_141 ? _slots_8_io_uop_stq_idx : _GEN_135 ? _slots_7_io_uop_stq_idx : _GEN_129 ? _slots_6_io_uop_stq_idx : _GEN_123 ? _slots_5_io_uop_stq_idx : _GEN_117 ? _slots_4_io_uop_stq_idx : _GEN_111 ? _slots_3_io_uop_stq_idx : _GEN_105 ? _slots_2_io_uop_stq_idx : _GEN_99 ? _slots_1_io_uop_stq_idx : _GEN_94 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_1_rxq_idx = _GEN_226 ? _slots_23_io_uop_rxq_idx : _GEN_224 ? _slots_22_io_uop_rxq_idx : _GEN_219 ? _slots_21_io_uop_rxq_idx : _GEN_213 ? _slots_20_io_uop_rxq_idx : _GEN_207 ? _slots_19_io_uop_rxq_idx : _GEN_201 ? _slots_18_io_uop_rxq_idx : _GEN_195 ? _slots_17_io_uop_rxq_idx : _GEN_189 ? _slots_16_io_uop_rxq_idx : _GEN_183 ? _slots_15_io_uop_rxq_idx : _GEN_177 ? _slots_14_io_uop_rxq_idx : _GEN_171 ? _slots_13_io_uop_rxq_idx : _GEN_165 ? _slots_12_io_uop_rxq_idx : _GEN_159 ? _slots_11_io_uop_rxq_idx : _GEN_153 ? _slots_10_io_uop_rxq_idx : _GEN_147 ? _slots_9_io_uop_rxq_idx : _GEN_141 ? _slots_8_io_uop_rxq_idx : _GEN_135 ? _slots_7_io_uop_rxq_idx : _GEN_129 ? _slots_6_io_uop_rxq_idx : _GEN_123 ? _slots_5_io_uop_rxq_idx : _GEN_117 ? _slots_4_io_uop_rxq_idx : _GEN_111 ? _slots_3_io_uop_rxq_idx : _GEN_105 ? _slots_2_io_uop_rxq_idx : _GEN_99 ? _slots_1_io_uop_rxq_idx : _GEN_94 ? _slots_0_io_uop_rxq_idx : 2'h0;
  assign io_iss_uops_1_pdst = _GEN_226 ? _slots_23_io_uop_pdst : _GEN_224 ? _slots_22_io_uop_pdst : _GEN_219 ? _slots_21_io_uop_pdst : _GEN_213 ? _slots_20_io_uop_pdst : _GEN_207 ? _slots_19_io_uop_pdst : _GEN_201 ? _slots_18_io_uop_pdst : _GEN_195 ? _slots_17_io_uop_pdst : _GEN_189 ? _slots_16_io_uop_pdst : _GEN_183 ? _slots_15_io_uop_pdst : _GEN_177 ? _slots_14_io_uop_pdst : _GEN_171 ? _slots_13_io_uop_pdst : _GEN_165 ? _slots_12_io_uop_pdst : _GEN_159 ? _slots_11_io_uop_pdst : _GEN_153 ? _slots_10_io_uop_pdst : _GEN_147 ? _slots_9_io_uop_pdst : _GEN_141 ? _slots_8_io_uop_pdst : _GEN_135 ? _slots_7_io_uop_pdst : _GEN_129 ? _slots_6_io_uop_pdst : _GEN_123 ? _slots_5_io_uop_pdst : _GEN_117 ? _slots_4_io_uop_pdst : _GEN_111 ? _slots_3_io_uop_pdst : _GEN_105 ? _slots_2_io_uop_pdst : _GEN_99 ? _slots_1_io_uop_pdst : _GEN_94 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_1_prs1 = _GEN_226 ? _slots_23_io_uop_prs1 : _GEN_224 ? _slots_22_io_uop_prs1 : _GEN_219 ? _slots_21_io_uop_prs1 : _GEN_213 ? _slots_20_io_uop_prs1 : _GEN_207 ? _slots_19_io_uop_prs1 : _GEN_201 ? _slots_18_io_uop_prs1 : _GEN_195 ? _slots_17_io_uop_prs1 : _GEN_189 ? _slots_16_io_uop_prs1 : _GEN_183 ? _slots_15_io_uop_prs1 : _GEN_177 ? _slots_14_io_uop_prs1 : _GEN_171 ? _slots_13_io_uop_prs1 : _GEN_165 ? _slots_12_io_uop_prs1 : _GEN_159 ? _slots_11_io_uop_prs1 : _GEN_153 ? _slots_10_io_uop_prs1 : _GEN_147 ? _slots_9_io_uop_prs1 : _GEN_141 ? _slots_8_io_uop_prs1 : _GEN_135 ? _slots_7_io_uop_prs1 : _GEN_129 ? _slots_6_io_uop_prs1 : _GEN_123 ? _slots_5_io_uop_prs1 : _GEN_117 ? _slots_4_io_uop_prs1 : _GEN_111 ? _slots_3_io_uop_prs1 : _GEN_105 ? _slots_2_io_uop_prs1 : _GEN_99 ? _slots_1_io_uop_prs1 : _GEN_94 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_1_prs2 = _GEN_226 ? _slots_23_io_uop_prs2 : _GEN_224 ? _slots_22_io_uop_prs2 : _GEN_219 ? _slots_21_io_uop_prs2 : _GEN_213 ? _slots_20_io_uop_prs2 : _GEN_207 ? _slots_19_io_uop_prs2 : _GEN_201 ? _slots_18_io_uop_prs2 : _GEN_195 ? _slots_17_io_uop_prs2 : _GEN_189 ? _slots_16_io_uop_prs2 : _GEN_183 ? _slots_15_io_uop_prs2 : _GEN_177 ? _slots_14_io_uop_prs2 : _GEN_171 ? _slots_13_io_uop_prs2 : _GEN_165 ? _slots_12_io_uop_prs2 : _GEN_159 ? _slots_11_io_uop_prs2 : _GEN_153 ? _slots_10_io_uop_prs2 : _GEN_147 ? _slots_9_io_uop_prs2 : _GEN_141 ? _slots_8_io_uop_prs2 : _GEN_135 ? _slots_7_io_uop_prs2 : _GEN_129 ? _slots_6_io_uop_prs2 : _GEN_123 ? _slots_5_io_uop_prs2 : _GEN_117 ? _slots_4_io_uop_prs2 : _GEN_111 ? _slots_3_io_uop_prs2 : _GEN_105 ? _slots_2_io_uop_prs2 : _GEN_99 ? _slots_1_io_uop_prs2 : _GEN_94 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_1_prs3 = _GEN_226 ? _slots_23_io_uop_prs3 : _GEN_224 ? _slots_22_io_uop_prs3 : _GEN_219 ? _slots_21_io_uop_prs3 : _GEN_213 ? _slots_20_io_uop_prs3 : _GEN_207 ? _slots_19_io_uop_prs3 : _GEN_201 ? _slots_18_io_uop_prs3 : _GEN_195 ? _slots_17_io_uop_prs3 : _GEN_189 ? _slots_16_io_uop_prs3 : _GEN_183 ? _slots_15_io_uop_prs3 : _GEN_177 ? _slots_14_io_uop_prs3 : _GEN_171 ? _slots_13_io_uop_prs3 : _GEN_165 ? _slots_12_io_uop_prs3 : _GEN_159 ? _slots_11_io_uop_prs3 : _GEN_153 ? _slots_10_io_uop_prs3 : _GEN_147 ? _slots_9_io_uop_prs3 : _GEN_141 ? _slots_8_io_uop_prs3 : _GEN_135 ? _slots_7_io_uop_prs3 : _GEN_129 ? _slots_6_io_uop_prs3 : _GEN_123 ? _slots_5_io_uop_prs3 : _GEN_117 ? _slots_4_io_uop_prs3 : _GEN_111 ? _slots_3_io_uop_prs3 : _GEN_105 ? _slots_2_io_uop_prs3 : _GEN_99 ? _slots_1_io_uop_prs3 : _GEN_94 ? _slots_0_io_uop_prs3 : 7'h0;
  assign io_iss_uops_1_ppred = _GEN_226 ? _slots_23_io_uop_ppred : _GEN_224 ? _slots_22_io_uop_ppred : _GEN_219 ? _slots_21_io_uop_ppred : _GEN_213 ? _slots_20_io_uop_ppred : _GEN_207 ? _slots_19_io_uop_ppred : _GEN_201 ? _slots_18_io_uop_ppred : _GEN_195 ? _slots_17_io_uop_ppred : _GEN_189 ? _slots_16_io_uop_ppred : _GEN_183 ? _slots_15_io_uop_ppred : _GEN_177 ? _slots_14_io_uop_ppred : _GEN_171 ? _slots_13_io_uop_ppred : _GEN_165 ? _slots_12_io_uop_ppred : _GEN_159 ? _slots_11_io_uop_ppred : _GEN_153 ? _slots_10_io_uop_ppred : _GEN_147 ? _slots_9_io_uop_ppred : _GEN_141 ? _slots_8_io_uop_ppred : _GEN_135 ? _slots_7_io_uop_ppred : _GEN_129 ? _slots_6_io_uop_ppred : _GEN_123 ? _slots_5_io_uop_ppred : _GEN_117 ? _slots_4_io_uop_ppred : _GEN_111 ? _slots_3_io_uop_ppred : _GEN_105 ? _slots_2_io_uop_ppred : _GEN_99 ? _slots_1_io_uop_ppred : _GEN_94 ? _slots_0_io_uop_ppred : 6'h0;
  assign io_iss_uops_1_prs1_busy = _GEN_226 ? _slots_23_io_uop_prs1_busy : _GEN_224 ? _slots_22_io_uop_prs1_busy : _GEN_219 ? _slots_21_io_uop_prs1_busy : _GEN_213 ? _slots_20_io_uop_prs1_busy : _GEN_207 ? _slots_19_io_uop_prs1_busy : _GEN_201 ? _slots_18_io_uop_prs1_busy : _GEN_195 ? _slots_17_io_uop_prs1_busy : _GEN_189 ? _slots_16_io_uop_prs1_busy : _GEN_183 ? _slots_15_io_uop_prs1_busy : _GEN_177 ? _slots_14_io_uop_prs1_busy : _GEN_171 ? _slots_13_io_uop_prs1_busy : _GEN_165 ? _slots_12_io_uop_prs1_busy : _GEN_159 ? _slots_11_io_uop_prs1_busy : _GEN_153 ? _slots_10_io_uop_prs1_busy : _GEN_147 ? _slots_9_io_uop_prs1_busy : _GEN_141 ? _slots_8_io_uop_prs1_busy : _GEN_135 ? _slots_7_io_uop_prs1_busy : _GEN_129 ? _slots_6_io_uop_prs1_busy : _GEN_123 ? _slots_5_io_uop_prs1_busy : _GEN_117 ? _slots_4_io_uop_prs1_busy : _GEN_111 ? _slots_3_io_uop_prs1_busy : _GEN_105 ? _slots_2_io_uop_prs1_busy : _GEN_99 ? _slots_1_io_uop_prs1_busy : _GEN_94 & _slots_0_io_uop_prs1_busy;
  assign io_iss_uops_1_prs2_busy = _GEN_226 ? _slots_23_io_uop_prs2_busy : _GEN_224 ? _slots_22_io_uop_prs2_busy : _GEN_219 ? _slots_21_io_uop_prs2_busy : _GEN_213 ? _slots_20_io_uop_prs2_busy : _GEN_207 ? _slots_19_io_uop_prs2_busy : _GEN_201 ? _slots_18_io_uop_prs2_busy : _GEN_195 ? _slots_17_io_uop_prs2_busy : _GEN_189 ? _slots_16_io_uop_prs2_busy : _GEN_183 ? _slots_15_io_uop_prs2_busy : _GEN_177 ? _slots_14_io_uop_prs2_busy : _GEN_171 ? _slots_13_io_uop_prs2_busy : _GEN_165 ? _slots_12_io_uop_prs2_busy : _GEN_159 ? _slots_11_io_uop_prs2_busy : _GEN_153 ? _slots_10_io_uop_prs2_busy : _GEN_147 ? _slots_9_io_uop_prs2_busy : _GEN_141 ? _slots_8_io_uop_prs2_busy : _GEN_135 ? _slots_7_io_uop_prs2_busy : _GEN_129 ? _slots_6_io_uop_prs2_busy : _GEN_123 ? _slots_5_io_uop_prs2_busy : _GEN_117 ? _slots_4_io_uop_prs2_busy : _GEN_111 ? _slots_3_io_uop_prs2_busy : _GEN_105 ? _slots_2_io_uop_prs2_busy : _GEN_99 ? _slots_1_io_uop_prs2_busy : _GEN_94 & _slots_0_io_uop_prs2_busy;
  assign io_iss_uops_1_prs3_busy = _GEN_226 ? _slots_23_io_uop_prs3_busy : _GEN_224 ? _slots_22_io_uop_prs3_busy : _GEN_219 ? _slots_21_io_uop_prs3_busy : _GEN_213 ? _slots_20_io_uop_prs3_busy : _GEN_207 ? _slots_19_io_uop_prs3_busy : _GEN_201 ? _slots_18_io_uop_prs3_busy : _GEN_195 ? _slots_17_io_uop_prs3_busy : _GEN_189 ? _slots_16_io_uop_prs3_busy : _GEN_183 ? _slots_15_io_uop_prs3_busy : _GEN_177 ? _slots_14_io_uop_prs3_busy : _GEN_171 ? _slots_13_io_uop_prs3_busy : _GEN_165 ? _slots_12_io_uop_prs3_busy : _GEN_159 ? _slots_11_io_uop_prs3_busy : _GEN_153 ? _slots_10_io_uop_prs3_busy : _GEN_147 ? _slots_9_io_uop_prs3_busy : _GEN_141 ? _slots_8_io_uop_prs3_busy : _GEN_135 ? _slots_7_io_uop_prs3_busy : _GEN_129 ? _slots_6_io_uop_prs3_busy : _GEN_123 ? _slots_5_io_uop_prs3_busy : _GEN_117 ? _slots_4_io_uop_prs3_busy : _GEN_111 ? _slots_3_io_uop_prs3_busy : _GEN_105 ? _slots_2_io_uop_prs3_busy : _GEN_99 ? _slots_1_io_uop_prs3_busy : _GEN_94 & _slots_0_io_uop_prs3_busy;
  assign io_iss_uops_1_ppred_busy = _GEN_226 ? _slots_23_io_uop_ppred_busy : _GEN_224 ? _slots_22_io_uop_ppred_busy : _GEN_219 ? _slots_21_io_uop_ppred_busy : _GEN_213 ? _slots_20_io_uop_ppred_busy : _GEN_207 ? _slots_19_io_uop_ppred_busy : _GEN_201 ? _slots_18_io_uop_ppred_busy : _GEN_195 ? _slots_17_io_uop_ppred_busy : _GEN_189 ? _slots_16_io_uop_ppred_busy : _GEN_183 ? _slots_15_io_uop_ppred_busy : _GEN_177 ? _slots_14_io_uop_ppred_busy : _GEN_171 ? _slots_13_io_uop_ppred_busy : _GEN_165 ? _slots_12_io_uop_ppred_busy : _GEN_159 ? _slots_11_io_uop_ppred_busy : _GEN_153 ? _slots_10_io_uop_ppred_busy : _GEN_147 ? _slots_9_io_uop_ppred_busy : _GEN_141 ? _slots_8_io_uop_ppred_busy : _GEN_135 ? _slots_7_io_uop_ppred_busy : _GEN_129 ? _slots_6_io_uop_ppred_busy : _GEN_123 ? _slots_5_io_uop_ppred_busy : _GEN_117 ? _slots_4_io_uop_ppred_busy : _GEN_111 ? _slots_3_io_uop_ppred_busy : _GEN_105 ? _slots_2_io_uop_ppred_busy : _GEN_99 ? _slots_1_io_uop_ppred_busy : _GEN_94 & _slots_0_io_uop_ppred_busy;
  assign io_iss_uops_1_stale_pdst = _GEN_226 ? _slots_23_io_uop_stale_pdst : _GEN_224 ? _slots_22_io_uop_stale_pdst : _GEN_219 ? _slots_21_io_uop_stale_pdst : _GEN_213 ? _slots_20_io_uop_stale_pdst : _GEN_207 ? _slots_19_io_uop_stale_pdst : _GEN_201 ? _slots_18_io_uop_stale_pdst : _GEN_195 ? _slots_17_io_uop_stale_pdst : _GEN_189 ? _slots_16_io_uop_stale_pdst : _GEN_183 ? _slots_15_io_uop_stale_pdst : _GEN_177 ? _slots_14_io_uop_stale_pdst : _GEN_171 ? _slots_13_io_uop_stale_pdst : _GEN_165 ? _slots_12_io_uop_stale_pdst : _GEN_159 ? _slots_11_io_uop_stale_pdst : _GEN_153 ? _slots_10_io_uop_stale_pdst : _GEN_147 ? _slots_9_io_uop_stale_pdst : _GEN_141 ? _slots_8_io_uop_stale_pdst : _GEN_135 ? _slots_7_io_uop_stale_pdst : _GEN_129 ? _slots_6_io_uop_stale_pdst : _GEN_123 ? _slots_5_io_uop_stale_pdst : _GEN_117 ? _slots_4_io_uop_stale_pdst : _GEN_111 ? _slots_3_io_uop_stale_pdst : _GEN_105 ? _slots_2_io_uop_stale_pdst : _GEN_99 ? _slots_1_io_uop_stale_pdst : _GEN_94 ? _slots_0_io_uop_stale_pdst : 7'h0;
  assign io_iss_uops_1_exception = _GEN_226 ? _slots_23_io_uop_exception : _GEN_224 ? _slots_22_io_uop_exception : _GEN_219 ? _slots_21_io_uop_exception : _GEN_213 ? _slots_20_io_uop_exception : _GEN_207 ? _slots_19_io_uop_exception : _GEN_201 ? _slots_18_io_uop_exception : _GEN_195 ? _slots_17_io_uop_exception : _GEN_189 ? _slots_16_io_uop_exception : _GEN_183 ? _slots_15_io_uop_exception : _GEN_177 ? _slots_14_io_uop_exception : _GEN_171 ? _slots_13_io_uop_exception : _GEN_165 ? _slots_12_io_uop_exception : _GEN_159 ? _slots_11_io_uop_exception : _GEN_153 ? _slots_10_io_uop_exception : _GEN_147 ? _slots_9_io_uop_exception : _GEN_141 ? _slots_8_io_uop_exception : _GEN_135 ? _slots_7_io_uop_exception : _GEN_129 ? _slots_6_io_uop_exception : _GEN_123 ? _slots_5_io_uop_exception : _GEN_117 ? _slots_4_io_uop_exception : _GEN_111 ? _slots_3_io_uop_exception : _GEN_105 ? _slots_2_io_uop_exception : _GEN_99 ? _slots_1_io_uop_exception : _GEN_94 & _slots_0_io_uop_exception;
  assign io_iss_uops_1_exc_cause = _GEN_226 ? _slots_23_io_uop_exc_cause : _GEN_224 ? _slots_22_io_uop_exc_cause : _GEN_219 ? _slots_21_io_uop_exc_cause : _GEN_213 ? _slots_20_io_uop_exc_cause : _GEN_207 ? _slots_19_io_uop_exc_cause : _GEN_201 ? _slots_18_io_uop_exc_cause : _GEN_195 ? _slots_17_io_uop_exc_cause : _GEN_189 ? _slots_16_io_uop_exc_cause : _GEN_183 ? _slots_15_io_uop_exc_cause : _GEN_177 ? _slots_14_io_uop_exc_cause : _GEN_171 ? _slots_13_io_uop_exc_cause : _GEN_165 ? _slots_12_io_uop_exc_cause : _GEN_159 ? _slots_11_io_uop_exc_cause : _GEN_153 ? _slots_10_io_uop_exc_cause : _GEN_147 ? _slots_9_io_uop_exc_cause : _GEN_141 ? _slots_8_io_uop_exc_cause : _GEN_135 ? _slots_7_io_uop_exc_cause : _GEN_129 ? _slots_6_io_uop_exc_cause : _GEN_123 ? _slots_5_io_uop_exc_cause : _GEN_117 ? _slots_4_io_uop_exc_cause : _GEN_111 ? _slots_3_io_uop_exc_cause : _GEN_105 ? _slots_2_io_uop_exc_cause : _GEN_99 ? _slots_1_io_uop_exc_cause : _GEN_94 ? _slots_0_io_uop_exc_cause : 64'h0;
  assign io_iss_uops_1_bypassable = _GEN_226 ? _slots_23_io_uop_bypassable : _GEN_224 ? _slots_22_io_uop_bypassable : _GEN_219 ? _slots_21_io_uop_bypassable : _GEN_213 ? _slots_20_io_uop_bypassable : _GEN_207 ? _slots_19_io_uop_bypassable : _GEN_201 ? _slots_18_io_uop_bypassable : _GEN_195 ? _slots_17_io_uop_bypassable : _GEN_189 ? _slots_16_io_uop_bypassable : _GEN_183 ? _slots_15_io_uop_bypassable : _GEN_177 ? _slots_14_io_uop_bypassable : _GEN_171 ? _slots_13_io_uop_bypassable : _GEN_165 ? _slots_12_io_uop_bypassable : _GEN_159 ? _slots_11_io_uop_bypassable : _GEN_153 ? _slots_10_io_uop_bypassable : _GEN_147 ? _slots_9_io_uop_bypassable : _GEN_141 ? _slots_8_io_uop_bypassable : _GEN_135 ? _slots_7_io_uop_bypassable : _GEN_129 ? _slots_6_io_uop_bypassable : _GEN_123 ? _slots_5_io_uop_bypassable : _GEN_117 ? _slots_4_io_uop_bypassable : _GEN_111 ? _slots_3_io_uop_bypassable : _GEN_105 ? _slots_2_io_uop_bypassable : _GEN_99 ? _slots_1_io_uop_bypassable : _GEN_94 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_1_mem_cmd = _GEN_226 ? _slots_23_io_uop_mem_cmd : _GEN_224 ? _slots_22_io_uop_mem_cmd : _GEN_219 ? _slots_21_io_uop_mem_cmd : _GEN_213 ? _slots_20_io_uop_mem_cmd : _GEN_207 ? _slots_19_io_uop_mem_cmd : _GEN_201 ? _slots_18_io_uop_mem_cmd : _GEN_195 ? _slots_17_io_uop_mem_cmd : _GEN_189 ? _slots_16_io_uop_mem_cmd : _GEN_183 ? _slots_15_io_uop_mem_cmd : _GEN_177 ? _slots_14_io_uop_mem_cmd : _GEN_171 ? _slots_13_io_uop_mem_cmd : _GEN_165 ? _slots_12_io_uop_mem_cmd : _GEN_159 ? _slots_11_io_uop_mem_cmd : _GEN_153 ? _slots_10_io_uop_mem_cmd : _GEN_147 ? _slots_9_io_uop_mem_cmd : _GEN_141 ? _slots_8_io_uop_mem_cmd : _GEN_135 ? _slots_7_io_uop_mem_cmd : _GEN_129 ? _slots_6_io_uop_mem_cmd : _GEN_123 ? _slots_5_io_uop_mem_cmd : _GEN_117 ? _slots_4_io_uop_mem_cmd : _GEN_111 ? _slots_3_io_uop_mem_cmd : _GEN_105 ? _slots_2_io_uop_mem_cmd : _GEN_99 ? _slots_1_io_uop_mem_cmd : _GEN_94 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_1_mem_size = _GEN_226 ? _slots_23_io_uop_mem_size : _GEN_224 ? _slots_22_io_uop_mem_size : _GEN_219 ? _slots_21_io_uop_mem_size : _GEN_213 ? _slots_20_io_uop_mem_size : _GEN_207 ? _slots_19_io_uop_mem_size : _GEN_201 ? _slots_18_io_uop_mem_size : _GEN_195 ? _slots_17_io_uop_mem_size : _GEN_189 ? _slots_16_io_uop_mem_size : _GEN_183 ? _slots_15_io_uop_mem_size : _GEN_177 ? _slots_14_io_uop_mem_size : _GEN_171 ? _slots_13_io_uop_mem_size : _GEN_165 ? _slots_12_io_uop_mem_size : _GEN_159 ? _slots_11_io_uop_mem_size : _GEN_153 ? _slots_10_io_uop_mem_size : _GEN_147 ? _slots_9_io_uop_mem_size : _GEN_141 ? _slots_8_io_uop_mem_size : _GEN_135 ? _slots_7_io_uop_mem_size : _GEN_129 ? _slots_6_io_uop_mem_size : _GEN_123 ? _slots_5_io_uop_mem_size : _GEN_117 ? _slots_4_io_uop_mem_size : _GEN_111 ? _slots_3_io_uop_mem_size : _GEN_105 ? _slots_2_io_uop_mem_size : _GEN_99 ? _slots_1_io_uop_mem_size : _GEN_94 ? _slots_0_io_uop_mem_size : 2'h0;
  assign io_iss_uops_1_mem_signed = _GEN_226 ? _slots_23_io_uop_mem_signed : _GEN_224 ? _slots_22_io_uop_mem_signed : _GEN_219 ? _slots_21_io_uop_mem_signed : _GEN_213 ? _slots_20_io_uop_mem_signed : _GEN_207 ? _slots_19_io_uop_mem_signed : _GEN_201 ? _slots_18_io_uop_mem_signed : _GEN_195 ? _slots_17_io_uop_mem_signed : _GEN_189 ? _slots_16_io_uop_mem_signed : _GEN_183 ? _slots_15_io_uop_mem_signed : _GEN_177 ? _slots_14_io_uop_mem_signed : _GEN_171 ? _slots_13_io_uop_mem_signed : _GEN_165 ? _slots_12_io_uop_mem_signed : _GEN_159 ? _slots_11_io_uop_mem_signed : _GEN_153 ? _slots_10_io_uop_mem_signed : _GEN_147 ? _slots_9_io_uop_mem_signed : _GEN_141 ? _slots_8_io_uop_mem_signed : _GEN_135 ? _slots_7_io_uop_mem_signed : _GEN_129 ? _slots_6_io_uop_mem_signed : _GEN_123 ? _slots_5_io_uop_mem_signed : _GEN_117 ? _slots_4_io_uop_mem_signed : _GEN_111 ? _slots_3_io_uop_mem_signed : _GEN_105 ? _slots_2_io_uop_mem_signed : _GEN_99 ? _slots_1_io_uop_mem_signed : _GEN_94 & _slots_0_io_uop_mem_signed;
  assign io_iss_uops_1_is_fence = _GEN_226 ? _slots_23_io_uop_is_fence : _GEN_224 ? _slots_22_io_uop_is_fence : _GEN_219 ? _slots_21_io_uop_is_fence : _GEN_213 ? _slots_20_io_uop_is_fence : _GEN_207 ? _slots_19_io_uop_is_fence : _GEN_201 ? _slots_18_io_uop_is_fence : _GEN_195 ? _slots_17_io_uop_is_fence : _GEN_189 ? _slots_16_io_uop_is_fence : _GEN_183 ? _slots_15_io_uop_is_fence : _GEN_177 ? _slots_14_io_uop_is_fence : _GEN_171 ? _slots_13_io_uop_is_fence : _GEN_165 ? _slots_12_io_uop_is_fence : _GEN_159 ? _slots_11_io_uop_is_fence : _GEN_153 ? _slots_10_io_uop_is_fence : _GEN_147 ? _slots_9_io_uop_is_fence : _GEN_141 ? _slots_8_io_uop_is_fence : _GEN_135 ? _slots_7_io_uop_is_fence : _GEN_129 ? _slots_6_io_uop_is_fence : _GEN_123 ? _slots_5_io_uop_is_fence : _GEN_117 ? _slots_4_io_uop_is_fence : _GEN_111 ? _slots_3_io_uop_is_fence : _GEN_105 ? _slots_2_io_uop_is_fence : _GEN_99 ? _slots_1_io_uop_is_fence : _GEN_94 & _slots_0_io_uop_is_fence;
  assign io_iss_uops_1_is_fencei = _GEN_226 ? _slots_23_io_uop_is_fencei : _GEN_224 ? _slots_22_io_uop_is_fencei : _GEN_219 ? _slots_21_io_uop_is_fencei : _GEN_213 ? _slots_20_io_uop_is_fencei : _GEN_207 ? _slots_19_io_uop_is_fencei : _GEN_201 ? _slots_18_io_uop_is_fencei : _GEN_195 ? _slots_17_io_uop_is_fencei : _GEN_189 ? _slots_16_io_uop_is_fencei : _GEN_183 ? _slots_15_io_uop_is_fencei : _GEN_177 ? _slots_14_io_uop_is_fencei : _GEN_171 ? _slots_13_io_uop_is_fencei : _GEN_165 ? _slots_12_io_uop_is_fencei : _GEN_159 ? _slots_11_io_uop_is_fencei : _GEN_153 ? _slots_10_io_uop_is_fencei : _GEN_147 ? _slots_9_io_uop_is_fencei : _GEN_141 ? _slots_8_io_uop_is_fencei : _GEN_135 ? _slots_7_io_uop_is_fencei : _GEN_129 ? _slots_6_io_uop_is_fencei : _GEN_123 ? _slots_5_io_uop_is_fencei : _GEN_117 ? _slots_4_io_uop_is_fencei : _GEN_111 ? _slots_3_io_uop_is_fencei : _GEN_105 ? _slots_2_io_uop_is_fencei : _GEN_99 ? _slots_1_io_uop_is_fencei : _GEN_94 & _slots_0_io_uop_is_fencei;
  assign io_iss_uops_1_is_amo = _GEN_226 ? _slots_23_io_uop_is_amo : _GEN_224 ? _slots_22_io_uop_is_amo : _GEN_219 ? _slots_21_io_uop_is_amo : _GEN_213 ? _slots_20_io_uop_is_amo : _GEN_207 ? _slots_19_io_uop_is_amo : _GEN_201 ? _slots_18_io_uop_is_amo : _GEN_195 ? _slots_17_io_uop_is_amo : _GEN_189 ? _slots_16_io_uop_is_amo : _GEN_183 ? _slots_15_io_uop_is_amo : _GEN_177 ? _slots_14_io_uop_is_amo : _GEN_171 ? _slots_13_io_uop_is_amo : _GEN_165 ? _slots_12_io_uop_is_amo : _GEN_159 ? _slots_11_io_uop_is_amo : _GEN_153 ? _slots_10_io_uop_is_amo : _GEN_147 ? _slots_9_io_uop_is_amo : _GEN_141 ? _slots_8_io_uop_is_amo : _GEN_135 ? _slots_7_io_uop_is_amo : _GEN_129 ? _slots_6_io_uop_is_amo : _GEN_123 ? _slots_5_io_uop_is_amo : _GEN_117 ? _slots_4_io_uop_is_amo : _GEN_111 ? _slots_3_io_uop_is_amo : _GEN_105 ? _slots_2_io_uop_is_amo : _GEN_99 ? _slots_1_io_uop_is_amo : _GEN_94 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_1_uses_ldq = _GEN_226 ? _slots_23_io_uop_uses_ldq : _GEN_224 ? _slots_22_io_uop_uses_ldq : _GEN_219 ? _slots_21_io_uop_uses_ldq : _GEN_213 ? _slots_20_io_uop_uses_ldq : _GEN_207 ? _slots_19_io_uop_uses_ldq : _GEN_201 ? _slots_18_io_uop_uses_ldq : _GEN_195 ? _slots_17_io_uop_uses_ldq : _GEN_189 ? _slots_16_io_uop_uses_ldq : _GEN_183 ? _slots_15_io_uop_uses_ldq : _GEN_177 ? _slots_14_io_uop_uses_ldq : _GEN_171 ? _slots_13_io_uop_uses_ldq : _GEN_165 ? _slots_12_io_uop_uses_ldq : _GEN_159 ? _slots_11_io_uop_uses_ldq : _GEN_153 ? _slots_10_io_uop_uses_ldq : _GEN_147 ? _slots_9_io_uop_uses_ldq : _GEN_141 ? _slots_8_io_uop_uses_ldq : _GEN_135 ? _slots_7_io_uop_uses_ldq : _GEN_129 ? _slots_6_io_uop_uses_ldq : _GEN_123 ? _slots_5_io_uop_uses_ldq : _GEN_117 ? _slots_4_io_uop_uses_ldq : _GEN_111 ? _slots_3_io_uop_uses_ldq : _GEN_105 ? _slots_2_io_uop_uses_ldq : _GEN_99 ? _slots_1_io_uop_uses_ldq : _GEN_94 & _slots_0_io_uop_uses_ldq;
  assign io_iss_uops_1_uses_stq = _GEN_226 ? _slots_23_io_uop_uses_stq : _GEN_224 ? _slots_22_io_uop_uses_stq : _GEN_219 ? _slots_21_io_uop_uses_stq : _GEN_213 ? _slots_20_io_uop_uses_stq : _GEN_207 ? _slots_19_io_uop_uses_stq : _GEN_201 ? _slots_18_io_uop_uses_stq : _GEN_195 ? _slots_17_io_uop_uses_stq : _GEN_189 ? _slots_16_io_uop_uses_stq : _GEN_183 ? _slots_15_io_uop_uses_stq : _GEN_177 ? _slots_14_io_uop_uses_stq : _GEN_171 ? _slots_13_io_uop_uses_stq : _GEN_165 ? _slots_12_io_uop_uses_stq : _GEN_159 ? _slots_11_io_uop_uses_stq : _GEN_153 ? _slots_10_io_uop_uses_stq : _GEN_147 ? _slots_9_io_uop_uses_stq : _GEN_141 ? _slots_8_io_uop_uses_stq : _GEN_135 ? _slots_7_io_uop_uses_stq : _GEN_129 ? _slots_6_io_uop_uses_stq : _GEN_123 ? _slots_5_io_uop_uses_stq : _GEN_117 ? _slots_4_io_uop_uses_stq : _GEN_111 ? _slots_3_io_uop_uses_stq : _GEN_105 ? _slots_2_io_uop_uses_stq : _GEN_99 ? _slots_1_io_uop_uses_stq : _GEN_94 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_1_is_sys_pc2epc = _GEN_226 ? _slots_23_io_uop_is_sys_pc2epc : _GEN_224 ? _slots_22_io_uop_is_sys_pc2epc : _GEN_219 ? _slots_21_io_uop_is_sys_pc2epc : _GEN_213 ? _slots_20_io_uop_is_sys_pc2epc : _GEN_207 ? _slots_19_io_uop_is_sys_pc2epc : _GEN_201 ? _slots_18_io_uop_is_sys_pc2epc : _GEN_195 ? _slots_17_io_uop_is_sys_pc2epc : _GEN_189 ? _slots_16_io_uop_is_sys_pc2epc : _GEN_183 ? _slots_15_io_uop_is_sys_pc2epc : _GEN_177 ? _slots_14_io_uop_is_sys_pc2epc : _GEN_171 ? _slots_13_io_uop_is_sys_pc2epc : _GEN_165 ? _slots_12_io_uop_is_sys_pc2epc : _GEN_159 ? _slots_11_io_uop_is_sys_pc2epc : _GEN_153 ? _slots_10_io_uop_is_sys_pc2epc : _GEN_147 ? _slots_9_io_uop_is_sys_pc2epc : _GEN_141 ? _slots_8_io_uop_is_sys_pc2epc : _GEN_135 ? _slots_7_io_uop_is_sys_pc2epc : _GEN_129 ? _slots_6_io_uop_is_sys_pc2epc : _GEN_123 ? _slots_5_io_uop_is_sys_pc2epc : _GEN_117 ? _slots_4_io_uop_is_sys_pc2epc : _GEN_111 ? _slots_3_io_uop_is_sys_pc2epc : _GEN_105 ? _slots_2_io_uop_is_sys_pc2epc : _GEN_99 ? _slots_1_io_uop_is_sys_pc2epc : _GEN_94 & _slots_0_io_uop_is_sys_pc2epc;
  assign io_iss_uops_1_is_unique = _GEN_226 ? _slots_23_io_uop_is_unique : _GEN_224 ? _slots_22_io_uop_is_unique : _GEN_219 ? _slots_21_io_uop_is_unique : _GEN_213 ? _slots_20_io_uop_is_unique : _GEN_207 ? _slots_19_io_uop_is_unique : _GEN_201 ? _slots_18_io_uop_is_unique : _GEN_195 ? _slots_17_io_uop_is_unique : _GEN_189 ? _slots_16_io_uop_is_unique : _GEN_183 ? _slots_15_io_uop_is_unique : _GEN_177 ? _slots_14_io_uop_is_unique : _GEN_171 ? _slots_13_io_uop_is_unique : _GEN_165 ? _slots_12_io_uop_is_unique : _GEN_159 ? _slots_11_io_uop_is_unique : _GEN_153 ? _slots_10_io_uop_is_unique : _GEN_147 ? _slots_9_io_uop_is_unique : _GEN_141 ? _slots_8_io_uop_is_unique : _GEN_135 ? _slots_7_io_uop_is_unique : _GEN_129 ? _slots_6_io_uop_is_unique : _GEN_123 ? _slots_5_io_uop_is_unique : _GEN_117 ? _slots_4_io_uop_is_unique : _GEN_111 ? _slots_3_io_uop_is_unique : _GEN_105 ? _slots_2_io_uop_is_unique : _GEN_99 ? _slots_1_io_uop_is_unique : _GEN_94 & _slots_0_io_uop_is_unique;
  assign io_iss_uops_1_flush_on_commit = _GEN_226 ? _slots_23_io_uop_flush_on_commit : _GEN_224 ? _slots_22_io_uop_flush_on_commit : _GEN_219 ? _slots_21_io_uop_flush_on_commit : _GEN_213 ? _slots_20_io_uop_flush_on_commit : _GEN_207 ? _slots_19_io_uop_flush_on_commit : _GEN_201 ? _slots_18_io_uop_flush_on_commit : _GEN_195 ? _slots_17_io_uop_flush_on_commit : _GEN_189 ? _slots_16_io_uop_flush_on_commit : _GEN_183 ? _slots_15_io_uop_flush_on_commit : _GEN_177 ? _slots_14_io_uop_flush_on_commit : _GEN_171 ? _slots_13_io_uop_flush_on_commit : _GEN_165 ? _slots_12_io_uop_flush_on_commit : _GEN_159 ? _slots_11_io_uop_flush_on_commit : _GEN_153 ? _slots_10_io_uop_flush_on_commit : _GEN_147 ? _slots_9_io_uop_flush_on_commit : _GEN_141 ? _slots_8_io_uop_flush_on_commit : _GEN_135 ? _slots_7_io_uop_flush_on_commit : _GEN_129 ? _slots_6_io_uop_flush_on_commit : _GEN_123 ? _slots_5_io_uop_flush_on_commit : _GEN_117 ? _slots_4_io_uop_flush_on_commit : _GEN_111 ? _slots_3_io_uop_flush_on_commit : _GEN_105 ? _slots_2_io_uop_flush_on_commit : _GEN_99 ? _slots_1_io_uop_flush_on_commit : _GEN_94 & _slots_0_io_uop_flush_on_commit;
  assign io_iss_uops_1_ldst_is_rs1 = _GEN_226 ? _slots_23_io_uop_ldst_is_rs1 : _GEN_224 ? _slots_22_io_uop_ldst_is_rs1 : _GEN_219 ? _slots_21_io_uop_ldst_is_rs1 : _GEN_213 ? _slots_20_io_uop_ldst_is_rs1 : _GEN_207 ? _slots_19_io_uop_ldst_is_rs1 : _GEN_201 ? _slots_18_io_uop_ldst_is_rs1 : _GEN_195 ? _slots_17_io_uop_ldst_is_rs1 : _GEN_189 ? _slots_16_io_uop_ldst_is_rs1 : _GEN_183 ? _slots_15_io_uop_ldst_is_rs1 : _GEN_177 ? _slots_14_io_uop_ldst_is_rs1 : _GEN_171 ? _slots_13_io_uop_ldst_is_rs1 : _GEN_165 ? _slots_12_io_uop_ldst_is_rs1 : _GEN_159 ? _slots_11_io_uop_ldst_is_rs1 : _GEN_153 ? _slots_10_io_uop_ldst_is_rs1 : _GEN_147 ? _slots_9_io_uop_ldst_is_rs1 : _GEN_141 ? _slots_8_io_uop_ldst_is_rs1 : _GEN_135 ? _slots_7_io_uop_ldst_is_rs1 : _GEN_129 ? _slots_6_io_uop_ldst_is_rs1 : _GEN_123 ? _slots_5_io_uop_ldst_is_rs1 : _GEN_117 ? _slots_4_io_uop_ldst_is_rs1 : _GEN_111 ? _slots_3_io_uop_ldst_is_rs1 : _GEN_105 ? _slots_2_io_uop_ldst_is_rs1 : _GEN_99 ? _slots_1_io_uop_ldst_is_rs1 : _GEN_94 & _slots_0_io_uop_ldst_is_rs1;
  assign io_iss_uops_1_ldst = _GEN_226 ? _slots_23_io_uop_ldst : _GEN_224 ? _slots_22_io_uop_ldst : _GEN_219 ? _slots_21_io_uop_ldst : _GEN_213 ? _slots_20_io_uop_ldst : _GEN_207 ? _slots_19_io_uop_ldst : _GEN_201 ? _slots_18_io_uop_ldst : _GEN_195 ? _slots_17_io_uop_ldst : _GEN_189 ? _slots_16_io_uop_ldst : _GEN_183 ? _slots_15_io_uop_ldst : _GEN_177 ? _slots_14_io_uop_ldst : _GEN_171 ? _slots_13_io_uop_ldst : _GEN_165 ? _slots_12_io_uop_ldst : _GEN_159 ? _slots_11_io_uop_ldst : _GEN_153 ? _slots_10_io_uop_ldst : _GEN_147 ? _slots_9_io_uop_ldst : _GEN_141 ? _slots_8_io_uop_ldst : _GEN_135 ? _slots_7_io_uop_ldst : _GEN_129 ? _slots_6_io_uop_ldst : _GEN_123 ? _slots_5_io_uop_ldst : _GEN_117 ? _slots_4_io_uop_ldst : _GEN_111 ? _slots_3_io_uop_ldst : _GEN_105 ? _slots_2_io_uop_ldst : _GEN_99 ? _slots_1_io_uop_ldst : _GEN_94 ? _slots_0_io_uop_ldst : 6'h0;
  assign io_iss_uops_1_lrs1 = _GEN_226 ? _slots_23_io_uop_lrs1 : _GEN_224 ? _slots_22_io_uop_lrs1 : _GEN_219 ? _slots_21_io_uop_lrs1 : _GEN_213 ? _slots_20_io_uop_lrs1 : _GEN_207 ? _slots_19_io_uop_lrs1 : _GEN_201 ? _slots_18_io_uop_lrs1 : _GEN_195 ? _slots_17_io_uop_lrs1 : _GEN_189 ? _slots_16_io_uop_lrs1 : _GEN_183 ? _slots_15_io_uop_lrs1 : _GEN_177 ? _slots_14_io_uop_lrs1 : _GEN_171 ? _slots_13_io_uop_lrs1 : _GEN_165 ? _slots_12_io_uop_lrs1 : _GEN_159 ? _slots_11_io_uop_lrs1 : _GEN_153 ? _slots_10_io_uop_lrs1 : _GEN_147 ? _slots_9_io_uop_lrs1 : _GEN_141 ? _slots_8_io_uop_lrs1 : _GEN_135 ? _slots_7_io_uop_lrs1 : _GEN_129 ? _slots_6_io_uop_lrs1 : _GEN_123 ? _slots_5_io_uop_lrs1 : _GEN_117 ? _slots_4_io_uop_lrs1 : _GEN_111 ? _slots_3_io_uop_lrs1 : _GEN_105 ? _slots_2_io_uop_lrs1 : _GEN_99 ? _slots_1_io_uop_lrs1 : _GEN_94 ? _slots_0_io_uop_lrs1 : 6'h0;
  assign io_iss_uops_1_lrs2 = _GEN_226 ? _slots_23_io_uop_lrs2 : _GEN_224 ? _slots_22_io_uop_lrs2 : _GEN_219 ? _slots_21_io_uop_lrs2 : _GEN_213 ? _slots_20_io_uop_lrs2 : _GEN_207 ? _slots_19_io_uop_lrs2 : _GEN_201 ? _slots_18_io_uop_lrs2 : _GEN_195 ? _slots_17_io_uop_lrs2 : _GEN_189 ? _slots_16_io_uop_lrs2 : _GEN_183 ? _slots_15_io_uop_lrs2 : _GEN_177 ? _slots_14_io_uop_lrs2 : _GEN_171 ? _slots_13_io_uop_lrs2 : _GEN_165 ? _slots_12_io_uop_lrs2 : _GEN_159 ? _slots_11_io_uop_lrs2 : _GEN_153 ? _slots_10_io_uop_lrs2 : _GEN_147 ? _slots_9_io_uop_lrs2 : _GEN_141 ? _slots_8_io_uop_lrs2 : _GEN_135 ? _slots_7_io_uop_lrs2 : _GEN_129 ? _slots_6_io_uop_lrs2 : _GEN_123 ? _slots_5_io_uop_lrs2 : _GEN_117 ? _slots_4_io_uop_lrs2 : _GEN_111 ? _slots_3_io_uop_lrs2 : _GEN_105 ? _slots_2_io_uop_lrs2 : _GEN_99 ? _slots_1_io_uop_lrs2 : _GEN_94 ? _slots_0_io_uop_lrs2 : 6'h0;
  assign io_iss_uops_1_lrs3 = _GEN_226 ? _slots_23_io_uop_lrs3 : _GEN_224 ? _slots_22_io_uop_lrs3 : _GEN_219 ? _slots_21_io_uop_lrs3 : _GEN_213 ? _slots_20_io_uop_lrs3 : _GEN_207 ? _slots_19_io_uop_lrs3 : _GEN_201 ? _slots_18_io_uop_lrs3 : _GEN_195 ? _slots_17_io_uop_lrs3 : _GEN_189 ? _slots_16_io_uop_lrs3 : _GEN_183 ? _slots_15_io_uop_lrs3 : _GEN_177 ? _slots_14_io_uop_lrs3 : _GEN_171 ? _slots_13_io_uop_lrs3 : _GEN_165 ? _slots_12_io_uop_lrs3 : _GEN_159 ? _slots_11_io_uop_lrs3 : _GEN_153 ? _slots_10_io_uop_lrs3 : _GEN_147 ? _slots_9_io_uop_lrs3 : _GEN_141 ? _slots_8_io_uop_lrs3 : _GEN_135 ? _slots_7_io_uop_lrs3 : _GEN_129 ? _slots_6_io_uop_lrs3 : _GEN_123 ? _slots_5_io_uop_lrs3 : _GEN_117 ? _slots_4_io_uop_lrs3 : _GEN_111 ? _slots_3_io_uop_lrs3 : _GEN_105 ? _slots_2_io_uop_lrs3 : _GEN_99 ? _slots_1_io_uop_lrs3 : _GEN_94 ? _slots_0_io_uop_lrs3 : 6'h0;
  assign io_iss_uops_1_ldst_val = _GEN_226 ? _slots_23_io_uop_ldst_val : _GEN_224 ? _slots_22_io_uop_ldst_val : _GEN_219 ? _slots_21_io_uop_ldst_val : _GEN_213 ? _slots_20_io_uop_ldst_val : _GEN_207 ? _slots_19_io_uop_ldst_val : _GEN_201 ? _slots_18_io_uop_ldst_val : _GEN_195 ? _slots_17_io_uop_ldst_val : _GEN_189 ? _slots_16_io_uop_ldst_val : _GEN_183 ? _slots_15_io_uop_ldst_val : _GEN_177 ? _slots_14_io_uop_ldst_val : _GEN_171 ? _slots_13_io_uop_ldst_val : _GEN_165 ? _slots_12_io_uop_ldst_val : _GEN_159 ? _slots_11_io_uop_ldst_val : _GEN_153 ? _slots_10_io_uop_ldst_val : _GEN_147 ? _slots_9_io_uop_ldst_val : _GEN_141 ? _slots_8_io_uop_ldst_val : _GEN_135 ? _slots_7_io_uop_ldst_val : _GEN_129 ? _slots_6_io_uop_ldst_val : _GEN_123 ? _slots_5_io_uop_ldst_val : _GEN_117 ? _slots_4_io_uop_ldst_val : _GEN_111 ? _slots_3_io_uop_ldst_val : _GEN_105 ? _slots_2_io_uop_ldst_val : _GEN_99 ? _slots_1_io_uop_ldst_val : _GEN_94 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_1_dst_rtype = _GEN_226 ? _slots_23_io_uop_dst_rtype : _GEN_224 ? _slots_22_io_uop_dst_rtype : _GEN_219 ? _slots_21_io_uop_dst_rtype : _GEN_213 ? _slots_20_io_uop_dst_rtype : _GEN_207 ? _slots_19_io_uop_dst_rtype : _GEN_201 ? _slots_18_io_uop_dst_rtype : _GEN_195 ? _slots_17_io_uop_dst_rtype : _GEN_189 ? _slots_16_io_uop_dst_rtype : _GEN_183 ? _slots_15_io_uop_dst_rtype : _GEN_177 ? _slots_14_io_uop_dst_rtype : _GEN_171 ? _slots_13_io_uop_dst_rtype : _GEN_165 ? _slots_12_io_uop_dst_rtype : _GEN_159 ? _slots_11_io_uop_dst_rtype : _GEN_153 ? _slots_10_io_uop_dst_rtype : _GEN_147 ? _slots_9_io_uop_dst_rtype : _GEN_141 ? _slots_8_io_uop_dst_rtype : _GEN_135 ? _slots_7_io_uop_dst_rtype : _GEN_129 ? _slots_6_io_uop_dst_rtype : _GEN_123 ? _slots_5_io_uop_dst_rtype : _GEN_117 ? _slots_4_io_uop_dst_rtype : _GEN_111 ? _slots_3_io_uop_dst_rtype : _GEN_105 ? _slots_2_io_uop_dst_rtype : _GEN_99 ? _slots_1_io_uop_dst_rtype : _GEN_94 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_1_lrs1_rtype = _GEN_226 ? _slots_23_io_uop_lrs1_rtype : _GEN_224 ? _slots_22_io_uop_lrs1_rtype : _GEN_219 ? _slots_21_io_uop_lrs1_rtype : _GEN_213 ? _slots_20_io_uop_lrs1_rtype : _GEN_207 ? _slots_19_io_uop_lrs1_rtype : _GEN_201 ? _slots_18_io_uop_lrs1_rtype : _GEN_195 ? _slots_17_io_uop_lrs1_rtype : _GEN_189 ? _slots_16_io_uop_lrs1_rtype : _GEN_183 ? _slots_15_io_uop_lrs1_rtype : _GEN_177 ? _slots_14_io_uop_lrs1_rtype : _GEN_171 ? _slots_13_io_uop_lrs1_rtype : _GEN_165 ? _slots_12_io_uop_lrs1_rtype : _GEN_159 ? _slots_11_io_uop_lrs1_rtype : _GEN_153 ? _slots_10_io_uop_lrs1_rtype : _GEN_147 ? _slots_9_io_uop_lrs1_rtype : _GEN_141 ? _slots_8_io_uop_lrs1_rtype : _GEN_135 ? _slots_7_io_uop_lrs1_rtype : _GEN_129 ? _slots_6_io_uop_lrs1_rtype : _GEN_123 ? _slots_5_io_uop_lrs1_rtype : _GEN_117 ? _slots_4_io_uop_lrs1_rtype : _GEN_111 ? _slots_3_io_uop_lrs1_rtype : _GEN_105 ? _slots_2_io_uop_lrs1_rtype : _GEN_99 ? _slots_1_io_uop_lrs1_rtype : _GEN_94 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_1_lrs2_rtype = _GEN_226 ? _slots_23_io_uop_lrs2_rtype : _GEN_224 ? _slots_22_io_uop_lrs2_rtype : _GEN_219 ? _slots_21_io_uop_lrs2_rtype : _GEN_213 ? _slots_20_io_uop_lrs2_rtype : _GEN_207 ? _slots_19_io_uop_lrs2_rtype : _GEN_201 ? _slots_18_io_uop_lrs2_rtype : _GEN_195 ? _slots_17_io_uop_lrs2_rtype : _GEN_189 ? _slots_16_io_uop_lrs2_rtype : _GEN_183 ? _slots_15_io_uop_lrs2_rtype : _GEN_177 ? _slots_14_io_uop_lrs2_rtype : _GEN_171 ? _slots_13_io_uop_lrs2_rtype : _GEN_165 ? _slots_12_io_uop_lrs2_rtype : _GEN_159 ? _slots_11_io_uop_lrs2_rtype : _GEN_153 ? _slots_10_io_uop_lrs2_rtype : _GEN_147 ? _slots_9_io_uop_lrs2_rtype : _GEN_141 ? _slots_8_io_uop_lrs2_rtype : _GEN_135 ? _slots_7_io_uop_lrs2_rtype : _GEN_129 ? _slots_6_io_uop_lrs2_rtype : _GEN_123 ? _slots_5_io_uop_lrs2_rtype : _GEN_117 ? _slots_4_io_uop_lrs2_rtype : _GEN_111 ? _slots_3_io_uop_lrs2_rtype : _GEN_105 ? _slots_2_io_uop_lrs2_rtype : _GEN_99 ? _slots_1_io_uop_lrs2_rtype : _GEN_94 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_1_frs3_en = _GEN_226 ? _slots_23_io_uop_frs3_en : _GEN_224 ? _slots_22_io_uop_frs3_en : _GEN_219 ? _slots_21_io_uop_frs3_en : _GEN_213 ? _slots_20_io_uop_frs3_en : _GEN_207 ? _slots_19_io_uop_frs3_en : _GEN_201 ? _slots_18_io_uop_frs3_en : _GEN_195 ? _slots_17_io_uop_frs3_en : _GEN_189 ? _slots_16_io_uop_frs3_en : _GEN_183 ? _slots_15_io_uop_frs3_en : _GEN_177 ? _slots_14_io_uop_frs3_en : _GEN_171 ? _slots_13_io_uop_frs3_en : _GEN_165 ? _slots_12_io_uop_frs3_en : _GEN_159 ? _slots_11_io_uop_frs3_en : _GEN_153 ? _slots_10_io_uop_frs3_en : _GEN_147 ? _slots_9_io_uop_frs3_en : _GEN_141 ? _slots_8_io_uop_frs3_en : _GEN_135 ? _slots_7_io_uop_frs3_en : _GEN_129 ? _slots_6_io_uop_frs3_en : _GEN_123 ? _slots_5_io_uop_frs3_en : _GEN_117 ? _slots_4_io_uop_frs3_en : _GEN_111 ? _slots_3_io_uop_frs3_en : _GEN_105 ? _slots_2_io_uop_frs3_en : _GEN_99 ? _slots_1_io_uop_frs3_en : _GEN_94 & _slots_0_io_uop_frs3_en;
  assign io_iss_uops_1_fp_val = _GEN_226 ? _slots_23_io_uop_fp_val : _GEN_224 ? _slots_22_io_uop_fp_val : _GEN_219 ? _slots_21_io_uop_fp_val : _GEN_213 ? _slots_20_io_uop_fp_val : _GEN_207 ? _slots_19_io_uop_fp_val : _GEN_201 ? _slots_18_io_uop_fp_val : _GEN_195 ? _slots_17_io_uop_fp_val : _GEN_189 ? _slots_16_io_uop_fp_val : _GEN_183 ? _slots_15_io_uop_fp_val : _GEN_177 ? _slots_14_io_uop_fp_val : _GEN_171 ? _slots_13_io_uop_fp_val : _GEN_165 ? _slots_12_io_uop_fp_val : _GEN_159 ? _slots_11_io_uop_fp_val : _GEN_153 ? _slots_10_io_uop_fp_val : _GEN_147 ? _slots_9_io_uop_fp_val : _GEN_141 ? _slots_8_io_uop_fp_val : _GEN_135 ? _slots_7_io_uop_fp_val : _GEN_129 ? _slots_6_io_uop_fp_val : _GEN_123 ? _slots_5_io_uop_fp_val : _GEN_117 ? _slots_4_io_uop_fp_val : _GEN_111 ? _slots_3_io_uop_fp_val : _GEN_105 ? _slots_2_io_uop_fp_val : _GEN_99 ? _slots_1_io_uop_fp_val : _GEN_94 & _slots_0_io_uop_fp_val;
  assign io_iss_uops_1_fp_single = _GEN_226 ? _slots_23_io_uop_fp_single : _GEN_224 ? _slots_22_io_uop_fp_single : _GEN_219 ? _slots_21_io_uop_fp_single : _GEN_213 ? _slots_20_io_uop_fp_single : _GEN_207 ? _slots_19_io_uop_fp_single : _GEN_201 ? _slots_18_io_uop_fp_single : _GEN_195 ? _slots_17_io_uop_fp_single : _GEN_189 ? _slots_16_io_uop_fp_single : _GEN_183 ? _slots_15_io_uop_fp_single : _GEN_177 ? _slots_14_io_uop_fp_single : _GEN_171 ? _slots_13_io_uop_fp_single : _GEN_165 ? _slots_12_io_uop_fp_single : _GEN_159 ? _slots_11_io_uop_fp_single : _GEN_153 ? _slots_10_io_uop_fp_single : _GEN_147 ? _slots_9_io_uop_fp_single : _GEN_141 ? _slots_8_io_uop_fp_single : _GEN_135 ? _slots_7_io_uop_fp_single : _GEN_129 ? _slots_6_io_uop_fp_single : _GEN_123 ? _slots_5_io_uop_fp_single : _GEN_117 ? _slots_4_io_uop_fp_single : _GEN_111 ? _slots_3_io_uop_fp_single : _GEN_105 ? _slots_2_io_uop_fp_single : _GEN_99 ? _slots_1_io_uop_fp_single : _GEN_94 & _slots_0_io_uop_fp_single;
  assign io_iss_uops_1_xcpt_pf_if = _GEN_226 ? _slots_23_io_uop_xcpt_pf_if : _GEN_224 ? _slots_22_io_uop_xcpt_pf_if : _GEN_219 ? _slots_21_io_uop_xcpt_pf_if : _GEN_213 ? _slots_20_io_uop_xcpt_pf_if : _GEN_207 ? _slots_19_io_uop_xcpt_pf_if : _GEN_201 ? _slots_18_io_uop_xcpt_pf_if : _GEN_195 ? _slots_17_io_uop_xcpt_pf_if : _GEN_189 ? _slots_16_io_uop_xcpt_pf_if : _GEN_183 ? _slots_15_io_uop_xcpt_pf_if : _GEN_177 ? _slots_14_io_uop_xcpt_pf_if : _GEN_171 ? _slots_13_io_uop_xcpt_pf_if : _GEN_165 ? _slots_12_io_uop_xcpt_pf_if : _GEN_159 ? _slots_11_io_uop_xcpt_pf_if : _GEN_153 ? _slots_10_io_uop_xcpt_pf_if : _GEN_147 ? _slots_9_io_uop_xcpt_pf_if : _GEN_141 ? _slots_8_io_uop_xcpt_pf_if : _GEN_135 ? _slots_7_io_uop_xcpt_pf_if : _GEN_129 ? _slots_6_io_uop_xcpt_pf_if : _GEN_123 ? _slots_5_io_uop_xcpt_pf_if : _GEN_117 ? _slots_4_io_uop_xcpt_pf_if : _GEN_111 ? _slots_3_io_uop_xcpt_pf_if : _GEN_105 ? _slots_2_io_uop_xcpt_pf_if : _GEN_99 ? _slots_1_io_uop_xcpt_pf_if : _GEN_94 & _slots_0_io_uop_xcpt_pf_if;
  assign io_iss_uops_1_xcpt_ae_if = _GEN_226 ? _slots_23_io_uop_xcpt_ae_if : _GEN_224 ? _slots_22_io_uop_xcpt_ae_if : _GEN_219 ? _slots_21_io_uop_xcpt_ae_if : _GEN_213 ? _slots_20_io_uop_xcpt_ae_if : _GEN_207 ? _slots_19_io_uop_xcpt_ae_if : _GEN_201 ? _slots_18_io_uop_xcpt_ae_if : _GEN_195 ? _slots_17_io_uop_xcpt_ae_if : _GEN_189 ? _slots_16_io_uop_xcpt_ae_if : _GEN_183 ? _slots_15_io_uop_xcpt_ae_if : _GEN_177 ? _slots_14_io_uop_xcpt_ae_if : _GEN_171 ? _slots_13_io_uop_xcpt_ae_if : _GEN_165 ? _slots_12_io_uop_xcpt_ae_if : _GEN_159 ? _slots_11_io_uop_xcpt_ae_if : _GEN_153 ? _slots_10_io_uop_xcpt_ae_if : _GEN_147 ? _slots_9_io_uop_xcpt_ae_if : _GEN_141 ? _slots_8_io_uop_xcpt_ae_if : _GEN_135 ? _slots_7_io_uop_xcpt_ae_if : _GEN_129 ? _slots_6_io_uop_xcpt_ae_if : _GEN_123 ? _slots_5_io_uop_xcpt_ae_if : _GEN_117 ? _slots_4_io_uop_xcpt_ae_if : _GEN_111 ? _slots_3_io_uop_xcpt_ae_if : _GEN_105 ? _slots_2_io_uop_xcpt_ae_if : _GEN_99 ? _slots_1_io_uop_xcpt_ae_if : _GEN_94 & _slots_0_io_uop_xcpt_ae_if;
  assign io_iss_uops_1_xcpt_ma_if = _GEN_226 ? _slots_23_io_uop_xcpt_ma_if : _GEN_224 ? _slots_22_io_uop_xcpt_ma_if : _GEN_219 ? _slots_21_io_uop_xcpt_ma_if : _GEN_213 ? _slots_20_io_uop_xcpt_ma_if : _GEN_207 ? _slots_19_io_uop_xcpt_ma_if : _GEN_201 ? _slots_18_io_uop_xcpt_ma_if : _GEN_195 ? _slots_17_io_uop_xcpt_ma_if : _GEN_189 ? _slots_16_io_uop_xcpt_ma_if : _GEN_183 ? _slots_15_io_uop_xcpt_ma_if : _GEN_177 ? _slots_14_io_uop_xcpt_ma_if : _GEN_171 ? _slots_13_io_uop_xcpt_ma_if : _GEN_165 ? _slots_12_io_uop_xcpt_ma_if : _GEN_159 ? _slots_11_io_uop_xcpt_ma_if : _GEN_153 ? _slots_10_io_uop_xcpt_ma_if : _GEN_147 ? _slots_9_io_uop_xcpt_ma_if : _GEN_141 ? _slots_8_io_uop_xcpt_ma_if : _GEN_135 ? _slots_7_io_uop_xcpt_ma_if : _GEN_129 ? _slots_6_io_uop_xcpt_ma_if : _GEN_123 ? _slots_5_io_uop_xcpt_ma_if : _GEN_117 ? _slots_4_io_uop_xcpt_ma_if : _GEN_111 ? _slots_3_io_uop_xcpt_ma_if : _GEN_105 ? _slots_2_io_uop_xcpt_ma_if : _GEN_99 ? _slots_1_io_uop_xcpt_ma_if : _GEN_94 & _slots_0_io_uop_xcpt_ma_if;
  assign io_iss_uops_1_bp_debug_if = _GEN_226 ? _slots_23_io_uop_bp_debug_if : _GEN_224 ? _slots_22_io_uop_bp_debug_if : _GEN_219 ? _slots_21_io_uop_bp_debug_if : _GEN_213 ? _slots_20_io_uop_bp_debug_if : _GEN_207 ? _slots_19_io_uop_bp_debug_if : _GEN_201 ? _slots_18_io_uop_bp_debug_if : _GEN_195 ? _slots_17_io_uop_bp_debug_if : _GEN_189 ? _slots_16_io_uop_bp_debug_if : _GEN_183 ? _slots_15_io_uop_bp_debug_if : _GEN_177 ? _slots_14_io_uop_bp_debug_if : _GEN_171 ? _slots_13_io_uop_bp_debug_if : _GEN_165 ? _slots_12_io_uop_bp_debug_if : _GEN_159 ? _slots_11_io_uop_bp_debug_if : _GEN_153 ? _slots_10_io_uop_bp_debug_if : _GEN_147 ? _slots_9_io_uop_bp_debug_if : _GEN_141 ? _slots_8_io_uop_bp_debug_if : _GEN_135 ? _slots_7_io_uop_bp_debug_if : _GEN_129 ? _slots_6_io_uop_bp_debug_if : _GEN_123 ? _slots_5_io_uop_bp_debug_if : _GEN_117 ? _slots_4_io_uop_bp_debug_if : _GEN_111 ? _slots_3_io_uop_bp_debug_if : _GEN_105 ? _slots_2_io_uop_bp_debug_if : _GEN_99 ? _slots_1_io_uop_bp_debug_if : _GEN_94 & _slots_0_io_uop_bp_debug_if;
  assign io_iss_uops_1_bp_xcpt_if = _GEN_226 ? _slots_23_io_uop_bp_xcpt_if : _GEN_224 ? _slots_22_io_uop_bp_xcpt_if : _GEN_219 ? _slots_21_io_uop_bp_xcpt_if : _GEN_213 ? _slots_20_io_uop_bp_xcpt_if : _GEN_207 ? _slots_19_io_uop_bp_xcpt_if : _GEN_201 ? _slots_18_io_uop_bp_xcpt_if : _GEN_195 ? _slots_17_io_uop_bp_xcpt_if : _GEN_189 ? _slots_16_io_uop_bp_xcpt_if : _GEN_183 ? _slots_15_io_uop_bp_xcpt_if : _GEN_177 ? _slots_14_io_uop_bp_xcpt_if : _GEN_171 ? _slots_13_io_uop_bp_xcpt_if : _GEN_165 ? _slots_12_io_uop_bp_xcpt_if : _GEN_159 ? _slots_11_io_uop_bp_xcpt_if : _GEN_153 ? _slots_10_io_uop_bp_xcpt_if : _GEN_147 ? _slots_9_io_uop_bp_xcpt_if : _GEN_141 ? _slots_8_io_uop_bp_xcpt_if : _GEN_135 ? _slots_7_io_uop_bp_xcpt_if : _GEN_129 ? _slots_6_io_uop_bp_xcpt_if : _GEN_123 ? _slots_5_io_uop_bp_xcpt_if : _GEN_117 ? _slots_4_io_uop_bp_xcpt_if : _GEN_111 ? _slots_3_io_uop_bp_xcpt_if : _GEN_105 ? _slots_2_io_uop_bp_xcpt_if : _GEN_99 ? _slots_1_io_uop_bp_xcpt_if : _GEN_94 & _slots_0_io_uop_bp_xcpt_if;
  assign io_iss_uops_1_debug_fsrc = _GEN_226 ? _slots_23_io_uop_debug_fsrc : _GEN_224 ? _slots_22_io_uop_debug_fsrc : _GEN_219 ? _slots_21_io_uop_debug_fsrc : _GEN_213 ? _slots_20_io_uop_debug_fsrc : _GEN_207 ? _slots_19_io_uop_debug_fsrc : _GEN_201 ? _slots_18_io_uop_debug_fsrc : _GEN_195 ? _slots_17_io_uop_debug_fsrc : _GEN_189 ? _slots_16_io_uop_debug_fsrc : _GEN_183 ? _slots_15_io_uop_debug_fsrc : _GEN_177 ? _slots_14_io_uop_debug_fsrc : _GEN_171 ? _slots_13_io_uop_debug_fsrc : _GEN_165 ? _slots_12_io_uop_debug_fsrc : _GEN_159 ? _slots_11_io_uop_debug_fsrc : _GEN_153 ? _slots_10_io_uop_debug_fsrc : _GEN_147 ? _slots_9_io_uop_debug_fsrc : _GEN_141 ? _slots_8_io_uop_debug_fsrc : _GEN_135 ? _slots_7_io_uop_debug_fsrc : _GEN_129 ? _slots_6_io_uop_debug_fsrc : _GEN_123 ? _slots_5_io_uop_debug_fsrc : _GEN_117 ? _slots_4_io_uop_debug_fsrc : _GEN_111 ? _slots_3_io_uop_debug_fsrc : _GEN_105 ? _slots_2_io_uop_debug_fsrc : _GEN_99 ? _slots_1_io_uop_debug_fsrc : _GEN_94 ? _slots_0_io_uop_debug_fsrc : 2'h0;
  assign io_iss_uops_1_debug_tsrc = _GEN_226 ? _slots_23_io_uop_debug_tsrc : _GEN_224 ? _slots_22_io_uop_debug_tsrc : _GEN_219 ? _slots_21_io_uop_debug_tsrc : _GEN_213 ? _slots_20_io_uop_debug_tsrc : _GEN_207 ? _slots_19_io_uop_debug_tsrc : _GEN_201 ? _slots_18_io_uop_debug_tsrc : _GEN_195 ? _slots_17_io_uop_debug_tsrc : _GEN_189 ? _slots_16_io_uop_debug_tsrc : _GEN_183 ? _slots_15_io_uop_debug_tsrc : _GEN_177 ? _slots_14_io_uop_debug_tsrc : _GEN_171 ? _slots_13_io_uop_debug_tsrc : _GEN_165 ? _slots_12_io_uop_debug_tsrc : _GEN_159 ? _slots_11_io_uop_debug_tsrc : _GEN_153 ? _slots_10_io_uop_debug_tsrc : _GEN_147 ? _slots_9_io_uop_debug_tsrc : _GEN_141 ? _slots_8_io_uop_debug_tsrc : _GEN_135 ? _slots_7_io_uop_debug_tsrc : _GEN_129 ? _slots_6_io_uop_debug_tsrc : _GEN_123 ? _slots_5_io_uop_debug_tsrc : _GEN_117 ? _slots_4_io_uop_debug_tsrc : _GEN_111 ? _slots_3_io_uop_debug_tsrc : _GEN_105 ? _slots_2_io_uop_debug_tsrc : _GEN_99 ? _slots_1_io_uop_debug_tsrc : _GEN_94 ? _slots_0_io_uop_debug_tsrc : 2'h0;
endmodule

