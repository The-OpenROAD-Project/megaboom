// Standard header to adapt well known macros for prints and assertions.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module ClockDivideOrPass(
  input        io_clockIn,
  input  [7:0] io_divisor,
  input        io_resetAsync,
  output       io_clockOut
);

  wire [7:0] _divider_io_divisor_chain_io_q;
  wire       _divider_io_clockOut;
  wire       _clock_mux_io_sel_T = io_divisor == 8'h0;
  ClockDivider divider (
    .clock       (io_clockIn),
    .reset       (io_resetAsync),
    .io_divisor  (_divider_io_divisor_chain_io_q),
    .io_clockOut (_divider_io_clockOut)
  );
  SynchronizerShiftReg_w8_d3 divider_io_divisor_chain (
    .clock (io_clockIn),
    .io_d  (_clock_mux_io_sel_T ? 8'h1 : io_divisor),
    .io_q  (_divider_io_divisor_chain_io_q)
  );
  ClockMutexMux clock_mux (
    .io_clocksIn_0 (_divider_io_clockOut),
    .io_clocksIn_1 (io_clockIn),
    .io_clockOut   (io_clockOut),
    .io_resetAsync (io_resetAsync),
    .io_sel        (_clock_mux_io_sel_T)
  );
endmodule

