// Standard header to adapt well known macros for prints and assertions.

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module IssueUnitCollapsing_2(
  input         clock,
                reset,
  output        io_dis_uops_0_ready,
  input         io_dis_uops_0_valid,
  input  [6:0]  io_dis_uops_0_bits_uopc,
  input  [31:0] io_dis_uops_0_bits_inst,
                io_dis_uops_0_bits_debug_inst,
  input         io_dis_uops_0_bits_is_rvc,
  input  [39:0] io_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_dis_uops_0_bits_iq_type,
  input  [9:0]  io_dis_uops_0_bits_fu_code,
  input         io_dis_uops_0_bits_is_br,
                io_dis_uops_0_bits_is_jalr,
                io_dis_uops_0_bits_is_jal,
                io_dis_uops_0_bits_is_sfb,
  input  [19:0] io_dis_uops_0_bits_br_mask,
  input  [4:0]  io_dis_uops_0_bits_br_tag,
  input  [5:0]  io_dis_uops_0_bits_ftq_idx,
  input         io_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_dis_uops_0_bits_pc_lob,
  input         io_dis_uops_0_bits_taken,
  input  [19:0] io_dis_uops_0_bits_imm_packed,
  input  [11:0] io_dis_uops_0_bits_csr_addr,
  input  [6:0]  io_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_dis_uops_0_bits_ldq_idx,
                io_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_dis_uops_0_bits_pdst,
                io_dis_uops_0_bits_prs1,
                io_dis_uops_0_bits_prs2,
                io_dis_uops_0_bits_prs3,
  input         io_dis_uops_0_bits_prs1_busy,
                io_dis_uops_0_bits_prs2_busy,
  input  [6:0]  io_dis_uops_0_bits_stale_pdst,
  input         io_dis_uops_0_bits_exception,
  input  [63:0] io_dis_uops_0_bits_exc_cause,
  input         io_dis_uops_0_bits_bypassable,
  input  [4:0]  io_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_dis_uops_0_bits_mem_size,
  input         io_dis_uops_0_bits_mem_signed,
                io_dis_uops_0_bits_is_fence,
                io_dis_uops_0_bits_is_fencei,
                io_dis_uops_0_bits_is_amo,
                io_dis_uops_0_bits_uses_ldq,
                io_dis_uops_0_bits_uses_stq,
                io_dis_uops_0_bits_is_sys_pc2epc,
                io_dis_uops_0_bits_is_unique,
                io_dis_uops_0_bits_flush_on_commit,
                io_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_0_bits_ldst,
                io_dis_uops_0_bits_lrs1,
                io_dis_uops_0_bits_lrs2,
                io_dis_uops_0_bits_lrs3,
  input         io_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_dis_uops_0_bits_dst_rtype,
                io_dis_uops_0_bits_lrs1_rtype,
                io_dis_uops_0_bits_lrs2_rtype,
  input         io_dis_uops_0_bits_frs3_en,
                io_dis_uops_0_bits_fp_val,
                io_dis_uops_0_bits_fp_single,
                io_dis_uops_0_bits_xcpt_pf_if,
                io_dis_uops_0_bits_xcpt_ae_if,
                io_dis_uops_0_bits_xcpt_ma_if,
                io_dis_uops_0_bits_bp_debug_if,
                io_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_0_bits_debug_fsrc,
                io_dis_uops_0_bits_debug_tsrc,
  output        io_dis_uops_1_ready,
  input         io_dis_uops_1_valid,
  input  [6:0]  io_dis_uops_1_bits_uopc,
  input  [31:0] io_dis_uops_1_bits_inst,
                io_dis_uops_1_bits_debug_inst,
  input         io_dis_uops_1_bits_is_rvc,
  input  [39:0] io_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_dis_uops_1_bits_iq_type,
  input  [9:0]  io_dis_uops_1_bits_fu_code,
  input         io_dis_uops_1_bits_is_br,
                io_dis_uops_1_bits_is_jalr,
                io_dis_uops_1_bits_is_jal,
                io_dis_uops_1_bits_is_sfb,
  input  [19:0] io_dis_uops_1_bits_br_mask,
  input  [4:0]  io_dis_uops_1_bits_br_tag,
  input  [5:0]  io_dis_uops_1_bits_ftq_idx,
  input         io_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_dis_uops_1_bits_pc_lob,
  input         io_dis_uops_1_bits_taken,
  input  [19:0] io_dis_uops_1_bits_imm_packed,
  input  [11:0] io_dis_uops_1_bits_csr_addr,
  input  [6:0]  io_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_dis_uops_1_bits_ldq_idx,
                io_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_dis_uops_1_bits_pdst,
                io_dis_uops_1_bits_prs1,
                io_dis_uops_1_bits_prs2,
                io_dis_uops_1_bits_prs3,
  input         io_dis_uops_1_bits_prs1_busy,
                io_dis_uops_1_bits_prs2_busy,
  input  [6:0]  io_dis_uops_1_bits_stale_pdst,
  input         io_dis_uops_1_bits_exception,
  input  [63:0] io_dis_uops_1_bits_exc_cause,
  input         io_dis_uops_1_bits_bypassable,
  input  [4:0]  io_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_dis_uops_1_bits_mem_size,
  input         io_dis_uops_1_bits_mem_signed,
                io_dis_uops_1_bits_is_fence,
                io_dis_uops_1_bits_is_fencei,
                io_dis_uops_1_bits_is_amo,
                io_dis_uops_1_bits_uses_ldq,
                io_dis_uops_1_bits_uses_stq,
                io_dis_uops_1_bits_is_sys_pc2epc,
                io_dis_uops_1_bits_is_unique,
                io_dis_uops_1_bits_flush_on_commit,
                io_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_1_bits_ldst,
                io_dis_uops_1_bits_lrs1,
                io_dis_uops_1_bits_lrs2,
                io_dis_uops_1_bits_lrs3,
  input         io_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_dis_uops_1_bits_dst_rtype,
                io_dis_uops_1_bits_lrs1_rtype,
                io_dis_uops_1_bits_lrs2_rtype,
  input         io_dis_uops_1_bits_frs3_en,
                io_dis_uops_1_bits_fp_val,
                io_dis_uops_1_bits_fp_single,
                io_dis_uops_1_bits_xcpt_pf_if,
                io_dis_uops_1_bits_xcpt_ae_if,
                io_dis_uops_1_bits_xcpt_ma_if,
                io_dis_uops_1_bits_bp_debug_if,
                io_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_1_bits_debug_fsrc,
                io_dis_uops_1_bits_debug_tsrc,
  output        io_dis_uops_2_ready,
  input         io_dis_uops_2_valid,
  input  [6:0]  io_dis_uops_2_bits_uopc,
  input  [31:0] io_dis_uops_2_bits_inst,
                io_dis_uops_2_bits_debug_inst,
  input         io_dis_uops_2_bits_is_rvc,
  input  [39:0] io_dis_uops_2_bits_debug_pc,
  input  [2:0]  io_dis_uops_2_bits_iq_type,
  input  [9:0]  io_dis_uops_2_bits_fu_code,
  input         io_dis_uops_2_bits_is_br,
                io_dis_uops_2_bits_is_jalr,
                io_dis_uops_2_bits_is_jal,
                io_dis_uops_2_bits_is_sfb,
  input  [19:0] io_dis_uops_2_bits_br_mask,
  input  [4:0]  io_dis_uops_2_bits_br_tag,
  input  [5:0]  io_dis_uops_2_bits_ftq_idx,
  input         io_dis_uops_2_bits_edge_inst,
  input  [5:0]  io_dis_uops_2_bits_pc_lob,
  input         io_dis_uops_2_bits_taken,
  input  [19:0] io_dis_uops_2_bits_imm_packed,
  input  [11:0] io_dis_uops_2_bits_csr_addr,
  input  [6:0]  io_dis_uops_2_bits_rob_idx,
  input  [4:0]  io_dis_uops_2_bits_ldq_idx,
                io_dis_uops_2_bits_stq_idx,
  input  [1:0]  io_dis_uops_2_bits_rxq_idx,
  input  [6:0]  io_dis_uops_2_bits_pdst,
                io_dis_uops_2_bits_prs1,
                io_dis_uops_2_bits_prs2,
                io_dis_uops_2_bits_prs3,
  input         io_dis_uops_2_bits_prs1_busy,
                io_dis_uops_2_bits_prs2_busy,
  input  [6:0]  io_dis_uops_2_bits_stale_pdst,
  input         io_dis_uops_2_bits_exception,
  input  [63:0] io_dis_uops_2_bits_exc_cause,
  input         io_dis_uops_2_bits_bypassable,
  input  [4:0]  io_dis_uops_2_bits_mem_cmd,
  input  [1:0]  io_dis_uops_2_bits_mem_size,
  input         io_dis_uops_2_bits_mem_signed,
                io_dis_uops_2_bits_is_fence,
                io_dis_uops_2_bits_is_fencei,
                io_dis_uops_2_bits_is_amo,
                io_dis_uops_2_bits_uses_ldq,
                io_dis_uops_2_bits_uses_stq,
                io_dis_uops_2_bits_is_sys_pc2epc,
                io_dis_uops_2_bits_is_unique,
                io_dis_uops_2_bits_flush_on_commit,
                io_dis_uops_2_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_2_bits_ldst,
                io_dis_uops_2_bits_lrs1,
                io_dis_uops_2_bits_lrs2,
                io_dis_uops_2_bits_lrs3,
  input         io_dis_uops_2_bits_ldst_val,
  input  [1:0]  io_dis_uops_2_bits_dst_rtype,
                io_dis_uops_2_bits_lrs1_rtype,
                io_dis_uops_2_bits_lrs2_rtype,
  input         io_dis_uops_2_bits_frs3_en,
                io_dis_uops_2_bits_fp_val,
                io_dis_uops_2_bits_fp_single,
                io_dis_uops_2_bits_xcpt_pf_if,
                io_dis_uops_2_bits_xcpt_ae_if,
                io_dis_uops_2_bits_xcpt_ma_if,
                io_dis_uops_2_bits_bp_debug_if,
                io_dis_uops_2_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_2_bits_debug_fsrc,
                io_dis_uops_2_bits_debug_tsrc,
  output        io_dis_uops_3_ready,
  input         io_dis_uops_3_valid,
  input  [6:0]  io_dis_uops_3_bits_uopc,
  input  [31:0] io_dis_uops_3_bits_inst,
                io_dis_uops_3_bits_debug_inst,
  input         io_dis_uops_3_bits_is_rvc,
  input  [39:0] io_dis_uops_3_bits_debug_pc,
  input  [2:0]  io_dis_uops_3_bits_iq_type,
  input  [9:0]  io_dis_uops_3_bits_fu_code,
  input         io_dis_uops_3_bits_is_br,
                io_dis_uops_3_bits_is_jalr,
                io_dis_uops_3_bits_is_jal,
                io_dis_uops_3_bits_is_sfb,
  input  [19:0] io_dis_uops_3_bits_br_mask,
  input  [4:0]  io_dis_uops_3_bits_br_tag,
  input  [5:0]  io_dis_uops_3_bits_ftq_idx,
  input         io_dis_uops_3_bits_edge_inst,
  input  [5:0]  io_dis_uops_3_bits_pc_lob,
  input         io_dis_uops_3_bits_taken,
  input  [19:0] io_dis_uops_3_bits_imm_packed,
  input  [11:0] io_dis_uops_3_bits_csr_addr,
  input  [6:0]  io_dis_uops_3_bits_rob_idx,
  input  [4:0]  io_dis_uops_3_bits_ldq_idx,
                io_dis_uops_3_bits_stq_idx,
  input  [1:0]  io_dis_uops_3_bits_rxq_idx,
  input  [6:0]  io_dis_uops_3_bits_pdst,
                io_dis_uops_3_bits_prs1,
                io_dis_uops_3_bits_prs2,
                io_dis_uops_3_bits_prs3,
  input         io_dis_uops_3_bits_prs1_busy,
                io_dis_uops_3_bits_prs2_busy,
  input  [6:0]  io_dis_uops_3_bits_stale_pdst,
  input         io_dis_uops_3_bits_exception,
  input  [63:0] io_dis_uops_3_bits_exc_cause,
  input         io_dis_uops_3_bits_bypassable,
  input  [4:0]  io_dis_uops_3_bits_mem_cmd,
  input  [1:0]  io_dis_uops_3_bits_mem_size,
  input         io_dis_uops_3_bits_mem_signed,
                io_dis_uops_3_bits_is_fence,
                io_dis_uops_3_bits_is_fencei,
                io_dis_uops_3_bits_is_amo,
                io_dis_uops_3_bits_uses_ldq,
                io_dis_uops_3_bits_uses_stq,
                io_dis_uops_3_bits_is_sys_pc2epc,
                io_dis_uops_3_bits_is_unique,
                io_dis_uops_3_bits_flush_on_commit,
                io_dis_uops_3_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_3_bits_ldst,
                io_dis_uops_3_bits_lrs1,
                io_dis_uops_3_bits_lrs2,
                io_dis_uops_3_bits_lrs3,
  input         io_dis_uops_3_bits_ldst_val,
  input  [1:0]  io_dis_uops_3_bits_dst_rtype,
                io_dis_uops_3_bits_lrs1_rtype,
                io_dis_uops_3_bits_lrs2_rtype,
  input         io_dis_uops_3_bits_frs3_en,
                io_dis_uops_3_bits_fp_val,
                io_dis_uops_3_bits_fp_single,
                io_dis_uops_3_bits_xcpt_pf_if,
                io_dis_uops_3_bits_xcpt_ae_if,
                io_dis_uops_3_bits_xcpt_ma_if,
                io_dis_uops_3_bits_bp_debug_if,
                io_dis_uops_3_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_3_bits_debug_fsrc,
                io_dis_uops_3_bits_debug_tsrc,
  output        io_iss_valids_0,
                io_iss_valids_1,
                io_iss_valids_2,
                io_iss_valids_3,
  output [6:0]  io_iss_uops_0_uopc,
  output [31:0] io_iss_uops_0_inst,
                io_iss_uops_0_debug_inst,
  output        io_iss_uops_0_is_rvc,
  output [39:0] io_iss_uops_0_debug_pc,
  output [2:0]  io_iss_uops_0_iq_type,
  output [9:0]  io_iss_uops_0_fu_code,
  output [1:0]  io_iss_uops_0_iw_state,
  output        io_iss_uops_0_iw_p1_poisoned,
                io_iss_uops_0_iw_p2_poisoned,
                io_iss_uops_0_is_br,
                io_iss_uops_0_is_jalr,
                io_iss_uops_0_is_jal,
                io_iss_uops_0_is_sfb,
  output [19:0] io_iss_uops_0_br_mask,
  output [4:0]  io_iss_uops_0_br_tag,
  output [5:0]  io_iss_uops_0_ftq_idx,
  output        io_iss_uops_0_edge_inst,
  output [5:0]  io_iss_uops_0_pc_lob,
  output        io_iss_uops_0_taken,
  output [19:0] io_iss_uops_0_imm_packed,
  output [11:0] io_iss_uops_0_csr_addr,
  output [6:0]  io_iss_uops_0_rob_idx,
  output [4:0]  io_iss_uops_0_ldq_idx,
                io_iss_uops_0_stq_idx,
  output [1:0]  io_iss_uops_0_rxq_idx,
  output [6:0]  io_iss_uops_0_pdst,
                io_iss_uops_0_prs1,
                io_iss_uops_0_prs2,
                io_iss_uops_0_prs3,
  output [5:0]  io_iss_uops_0_ppred,
  output        io_iss_uops_0_prs1_busy,
                io_iss_uops_0_prs2_busy,
                io_iss_uops_0_prs3_busy,
                io_iss_uops_0_ppred_busy,
  output [6:0]  io_iss_uops_0_stale_pdst,
  output        io_iss_uops_0_exception,
  output [63:0] io_iss_uops_0_exc_cause,
  output        io_iss_uops_0_bypassable,
  output [4:0]  io_iss_uops_0_mem_cmd,
  output [1:0]  io_iss_uops_0_mem_size,
  output        io_iss_uops_0_mem_signed,
                io_iss_uops_0_is_fence,
                io_iss_uops_0_is_fencei,
                io_iss_uops_0_is_amo,
                io_iss_uops_0_uses_ldq,
                io_iss_uops_0_uses_stq,
                io_iss_uops_0_is_sys_pc2epc,
                io_iss_uops_0_is_unique,
                io_iss_uops_0_flush_on_commit,
                io_iss_uops_0_ldst_is_rs1,
  output [5:0]  io_iss_uops_0_ldst,
                io_iss_uops_0_lrs1,
                io_iss_uops_0_lrs2,
                io_iss_uops_0_lrs3,
  output        io_iss_uops_0_ldst_val,
  output [1:0]  io_iss_uops_0_dst_rtype,
                io_iss_uops_0_lrs1_rtype,
                io_iss_uops_0_lrs2_rtype,
  output        io_iss_uops_0_frs3_en,
                io_iss_uops_0_fp_val,
                io_iss_uops_0_fp_single,
                io_iss_uops_0_xcpt_pf_if,
                io_iss_uops_0_xcpt_ae_if,
                io_iss_uops_0_xcpt_ma_if,
                io_iss_uops_0_bp_debug_if,
                io_iss_uops_0_bp_xcpt_if,
  output [1:0]  io_iss_uops_0_debug_fsrc,
                io_iss_uops_0_debug_tsrc,
  output [6:0]  io_iss_uops_1_uopc,
  output        io_iss_uops_1_is_rvc,
  output [9:0]  io_iss_uops_1_fu_code,
  output        io_iss_uops_1_iw_p1_poisoned,
                io_iss_uops_1_iw_p2_poisoned,
                io_iss_uops_1_is_br,
                io_iss_uops_1_is_jalr,
                io_iss_uops_1_is_jal,
                io_iss_uops_1_is_sfb,
  output [19:0] io_iss_uops_1_br_mask,
  output [4:0]  io_iss_uops_1_br_tag,
  output [5:0]  io_iss_uops_1_ftq_idx,
  output        io_iss_uops_1_edge_inst,
  output [5:0]  io_iss_uops_1_pc_lob,
  output        io_iss_uops_1_taken,
  output [19:0] io_iss_uops_1_imm_packed,
  output [6:0]  io_iss_uops_1_rob_idx,
  output [4:0]  io_iss_uops_1_ldq_idx,
                io_iss_uops_1_stq_idx,
  output [6:0]  io_iss_uops_1_pdst,
                io_iss_uops_1_prs1,
                io_iss_uops_1_prs2,
  output        io_iss_uops_1_bypassable,
  output [4:0]  io_iss_uops_1_mem_cmd,
  output        io_iss_uops_1_is_amo,
                io_iss_uops_1_uses_stq,
                io_iss_uops_1_ldst_val,
  output [1:0]  io_iss_uops_1_dst_rtype,
                io_iss_uops_1_lrs1_rtype,
                io_iss_uops_1_lrs2_rtype,
  output [6:0]  io_iss_uops_2_uopc,
  output        io_iss_uops_2_is_rvc,
  output [9:0]  io_iss_uops_2_fu_code,
  output        io_iss_uops_2_iw_p1_poisoned,
                io_iss_uops_2_iw_p2_poisoned,
                io_iss_uops_2_is_br,
                io_iss_uops_2_is_jalr,
                io_iss_uops_2_is_jal,
                io_iss_uops_2_is_sfb,
  output [19:0] io_iss_uops_2_br_mask,
  output [4:0]  io_iss_uops_2_br_tag,
  output [5:0]  io_iss_uops_2_ftq_idx,
  output        io_iss_uops_2_edge_inst,
  output [5:0]  io_iss_uops_2_pc_lob,
  output        io_iss_uops_2_taken,
  output [19:0] io_iss_uops_2_imm_packed,
  output [6:0]  io_iss_uops_2_rob_idx,
  output [4:0]  io_iss_uops_2_ldq_idx,
                io_iss_uops_2_stq_idx,
  output [6:0]  io_iss_uops_2_pdst,
                io_iss_uops_2_prs1,
                io_iss_uops_2_prs2,
  output        io_iss_uops_2_bypassable,
  output [4:0]  io_iss_uops_2_mem_cmd,
  output        io_iss_uops_2_is_amo,
                io_iss_uops_2_uses_stq,
                io_iss_uops_2_ldst_val,
  output [1:0]  io_iss_uops_2_dst_rtype,
                io_iss_uops_2_lrs1_rtype,
                io_iss_uops_2_lrs2_rtype,
  output [6:0]  io_iss_uops_3_uopc,
  output        io_iss_uops_3_is_rvc,
  output [9:0]  io_iss_uops_3_fu_code,
  output        io_iss_uops_3_iw_p1_poisoned,
                io_iss_uops_3_iw_p2_poisoned,
                io_iss_uops_3_is_br,
                io_iss_uops_3_is_jalr,
                io_iss_uops_3_is_jal,
                io_iss_uops_3_is_sfb,
  output [19:0] io_iss_uops_3_br_mask,
  output [4:0]  io_iss_uops_3_br_tag,
  output [5:0]  io_iss_uops_3_ftq_idx,
  output        io_iss_uops_3_edge_inst,
  output [5:0]  io_iss_uops_3_pc_lob,
  output        io_iss_uops_3_taken,
  output [19:0] io_iss_uops_3_imm_packed,
  output [6:0]  io_iss_uops_3_rob_idx,
  output [4:0]  io_iss_uops_3_ldq_idx,
                io_iss_uops_3_stq_idx,
  output [6:0]  io_iss_uops_3_pdst,
                io_iss_uops_3_prs1,
                io_iss_uops_3_prs2,
  output        io_iss_uops_3_bypassable,
  output [4:0]  io_iss_uops_3_mem_cmd,
  output        io_iss_uops_3_is_amo,
                io_iss_uops_3_uses_stq,
                io_iss_uops_3_ldst_val,
  output [1:0]  io_iss_uops_3_dst_rtype,
                io_iss_uops_3_lrs1_rtype,
                io_iss_uops_3_lrs2_rtype,
  input         io_wakeup_ports_0_valid,
  input  [6:0]  io_wakeup_ports_0_bits_pdst,
  input         io_wakeup_ports_1_valid,
  input  [6:0]  io_wakeup_ports_1_bits_pdst,
  input         io_wakeup_ports_2_valid,
  input  [6:0]  io_wakeup_ports_2_bits_pdst,
  input         io_wakeup_ports_3_valid,
  input  [6:0]  io_wakeup_ports_3_bits_pdst,
  input         io_wakeup_ports_4_valid,
  input  [6:0]  io_wakeup_ports_4_bits_pdst,
  input         io_wakeup_ports_5_valid,
  input  [6:0]  io_wakeup_ports_5_bits_pdst,
  input         io_wakeup_ports_6_valid,
  input  [6:0]  io_wakeup_ports_6_bits_pdst,
  input         io_wakeup_ports_7_valid,
  input  [6:0]  io_wakeup_ports_7_bits_pdst,
  input         io_wakeup_ports_8_valid,
  input  [6:0]  io_wakeup_ports_8_bits_pdst,
  input         io_wakeup_ports_9_valid,
  input  [6:0]  io_wakeup_ports_9_bits_pdst,
  input         io_spec_ld_wakeup_0_valid,
  input  [6:0]  io_spec_ld_wakeup_0_bits,
  input         io_spec_ld_wakeup_1_valid,
  input  [6:0]  io_spec_ld_wakeup_1_bits,
  input  [9:0]  io_fu_types_0,
                io_fu_types_2,
                io_fu_types_3,
  input  [19:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input         io_flush_pipeline,
                io_ld_miss
);

  wire        issue_slots_39_grant;
  wire        issue_slots_38_grant;
  wire        issue_slots_37_grant;
  wire        issue_slots_36_grant;
  wire        issue_slots_35_grant;
  wire        issue_slots_34_grant;
  wire        issue_slots_33_grant;
  wire        issue_slots_32_grant;
  wire        issue_slots_31_grant;
  wire        issue_slots_30_grant;
  wire        issue_slots_29_grant;
  wire        issue_slots_28_grant;
  wire        issue_slots_27_grant;
  wire        issue_slots_26_grant;
  wire        issue_slots_25_grant;
  wire        issue_slots_24_grant;
  wire        issue_slots_23_grant;
  wire        issue_slots_22_grant;
  wire        issue_slots_21_grant;
  wire        issue_slots_20_grant;
  wire        issue_slots_19_grant;
  wire        issue_slots_18_grant;
  wire        issue_slots_17_grant;
  wire        issue_slots_16_grant;
  wire        issue_slots_15_grant;
  wire        issue_slots_14_grant;
  wire        issue_slots_13_grant;
  wire        issue_slots_12_grant;
  wire        issue_slots_11_grant;
  wire        issue_slots_10_grant;
  wire        issue_slots_9_grant;
  wire        issue_slots_8_grant;
  wire        issue_slots_7_grant;
  wire        issue_slots_6_grant;
  wire        issue_slots_5_grant;
  wire        issue_slots_4_grant;
  wire        issue_slots_3_grant;
  wire        issue_slots_2_grant;
  wire        issue_slots_1_grant;
  wire        issue_slots_0_grant;
  wire [3:0]  next_38;
  wire [3:0]  next_37;
  wire [3:0]  next_36;
  wire [3:0]  next_35;
  wire [3:0]  next_34;
  wire [3:0]  next_33;
  wire [3:0]  next_32;
  wire [3:0]  next_31;
  wire [3:0]  next_30;
  wire [3:0]  next_29;
  wire [3:0]  next_28;
  wire [3:0]  next_27;
  wire [3:0]  next_26;
  wire [3:0]  next_25;
  wire [3:0]  next_24;
  wire [3:0]  next_23;
  wire [3:0]  next_22;
  wire [3:0]  next_21;
  wire [3:0]  next_20;
  wire [3:0]  next_19;
  wire [3:0]  next_18;
  wire [3:0]  next_17;
  wire [3:0]  next_16;
  wire [3:0]  next_15;
  wire [3:0]  next_14;
  wire [3:0]  next_13;
  wire [3:0]  next_12;
  wire [3:0]  next_11;
  wire [3:0]  next_10;
  wire [3:0]  next_9;
  wire [3:0]  next_8;
  wire [3:0]  next_7;
  wire [3:0]  next_6;
  wire [3:0]  next_5;
  wire [3:0]  next_4;
  wire [3:0]  next_3;
  wire [3:0]  next_2;
  wire [1:0]  _next_1_1to0;
  wire        _slots_39_io_valid;
  wire        _slots_39_io_will_be_valid;
  wire        _slots_39_io_request;
  wire [6:0]  _slots_39_io_out_uop_uopc;
  wire [31:0] _slots_39_io_out_uop_inst;
  wire [31:0] _slots_39_io_out_uop_debug_inst;
  wire        _slots_39_io_out_uop_is_rvc;
  wire [39:0] _slots_39_io_out_uop_debug_pc;
  wire [2:0]  _slots_39_io_out_uop_iq_type;
  wire [9:0]  _slots_39_io_out_uop_fu_code;
  wire [1:0]  _slots_39_io_out_uop_iw_state;
  wire        _slots_39_io_out_uop_iw_p1_poisoned;
  wire        _slots_39_io_out_uop_iw_p2_poisoned;
  wire        _slots_39_io_out_uop_is_br;
  wire        _slots_39_io_out_uop_is_jalr;
  wire        _slots_39_io_out_uop_is_jal;
  wire        _slots_39_io_out_uop_is_sfb;
  wire [19:0] _slots_39_io_out_uop_br_mask;
  wire [4:0]  _slots_39_io_out_uop_br_tag;
  wire [5:0]  _slots_39_io_out_uop_ftq_idx;
  wire        _slots_39_io_out_uop_edge_inst;
  wire [5:0]  _slots_39_io_out_uop_pc_lob;
  wire        _slots_39_io_out_uop_taken;
  wire [19:0] _slots_39_io_out_uop_imm_packed;
  wire [11:0] _slots_39_io_out_uop_csr_addr;
  wire [6:0]  _slots_39_io_out_uop_rob_idx;
  wire [4:0]  _slots_39_io_out_uop_ldq_idx;
  wire [4:0]  _slots_39_io_out_uop_stq_idx;
  wire [1:0]  _slots_39_io_out_uop_rxq_idx;
  wire [6:0]  _slots_39_io_out_uop_pdst;
  wire [6:0]  _slots_39_io_out_uop_prs1;
  wire [6:0]  _slots_39_io_out_uop_prs2;
  wire [6:0]  _slots_39_io_out_uop_prs3;
  wire [5:0]  _slots_39_io_out_uop_ppred;
  wire        _slots_39_io_out_uop_prs1_busy;
  wire        _slots_39_io_out_uop_prs2_busy;
  wire        _slots_39_io_out_uop_prs3_busy;
  wire        _slots_39_io_out_uop_ppred_busy;
  wire [6:0]  _slots_39_io_out_uop_stale_pdst;
  wire        _slots_39_io_out_uop_exception;
  wire [63:0] _slots_39_io_out_uop_exc_cause;
  wire        _slots_39_io_out_uop_bypassable;
  wire [4:0]  _slots_39_io_out_uop_mem_cmd;
  wire [1:0]  _slots_39_io_out_uop_mem_size;
  wire        _slots_39_io_out_uop_mem_signed;
  wire        _slots_39_io_out_uop_is_fence;
  wire        _slots_39_io_out_uop_is_fencei;
  wire        _slots_39_io_out_uop_is_amo;
  wire        _slots_39_io_out_uop_uses_ldq;
  wire        _slots_39_io_out_uop_uses_stq;
  wire        _slots_39_io_out_uop_is_sys_pc2epc;
  wire        _slots_39_io_out_uop_is_unique;
  wire        _slots_39_io_out_uop_flush_on_commit;
  wire        _slots_39_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_39_io_out_uop_ldst;
  wire [5:0]  _slots_39_io_out_uop_lrs1;
  wire [5:0]  _slots_39_io_out_uop_lrs2;
  wire [5:0]  _slots_39_io_out_uop_lrs3;
  wire        _slots_39_io_out_uop_ldst_val;
  wire [1:0]  _slots_39_io_out_uop_dst_rtype;
  wire [1:0]  _slots_39_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_39_io_out_uop_lrs2_rtype;
  wire        _slots_39_io_out_uop_frs3_en;
  wire        _slots_39_io_out_uop_fp_val;
  wire        _slots_39_io_out_uop_fp_single;
  wire        _slots_39_io_out_uop_xcpt_pf_if;
  wire        _slots_39_io_out_uop_xcpt_ae_if;
  wire        _slots_39_io_out_uop_xcpt_ma_if;
  wire        _slots_39_io_out_uop_bp_debug_if;
  wire        _slots_39_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_39_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_39_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_39_io_uop_uopc;
  wire [31:0] _slots_39_io_uop_inst;
  wire [31:0] _slots_39_io_uop_debug_inst;
  wire        _slots_39_io_uop_is_rvc;
  wire [39:0] _slots_39_io_uop_debug_pc;
  wire [2:0]  _slots_39_io_uop_iq_type;
  wire [9:0]  _slots_39_io_uop_fu_code;
  wire [1:0]  _slots_39_io_uop_iw_state;
  wire        _slots_39_io_uop_iw_p1_poisoned;
  wire        _slots_39_io_uop_iw_p2_poisoned;
  wire        _slots_39_io_uop_is_br;
  wire        _slots_39_io_uop_is_jalr;
  wire        _slots_39_io_uop_is_jal;
  wire        _slots_39_io_uop_is_sfb;
  wire [19:0] _slots_39_io_uop_br_mask;
  wire [4:0]  _slots_39_io_uop_br_tag;
  wire [5:0]  _slots_39_io_uop_ftq_idx;
  wire        _slots_39_io_uop_edge_inst;
  wire [5:0]  _slots_39_io_uop_pc_lob;
  wire        _slots_39_io_uop_taken;
  wire [19:0] _slots_39_io_uop_imm_packed;
  wire [11:0] _slots_39_io_uop_csr_addr;
  wire [6:0]  _slots_39_io_uop_rob_idx;
  wire [4:0]  _slots_39_io_uop_ldq_idx;
  wire [4:0]  _slots_39_io_uop_stq_idx;
  wire [1:0]  _slots_39_io_uop_rxq_idx;
  wire [6:0]  _slots_39_io_uop_pdst;
  wire [6:0]  _slots_39_io_uop_prs1;
  wire [6:0]  _slots_39_io_uop_prs2;
  wire [6:0]  _slots_39_io_uop_prs3;
  wire [5:0]  _slots_39_io_uop_ppred;
  wire        _slots_39_io_uop_prs1_busy;
  wire        _slots_39_io_uop_prs2_busy;
  wire        _slots_39_io_uop_prs3_busy;
  wire        _slots_39_io_uop_ppred_busy;
  wire [6:0]  _slots_39_io_uop_stale_pdst;
  wire        _slots_39_io_uop_exception;
  wire [63:0] _slots_39_io_uop_exc_cause;
  wire        _slots_39_io_uop_bypassable;
  wire [4:0]  _slots_39_io_uop_mem_cmd;
  wire [1:0]  _slots_39_io_uop_mem_size;
  wire        _slots_39_io_uop_mem_signed;
  wire        _slots_39_io_uop_is_fence;
  wire        _slots_39_io_uop_is_fencei;
  wire        _slots_39_io_uop_is_amo;
  wire        _slots_39_io_uop_uses_ldq;
  wire        _slots_39_io_uop_uses_stq;
  wire        _slots_39_io_uop_is_sys_pc2epc;
  wire        _slots_39_io_uop_is_unique;
  wire        _slots_39_io_uop_flush_on_commit;
  wire        _slots_39_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_39_io_uop_ldst;
  wire [5:0]  _slots_39_io_uop_lrs1;
  wire [5:0]  _slots_39_io_uop_lrs2;
  wire [5:0]  _slots_39_io_uop_lrs3;
  wire        _slots_39_io_uop_ldst_val;
  wire [1:0]  _slots_39_io_uop_dst_rtype;
  wire [1:0]  _slots_39_io_uop_lrs1_rtype;
  wire [1:0]  _slots_39_io_uop_lrs2_rtype;
  wire        _slots_39_io_uop_frs3_en;
  wire        _slots_39_io_uop_fp_val;
  wire        _slots_39_io_uop_fp_single;
  wire        _slots_39_io_uop_xcpt_pf_if;
  wire        _slots_39_io_uop_xcpt_ae_if;
  wire        _slots_39_io_uop_xcpt_ma_if;
  wire        _slots_39_io_uop_bp_debug_if;
  wire        _slots_39_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_39_io_uop_debug_fsrc;
  wire [1:0]  _slots_39_io_uop_debug_tsrc;
  wire        _slots_38_io_valid;
  wire        _slots_38_io_will_be_valid;
  wire        _slots_38_io_request;
  wire [6:0]  _slots_38_io_out_uop_uopc;
  wire [31:0] _slots_38_io_out_uop_inst;
  wire [31:0] _slots_38_io_out_uop_debug_inst;
  wire        _slots_38_io_out_uop_is_rvc;
  wire [39:0] _slots_38_io_out_uop_debug_pc;
  wire [2:0]  _slots_38_io_out_uop_iq_type;
  wire [9:0]  _slots_38_io_out_uop_fu_code;
  wire [1:0]  _slots_38_io_out_uop_iw_state;
  wire        _slots_38_io_out_uop_iw_p1_poisoned;
  wire        _slots_38_io_out_uop_iw_p2_poisoned;
  wire        _slots_38_io_out_uop_is_br;
  wire        _slots_38_io_out_uop_is_jalr;
  wire        _slots_38_io_out_uop_is_jal;
  wire        _slots_38_io_out_uop_is_sfb;
  wire [19:0] _slots_38_io_out_uop_br_mask;
  wire [4:0]  _slots_38_io_out_uop_br_tag;
  wire [5:0]  _slots_38_io_out_uop_ftq_idx;
  wire        _slots_38_io_out_uop_edge_inst;
  wire [5:0]  _slots_38_io_out_uop_pc_lob;
  wire        _slots_38_io_out_uop_taken;
  wire [19:0] _slots_38_io_out_uop_imm_packed;
  wire [11:0] _slots_38_io_out_uop_csr_addr;
  wire [6:0]  _slots_38_io_out_uop_rob_idx;
  wire [4:0]  _slots_38_io_out_uop_ldq_idx;
  wire [4:0]  _slots_38_io_out_uop_stq_idx;
  wire [1:0]  _slots_38_io_out_uop_rxq_idx;
  wire [6:0]  _slots_38_io_out_uop_pdst;
  wire [6:0]  _slots_38_io_out_uop_prs1;
  wire [6:0]  _slots_38_io_out_uop_prs2;
  wire [6:0]  _slots_38_io_out_uop_prs3;
  wire [5:0]  _slots_38_io_out_uop_ppred;
  wire        _slots_38_io_out_uop_prs1_busy;
  wire        _slots_38_io_out_uop_prs2_busy;
  wire        _slots_38_io_out_uop_prs3_busy;
  wire        _slots_38_io_out_uop_ppred_busy;
  wire [6:0]  _slots_38_io_out_uop_stale_pdst;
  wire        _slots_38_io_out_uop_exception;
  wire [63:0] _slots_38_io_out_uop_exc_cause;
  wire        _slots_38_io_out_uop_bypassable;
  wire [4:0]  _slots_38_io_out_uop_mem_cmd;
  wire [1:0]  _slots_38_io_out_uop_mem_size;
  wire        _slots_38_io_out_uop_mem_signed;
  wire        _slots_38_io_out_uop_is_fence;
  wire        _slots_38_io_out_uop_is_fencei;
  wire        _slots_38_io_out_uop_is_amo;
  wire        _slots_38_io_out_uop_uses_ldq;
  wire        _slots_38_io_out_uop_uses_stq;
  wire        _slots_38_io_out_uop_is_sys_pc2epc;
  wire        _slots_38_io_out_uop_is_unique;
  wire        _slots_38_io_out_uop_flush_on_commit;
  wire        _slots_38_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_38_io_out_uop_ldst;
  wire [5:0]  _slots_38_io_out_uop_lrs1;
  wire [5:0]  _slots_38_io_out_uop_lrs2;
  wire [5:0]  _slots_38_io_out_uop_lrs3;
  wire        _slots_38_io_out_uop_ldst_val;
  wire [1:0]  _slots_38_io_out_uop_dst_rtype;
  wire [1:0]  _slots_38_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_38_io_out_uop_lrs2_rtype;
  wire        _slots_38_io_out_uop_frs3_en;
  wire        _slots_38_io_out_uop_fp_val;
  wire        _slots_38_io_out_uop_fp_single;
  wire        _slots_38_io_out_uop_xcpt_pf_if;
  wire        _slots_38_io_out_uop_xcpt_ae_if;
  wire        _slots_38_io_out_uop_xcpt_ma_if;
  wire        _slots_38_io_out_uop_bp_debug_if;
  wire        _slots_38_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_38_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_38_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_38_io_uop_uopc;
  wire [31:0] _slots_38_io_uop_inst;
  wire [31:0] _slots_38_io_uop_debug_inst;
  wire        _slots_38_io_uop_is_rvc;
  wire [39:0] _slots_38_io_uop_debug_pc;
  wire [2:0]  _slots_38_io_uop_iq_type;
  wire [9:0]  _slots_38_io_uop_fu_code;
  wire [1:0]  _slots_38_io_uop_iw_state;
  wire        _slots_38_io_uop_iw_p1_poisoned;
  wire        _slots_38_io_uop_iw_p2_poisoned;
  wire        _slots_38_io_uop_is_br;
  wire        _slots_38_io_uop_is_jalr;
  wire        _slots_38_io_uop_is_jal;
  wire        _slots_38_io_uop_is_sfb;
  wire [19:0] _slots_38_io_uop_br_mask;
  wire [4:0]  _slots_38_io_uop_br_tag;
  wire [5:0]  _slots_38_io_uop_ftq_idx;
  wire        _slots_38_io_uop_edge_inst;
  wire [5:0]  _slots_38_io_uop_pc_lob;
  wire        _slots_38_io_uop_taken;
  wire [19:0] _slots_38_io_uop_imm_packed;
  wire [11:0] _slots_38_io_uop_csr_addr;
  wire [6:0]  _slots_38_io_uop_rob_idx;
  wire [4:0]  _slots_38_io_uop_ldq_idx;
  wire [4:0]  _slots_38_io_uop_stq_idx;
  wire [1:0]  _slots_38_io_uop_rxq_idx;
  wire [6:0]  _slots_38_io_uop_pdst;
  wire [6:0]  _slots_38_io_uop_prs1;
  wire [6:0]  _slots_38_io_uop_prs2;
  wire [6:0]  _slots_38_io_uop_prs3;
  wire [5:0]  _slots_38_io_uop_ppred;
  wire        _slots_38_io_uop_prs1_busy;
  wire        _slots_38_io_uop_prs2_busy;
  wire        _slots_38_io_uop_prs3_busy;
  wire        _slots_38_io_uop_ppred_busy;
  wire [6:0]  _slots_38_io_uop_stale_pdst;
  wire        _slots_38_io_uop_exception;
  wire [63:0] _slots_38_io_uop_exc_cause;
  wire        _slots_38_io_uop_bypassable;
  wire [4:0]  _slots_38_io_uop_mem_cmd;
  wire [1:0]  _slots_38_io_uop_mem_size;
  wire        _slots_38_io_uop_mem_signed;
  wire        _slots_38_io_uop_is_fence;
  wire        _slots_38_io_uop_is_fencei;
  wire        _slots_38_io_uop_is_amo;
  wire        _slots_38_io_uop_uses_ldq;
  wire        _slots_38_io_uop_uses_stq;
  wire        _slots_38_io_uop_is_sys_pc2epc;
  wire        _slots_38_io_uop_is_unique;
  wire        _slots_38_io_uop_flush_on_commit;
  wire        _slots_38_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_38_io_uop_ldst;
  wire [5:0]  _slots_38_io_uop_lrs1;
  wire [5:0]  _slots_38_io_uop_lrs2;
  wire [5:0]  _slots_38_io_uop_lrs3;
  wire        _slots_38_io_uop_ldst_val;
  wire [1:0]  _slots_38_io_uop_dst_rtype;
  wire [1:0]  _slots_38_io_uop_lrs1_rtype;
  wire [1:0]  _slots_38_io_uop_lrs2_rtype;
  wire        _slots_38_io_uop_frs3_en;
  wire        _slots_38_io_uop_fp_val;
  wire        _slots_38_io_uop_fp_single;
  wire        _slots_38_io_uop_xcpt_pf_if;
  wire        _slots_38_io_uop_xcpt_ae_if;
  wire        _slots_38_io_uop_xcpt_ma_if;
  wire        _slots_38_io_uop_bp_debug_if;
  wire        _slots_38_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_38_io_uop_debug_fsrc;
  wire [1:0]  _slots_38_io_uop_debug_tsrc;
  wire        _slots_37_io_valid;
  wire        _slots_37_io_will_be_valid;
  wire        _slots_37_io_request;
  wire [6:0]  _slots_37_io_out_uop_uopc;
  wire [31:0] _slots_37_io_out_uop_inst;
  wire [31:0] _slots_37_io_out_uop_debug_inst;
  wire        _slots_37_io_out_uop_is_rvc;
  wire [39:0] _slots_37_io_out_uop_debug_pc;
  wire [2:0]  _slots_37_io_out_uop_iq_type;
  wire [9:0]  _slots_37_io_out_uop_fu_code;
  wire [1:0]  _slots_37_io_out_uop_iw_state;
  wire        _slots_37_io_out_uop_iw_p1_poisoned;
  wire        _slots_37_io_out_uop_iw_p2_poisoned;
  wire        _slots_37_io_out_uop_is_br;
  wire        _slots_37_io_out_uop_is_jalr;
  wire        _slots_37_io_out_uop_is_jal;
  wire        _slots_37_io_out_uop_is_sfb;
  wire [19:0] _slots_37_io_out_uop_br_mask;
  wire [4:0]  _slots_37_io_out_uop_br_tag;
  wire [5:0]  _slots_37_io_out_uop_ftq_idx;
  wire        _slots_37_io_out_uop_edge_inst;
  wire [5:0]  _slots_37_io_out_uop_pc_lob;
  wire        _slots_37_io_out_uop_taken;
  wire [19:0] _slots_37_io_out_uop_imm_packed;
  wire [11:0] _slots_37_io_out_uop_csr_addr;
  wire [6:0]  _slots_37_io_out_uop_rob_idx;
  wire [4:0]  _slots_37_io_out_uop_ldq_idx;
  wire [4:0]  _slots_37_io_out_uop_stq_idx;
  wire [1:0]  _slots_37_io_out_uop_rxq_idx;
  wire [6:0]  _slots_37_io_out_uop_pdst;
  wire [6:0]  _slots_37_io_out_uop_prs1;
  wire [6:0]  _slots_37_io_out_uop_prs2;
  wire [6:0]  _slots_37_io_out_uop_prs3;
  wire [5:0]  _slots_37_io_out_uop_ppred;
  wire        _slots_37_io_out_uop_prs1_busy;
  wire        _slots_37_io_out_uop_prs2_busy;
  wire        _slots_37_io_out_uop_prs3_busy;
  wire        _slots_37_io_out_uop_ppred_busy;
  wire [6:0]  _slots_37_io_out_uop_stale_pdst;
  wire        _slots_37_io_out_uop_exception;
  wire [63:0] _slots_37_io_out_uop_exc_cause;
  wire        _slots_37_io_out_uop_bypassable;
  wire [4:0]  _slots_37_io_out_uop_mem_cmd;
  wire [1:0]  _slots_37_io_out_uop_mem_size;
  wire        _slots_37_io_out_uop_mem_signed;
  wire        _slots_37_io_out_uop_is_fence;
  wire        _slots_37_io_out_uop_is_fencei;
  wire        _slots_37_io_out_uop_is_amo;
  wire        _slots_37_io_out_uop_uses_ldq;
  wire        _slots_37_io_out_uop_uses_stq;
  wire        _slots_37_io_out_uop_is_sys_pc2epc;
  wire        _slots_37_io_out_uop_is_unique;
  wire        _slots_37_io_out_uop_flush_on_commit;
  wire        _slots_37_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_37_io_out_uop_ldst;
  wire [5:0]  _slots_37_io_out_uop_lrs1;
  wire [5:0]  _slots_37_io_out_uop_lrs2;
  wire [5:0]  _slots_37_io_out_uop_lrs3;
  wire        _slots_37_io_out_uop_ldst_val;
  wire [1:0]  _slots_37_io_out_uop_dst_rtype;
  wire [1:0]  _slots_37_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_37_io_out_uop_lrs2_rtype;
  wire        _slots_37_io_out_uop_frs3_en;
  wire        _slots_37_io_out_uop_fp_val;
  wire        _slots_37_io_out_uop_fp_single;
  wire        _slots_37_io_out_uop_xcpt_pf_if;
  wire        _slots_37_io_out_uop_xcpt_ae_if;
  wire        _slots_37_io_out_uop_xcpt_ma_if;
  wire        _slots_37_io_out_uop_bp_debug_if;
  wire        _slots_37_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_37_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_37_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_37_io_uop_uopc;
  wire [31:0] _slots_37_io_uop_inst;
  wire [31:0] _slots_37_io_uop_debug_inst;
  wire        _slots_37_io_uop_is_rvc;
  wire [39:0] _slots_37_io_uop_debug_pc;
  wire [2:0]  _slots_37_io_uop_iq_type;
  wire [9:0]  _slots_37_io_uop_fu_code;
  wire [1:0]  _slots_37_io_uop_iw_state;
  wire        _slots_37_io_uop_iw_p1_poisoned;
  wire        _slots_37_io_uop_iw_p2_poisoned;
  wire        _slots_37_io_uop_is_br;
  wire        _slots_37_io_uop_is_jalr;
  wire        _slots_37_io_uop_is_jal;
  wire        _slots_37_io_uop_is_sfb;
  wire [19:0] _slots_37_io_uop_br_mask;
  wire [4:0]  _slots_37_io_uop_br_tag;
  wire [5:0]  _slots_37_io_uop_ftq_idx;
  wire        _slots_37_io_uop_edge_inst;
  wire [5:0]  _slots_37_io_uop_pc_lob;
  wire        _slots_37_io_uop_taken;
  wire [19:0] _slots_37_io_uop_imm_packed;
  wire [11:0] _slots_37_io_uop_csr_addr;
  wire [6:0]  _slots_37_io_uop_rob_idx;
  wire [4:0]  _slots_37_io_uop_ldq_idx;
  wire [4:0]  _slots_37_io_uop_stq_idx;
  wire [1:0]  _slots_37_io_uop_rxq_idx;
  wire [6:0]  _slots_37_io_uop_pdst;
  wire [6:0]  _slots_37_io_uop_prs1;
  wire [6:0]  _slots_37_io_uop_prs2;
  wire [6:0]  _slots_37_io_uop_prs3;
  wire [5:0]  _slots_37_io_uop_ppred;
  wire        _slots_37_io_uop_prs1_busy;
  wire        _slots_37_io_uop_prs2_busy;
  wire        _slots_37_io_uop_prs3_busy;
  wire        _slots_37_io_uop_ppred_busy;
  wire [6:0]  _slots_37_io_uop_stale_pdst;
  wire        _slots_37_io_uop_exception;
  wire [63:0] _slots_37_io_uop_exc_cause;
  wire        _slots_37_io_uop_bypassable;
  wire [4:0]  _slots_37_io_uop_mem_cmd;
  wire [1:0]  _slots_37_io_uop_mem_size;
  wire        _slots_37_io_uop_mem_signed;
  wire        _slots_37_io_uop_is_fence;
  wire        _slots_37_io_uop_is_fencei;
  wire        _slots_37_io_uop_is_amo;
  wire        _slots_37_io_uop_uses_ldq;
  wire        _slots_37_io_uop_uses_stq;
  wire        _slots_37_io_uop_is_sys_pc2epc;
  wire        _slots_37_io_uop_is_unique;
  wire        _slots_37_io_uop_flush_on_commit;
  wire        _slots_37_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_37_io_uop_ldst;
  wire [5:0]  _slots_37_io_uop_lrs1;
  wire [5:0]  _slots_37_io_uop_lrs2;
  wire [5:0]  _slots_37_io_uop_lrs3;
  wire        _slots_37_io_uop_ldst_val;
  wire [1:0]  _slots_37_io_uop_dst_rtype;
  wire [1:0]  _slots_37_io_uop_lrs1_rtype;
  wire [1:0]  _slots_37_io_uop_lrs2_rtype;
  wire        _slots_37_io_uop_frs3_en;
  wire        _slots_37_io_uop_fp_val;
  wire        _slots_37_io_uop_fp_single;
  wire        _slots_37_io_uop_xcpt_pf_if;
  wire        _slots_37_io_uop_xcpt_ae_if;
  wire        _slots_37_io_uop_xcpt_ma_if;
  wire        _slots_37_io_uop_bp_debug_if;
  wire        _slots_37_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_37_io_uop_debug_fsrc;
  wire [1:0]  _slots_37_io_uop_debug_tsrc;
  wire        _slots_36_io_valid;
  wire        _slots_36_io_will_be_valid;
  wire        _slots_36_io_request;
  wire [6:0]  _slots_36_io_out_uop_uopc;
  wire [31:0] _slots_36_io_out_uop_inst;
  wire [31:0] _slots_36_io_out_uop_debug_inst;
  wire        _slots_36_io_out_uop_is_rvc;
  wire [39:0] _slots_36_io_out_uop_debug_pc;
  wire [2:0]  _slots_36_io_out_uop_iq_type;
  wire [9:0]  _slots_36_io_out_uop_fu_code;
  wire [1:0]  _slots_36_io_out_uop_iw_state;
  wire        _slots_36_io_out_uop_iw_p1_poisoned;
  wire        _slots_36_io_out_uop_iw_p2_poisoned;
  wire        _slots_36_io_out_uop_is_br;
  wire        _slots_36_io_out_uop_is_jalr;
  wire        _slots_36_io_out_uop_is_jal;
  wire        _slots_36_io_out_uop_is_sfb;
  wire [19:0] _slots_36_io_out_uop_br_mask;
  wire [4:0]  _slots_36_io_out_uop_br_tag;
  wire [5:0]  _slots_36_io_out_uop_ftq_idx;
  wire        _slots_36_io_out_uop_edge_inst;
  wire [5:0]  _slots_36_io_out_uop_pc_lob;
  wire        _slots_36_io_out_uop_taken;
  wire [19:0] _slots_36_io_out_uop_imm_packed;
  wire [11:0] _slots_36_io_out_uop_csr_addr;
  wire [6:0]  _slots_36_io_out_uop_rob_idx;
  wire [4:0]  _slots_36_io_out_uop_ldq_idx;
  wire [4:0]  _slots_36_io_out_uop_stq_idx;
  wire [1:0]  _slots_36_io_out_uop_rxq_idx;
  wire [6:0]  _slots_36_io_out_uop_pdst;
  wire [6:0]  _slots_36_io_out_uop_prs1;
  wire [6:0]  _slots_36_io_out_uop_prs2;
  wire [6:0]  _slots_36_io_out_uop_prs3;
  wire [5:0]  _slots_36_io_out_uop_ppred;
  wire        _slots_36_io_out_uop_prs1_busy;
  wire        _slots_36_io_out_uop_prs2_busy;
  wire        _slots_36_io_out_uop_prs3_busy;
  wire        _slots_36_io_out_uop_ppred_busy;
  wire [6:0]  _slots_36_io_out_uop_stale_pdst;
  wire        _slots_36_io_out_uop_exception;
  wire [63:0] _slots_36_io_out_uop_exc_cause;
  wire        _slots_36_io_out_uop_bypassable;
  wire [4:0]  _slots_36_io_out_uop_mem_cmd;
  wire [1:0]  _slots_36_io_out_uop_mem_size;
  wire        _slots_36_io_out_uop_mem_signed;
  wire        _slots_36_io_out_uop_is_fence;
  wire        _slots_36_io_out_uop_is_fencei;
  wire        _slots_36_io_out_uop_is_amo;
  wire        _slots_36_io_out_uop_uses_ldq;
  wire        _slots_36_io_out_uop_uses_stq;
  wire        _slots_36_io_out_uop_is_sys_pc2epc;
  wire        _slots_36_io_out_uop_is_unique;
  wire        _slots_36_io_out_uop_flush_on_commit;
  wire        _slots_36_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_36_io_out_uop_ldst;
  wire [5:0]  _slots_36_io_out_uop_lrs1;
  wire [5:0]  _slots_36_io_out_uop_lrs2;
  wire [5:0]  _slots_36_io_out_uop_lrs3;
  wire        _slots_36_io_out_uop_ldst_val;
  wire [1:0]  _slots_36_io_out_uop_dst_rtype;
  wire [1:0]  _slots_36_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_36_io_out_uop_lrs2_rtype;
  wire        _slots_36_io_out_uop_frs3_en;
  wire        _slots_36_io_out_uop_fp_val;
  wire        _slots_36_io_out_uop_fp_single;
  wire        _slots_36_io_out_uop_xcpt_pf_if;
  wire        _slots_36_io_out_uop_xcpt_ae_if;
  wire        _slots_36_io_out_uop_xcpt_ma_if;
  wire        _slots_36_io_out_uop_bp_debug_if;
  wire        _slots_36_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_36_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_36_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_36_io_uop_uopc;
  wire [31:0] _slots_36_io_uop_inst;
  wire [31:0] _slots_36_io_uop_debug_inst;
  wire        _slots_36_io_uop_is_rvc;
  wire [39:0] _slots_36_io_uop_debug_pc;
  wire [2:0]  _slots_36_io_uop_iq_type;
  wire [9:0]  _slots_36_io_uop_fu_code;
  wire [1:0]  _slots_36_io_uop_iw_state;
  wire        _slots_36_io_uop_iw_p1_poisoned;
  wire        _slots_36_io_uop_iw_p2_poisoned;
  wire        _slots_36_io_uop_is_br;
  wire        _slots_36_io_uop_is_jalr;
  wire        _slots_36_io_uop_is_jal;
  wire        _slots_36_io_uop_is_sfb;
  wire [19:0] _slots_36_io_uop_br_mask;
  wire [4:0]  _slots_36_io_uop_br_tag;
  wire [5:0]  _slots_36_io_uop_ftq_idx;
  wire        _slots_36_io_uop_edge_inst;
  wire [5:0]  _slots_36_io_uop_pc_lob;
  wire        _slots_36_io_uop_taken;
  wire [19:0] _slots_36_io_uop_imm_packed;
  wire [11:0] _slots_36_io_uop_csr_addr;
  wire [6:0]  _slots_36_io_uop_rob_idx;
  wire [4:0]  _slots_36_io_uop_ldq_idx;
  wire [4:0]  _slots_36_io_uop_stq_idx;
  wire [1:0]  _slots_36_io_uop_rxq_idx;
  wire [6:0]  _slots_36_io_uop_pdst;
  wire [6:0]  _slots_36_io_uop_prs1;
  wire [6:0]  _slots_36_io_uop_prs2;
  wire [6:0]  _slots_36_io_uop_prs3;
  wire [5:0]  _slots_36_io_uop_ppred;
  wire        _slots_36_io_uop_prs1_busy;
  wire        _slots_36_io_uop_prs2_busy;
  wire        _slots_36_io_uop_prs3_busy;
  wire        _slots_36_io_uop_ppred_busy;
  wire [6:0]  _slots_36_io_uop_stale_pdst;
  wire        _slots_36_io_uop_exception;
  wire [63:0] _slots_36_io_uop_exc_cause;
  wire        _slots_36_io_uop_bypassable;
  wire [4:0]  _slots_36_io_uop_mem_cmd;
  wire [1:0]  _slots_36_io_uop_mem_size;
  wire        _slots_36_io_uop_mem_signed;
  wire        _slots_36_io_uop_is_fence;
  wire        _slots_36_io_uop_is_fencei;
  wire        _slots_36_io_uop_is_amo;
  wire        _slots_36_io_uop_uses_ldq;
  wire        _slots_36_io_uop_uses_stq;
  wire        _slots_36_io_uop_is_sys_pc2epc;
  wire        _slots_36_io_uop_is_unique;
  wire        _slots_36_io_uop_flush_on_commit;
  wire        _slots_36_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_36_io_uop_ldst;
  wire [5:0]  _slots_36_io_uop_lrs1;
  wire [5:0]  _slots_36_io_uop_lrs2;
  wire [5:0]  _slots_36_io_uop_lrs3;
  wire        _slots_36_io_uop_ldst_val;
  wire [1:0]  _slots_36_io_uop_dst_rtype;
  wire [1:0]  _slots_36_io_uop_lrs1_rtype;
  wire [1:0]  _slots_36_io_uop_lrs2_rtype;
  wire        _slots_36_io_uop_frs3_en;
  wire        _slots_36_io_uop_fp_val;
  wire        _slots_36_io_uop_fp_single;
  wire        _slots_36_io_uop_xcpt_pf_if;
  wire        _slots_36_io_uop_xcpt_ae_if;
  wire        _slots_36_io_uop_xcpt_ma_if;
  wire        _slots_36_io_uop_bp_debug_if;
  wire        _slots_36_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_36_io_uop_debug_fsrc;
  wire [1:0]  _slots_36_io_uop_debug_tsrc;
  wire        _slots_35_io_valid;
  wire        _slots_35_io_will_be_valid;
  wire        _slots_35_io_request;
  wire [6:0]  _slots_35_io_out_uop_uopc;
  wire [31:0] _slots_35_io_out_uop_inst;
  wire [31:0] _slots_35_io_out_uop_debug_inst;
  wire        _slots_35_io_out_uop_is_rvc;
  wire [39:0] _slots_35_io_out_uop_debug_pc;
  wire [2:0]  _slots_35_io_out_uop_iq_type;
  wire [9:0]  _slots_35_io_out_uop_fu_code;
  wire [1:0]  _slots_35_io_out_uop_iw_state;
  wire        _slots_35_io_out_uop_iw_p1_poisoned;
  wire        _slots_35_io_out_uop_iw_p2_poisoned;
  wire        _slots_35_io_out_uop_is_br;
  wire        _slots_35_io_out_uop_is_jalr;
  wire        _slots_35_io_out_uop_is_jal;
  wire        _slots_35_io_out_uop_is_sfb;
  wire [19:0] _slots_35_io_out_uop_br_mask;
  wire [4:0]  _slots_35_io_out_uop_br_tag;
  wire [5:0]  _slots_35_io_out_uop_ftq_idx;
  wire        _slots_35_io_out_uop_edge_inst;
  wire [5:0]  _slots_35_io_out_uop_pc_lob;
  wire        _slots_35_io_out_uop_taken;
  wire [19:0] _slots_35_io_out_uop_imm_packed;
  wire [11:0] _slots_35_io_out_uop_csr_addr;
  wire [6:0]  _slots_35_io_out_uop_rob_idx;
  wire [4:0]  _slots_35_io_out_uop_ldq_idx;
  wire [4:0]  _slots_35_io_out_uop_stq_idx;
  wire [1:0]  _slots_35_io_out_uop_rxq_idx;
  wire [6:0]  _slots_35_io_out_uop_pdst;
  wire [6:0]  _slots_35_io_out_uop_prs1;
  wire [6:0]  _slots_35_io_out_uop_prs2;
  wire [6:0]  _slots_35_io_out_uop_prs3;
  wire [5:0]  _slots_35_io_out_uop_ppred;
  wire        _slots_35_io_out_uop_prs1_busy;
  wire        _slots_35_io_out_uop_prs2_busy;
  wire        _slots_35_io_out_uop_prs3_busy;
  wire        _slots_35_io_out_uop_ppred_busy;
  wire [6:0]  _slots_35_io_out_uop_stale_pdst;
  wire        _slots_35_io_out_uop_exception;
  wire [63:0] _slots_35_io_out_uop_exc_cause;
  wire        _slots_35_io_out_uop_bypassable;
  wire [4:0]  _slots_35_io_out_uop_mem_cmd;
  wire [1:0]  _slots_35_io_out_uop_mem_size;
  wire        _slots_35_io_out_uop_mem_signed;
  wire        _slots_35_io_out_uop_is_fence;
  wire        _slots_35_io_out_uop_is_fencei;
  wire        _slots_35_io_out_uop_is_amo;
  wire        _slots_35_io_out_uop_uses_ldq;
  wire        _slots_35_io_out_uop_uses_stq;
  wire        _slots_35_io_out_uop_is_sys_pc2epc;
  wire        _slots_35_io_out_uop_is_unique;
  wire        _slots_35_io_out_uop_flush_on_commit;
  wire        _slots_35_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_35_io_out_uop_ldst;
  wire [5:0]  _slots_35_io_out_uop_lrs1;
  wire [5:0]  _slots_35_io_out_uop_lrs2;
  wire [5:0]  _slots_35_io_out_uop_lrs3;
  wire        _slots_35_io_out_uop_ldst_val;
  wire [1:0]  _slots_35_io_out_uop_dst_rtype;
  wire [1:0]  _slots_35_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_35_io_out_uop_lrs2_rtype;
  wire        _slots_35_io_out_uop_frs3_en;
  wire        _slots_35_io_out_uop_fp_val;
  wire        _slots_35_io_out_uop_fp_single;
  wire        _slots_35_io_out_uop_xcpt_pf_if;
  wire        _slots_35_io_out_uop_xcpt_ae_if;
  wire        _slots_35_io_out_uop_xcpt_ma_if;
  wire        _slots_35_io_out_uop_bp_debug_if;
  wire        _slots_35_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_35_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_35_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_35_io_uop_uopc;
  wire [31:0] _slots_35_io_uop_inst;
  wire [31:0] _slots_35_io_uop_debug_inst;
  wire        _slots_35_io_uop_is_rvc;
  wire [39:0] _slots_35_io_uop_debug_pc;
  wire [2:0]  _slots_35_io_uop_iq_type;
  wire [9:0]  _slots_35_io_uop_fu_code;
  wire [1:0]  _slots_35_io_uop_iw_state;
  wire        _slots_35_io_uop_iw_p1_poisoned;
  wire        _slots_35_io_uop_iw_p2_poisoned;
  wire        _slots_35_io_uop_is_br;
  wire        _slots_35_io_uop_is_jalr;
  wire        _slots_35_io_uop_is_jal;
  wire        _slots_35_io_uop_is_sfb;
  wire [19:0] _slots_35_io_uop_br_mask;
  wire [4:0]  _slots_35_io_uop_br_tag;
  wire [5:0]  _slots_35_io_uop_ftq_idx;
  wire        _slots_35_io_uop_edge_inst;
  wire [5:0]  _slots_35_io_uop_pc_lob;
  wire        _slots_35_io_uop_taken;
  wire [19:0] _slots_35_io_uop_imm_packed;
  wire [11:0] _slots_35_io_uop_csr_addr;
  wire [6:0]  _slots_35_io_uop_rob_idx;
  wire [4:0]  _slots_35_io_uop_ldq_idx;
  wire [4:0]  _slots_35_io_uop_stq_idx;
  wire [1:0]  _slots_35_io_uop_rxq_idx;
  wire [6:0]  _slots_35_io_uop_pdst;
  wire [6:0]  _slots_35_io_uop_prs1;
  wire [6:0]  _slots_35_io_uop_prs2;
  wire [6:0]  _slots_35_io_uop_prs3;
  wire [5:0]  _slots_35_io_uop_ppred;
  wire        _slots_35_io_uop_prs1_busy;
  wire        _slots_35_io_uop_prs2_busy;
  wire        _slots_35_io_uop_prs3_busy;
  wire        _slots_35_io_uop_ppred_busy;
  wire [6:0]  _slots_35_io_uop_stale_pdst;
  wire        _slots_35_io_uop_exception;
  wire [63:0] _slots_35_io_uop_exc_cause;
  wire        _slots_35_io_uop_bypassable;
  wire [4:0]  _slots_35_io_uop_mem_cmd;
  wire [1:0]  _slots_35_io_uop_mem_size;
  wire        _slots_35_io_uop_mem_signed;
  wire        _slots_35_io_uop_is_fence;
  wire        _slots_35_io_uop_is_fencei;
  wire        _slots_35_io_uop_is_amo;
  wire        _slots_35_io_uop_uses_ldq;
  wire        _slots_35_io_uop_uses_stq;
  wire        _slots_35_io_uop_is_sys_pc2epc;
  wire        _slots_35_io_uop_is_unique;
  wire        _slots_35_io_uop_flush_on_commit;
  wire        _slots_35_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_35_io_uop_ldst;
  wire [5:0]  _slots_35_io_uop_lrs1;
  wire [5:0]  _slots_35_io_uop_lrs2;
  wire [5:0]  _slots_35_io_uop_lrs3;
  wire        _slots_35_io_uop_ldst_val;
  wire [1:0]  _slots_35_io_uop_dst_rtype;
  wire [1:0]  _slots_35_io_uop_lrs1_rtype;
  wire [1:0]  _slots_35_io_uop_lrs2_rtype;
  wire        _slots_35_io_uop_frs3_en;
  wire        _slots_35_io_uop_fp_val;
  wire        _slots_35_io_uop_fp_single;
  wire        _slots_35_io_uop_xcpt_pf_if;
  wire        _slots_35_io_uop_xcpt_ae_if;
  wire        _slots_35_io_uop_xcpt_ma_if;
  wire        _slots_35_io_uop_bp_debug_if;
  wire        _slots_35_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_35_io_uop_debug_fsrc;
  wire [1:0]  _slots_35_io_uop_debug_tsrc;
  wire        _slots_34_io_valid;
  wire        _slots_34_io_will_be_valid;
  wire        _slots_34_io_request;
  wire [6:0]  _slots_34_io_out_uop_uopc;
  wire [31:0] _slots_34_io_out_uop_inst;
  wire [31:0] _slots_34_io_out_uop_debug_inst;
  wire        _slots_34_io_out_uop_is_rvc;
  wire [39:0] _slots_34_io_out_uop_debug_pc;
  wire [2:0]  _slots_34_io_out_uop_iq_type;
  wire [9:0]  _slots_34_io_out_uop_fu_code;
  wire [1:0]  _slots_34_io_out_uop_iw_state;
  wire        _slots_34_io_out_uop_iw_p1_poisoned;
  wire        _slots_34_io_out_uop_iw_p2_poisoned;
  wire        _slots_34_io_out_uop_is_br;
  wire        _slots_34_io_out_uop_is_jalr;
  wire        _slots_34_io_out_uop_is_jal;
  wire        _slots_34_io_out_uop_is_sfb;
  wire [19:0] _slots_34_io_out_uop_br_mask;
  wire [4:0]  _slots_34_io_out_uop_br_tag;
  wire [5:0]  _slots_34_io_out_uop_ftq_idx;
  wire        _slots_34_io_out_uop_edge_inst;
  wire [5:0]  _slots_34_io_out_uop_pc_lob;
  wire        _slots_34_io_out_uop_taken;
  wire [19:0] _slots_34_io_out_uop_imm_packed;
  wire [11:0] _slots_34_io_out_uop_csr_addr;
  wire [6:0]  _slots_34_io_out_uop_rob_idx;
  wire [4:0]  _slots_34_io_out_uop_ldq_idx;
  wire [4:0]  _slots_34_io_out_uop_stq_idx;
  wire [1:0]  _slots_34_io_out_uop_rxq_idx;
  wire [6:0]  _slots_34_io_out_uop_pdst;
  wire [6:0]  _slots_34_io_out_uop_prs1;
  wire [6:0]  _slots_34_io_out_uop_prs2;
  wire [6:0]  _slots_34_io_out_uop_prs3;
  wire [5:0]  _slots_34_io_out_uop_ppred;
  wire        _slots_34_io_out_uop_prs1_busy;
  wire        _slots_34_io_out_uop_prs2_busy;
  wire        _slots_34_io_out_uop_prs3_busy;
  wire        _slots_34_io_out_uop_ppred_busy;
  wire [6:0]  _slots_34_io_out_uop_stale_pdst;
  wire        _slots_34_io_out_uop_exception;
  wire [63:0] _slots_34_io_out_uop_exc_cause;
  wire        _slots_34_io_out_uop_bypassable;
  wire [4:0]  _slots_34_io_out_uop_mem_cmd;
  wire [1:0]  _slots_34_io_out_uop_mem_size;
  wire        _slots_34_io_out_uop_mem_signed;
  wire        _slots_34_io_out_uop_is_fence;
  wire        _slots_34_io_out_uop_is_fencei;
  wire        _slots_34_io_out_uop_is_amo;
  wire        _slots_34_io_out_uop_uses_ldq;
  wire        _slots_34_io_out_uop_uses_stq;
  wire        _slots_34_io_out_uop_is_sys_pc2epc;
  wire        _slots_34_io_out_uop_is_unique;
  wire        _slots_34_io_out_uop_flush_on_commit;
  wire        _slots_34_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_34_io_out_uop_ldst;
  wire [5:0]  _slots_34_io_out_uop_lrs1;
  wire [5:0]  _slots_34_io_out_uop_lrs2;
  wire [5:0]  _slots_34_io_out_uop_lrs3;
  wire        _slots_34_io_out_uop_ldst_val;
  wire [1:0]  _slots_34_io_out_uop_dst_rtype;
  wire [1:0]  _slots_34_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_34_io_out_uop_lrs2_rtype;
  wire        _slots_34_io_out_uop_frs3_en;
  wire        _slots_34_io_out_uop_fp_val;
  wire        _slots_34_io_out_uop_fp_single;
  wire        _slots_34_io_out_uop_xcpt_pf_if;
  wire        _slots_34_io_out_uop_xcpt_ae_if;
  wire        _slots_34_io_out_uop_xcpt_ma_if;
  wire        _slots_34_io_out_uop_bp_debug_if;
  wire        _slots_34_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_34_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_34_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_34_io_uop_uopc;
  wire [31:0] _slots_34_io_uop_inst;
  wire [31:0] _slots_34_io_uop_debug_inst;
  wire        _slots_34_io_uop_is_rvc;
  wire [39:0] _slots_34_io_uop_debug_pc;
  wire [2:0]  _slots_34_io_uop_iq_type;
  wire [9:0]  _slots_34_io_uop_fu_code;
  wire [1:0]  _slots_34_io_uop_iw_state;
  wire        _slots_34_io_uop_iw_p1_poisoned;
  wire        _slots_34_io_uop_iw_p2_poisoned;
  wire        _slots_34_io_uop_is_br;
  wire        _slots_34_io_uop_is_jalr;
  wire        _slots_34_io_uop_is_jal;
  wire        _slots_34_io_uop_is_sfb;
  wire [19:0] _slots_34_io_uop_br_mask;
  wire [4:0]  _slots_34_io_uop_br_tag;
  wire [5:0]  _slots_34_io_uop_ftq_idx;
  wire        _slots_34_io_uop_edge_inst;
  wire [5:0]  _slots_34_io_uop_pc_lob;
  wire        _slots_34_io_uop_taken;
  wire [19:0] _slots_34_io_uop_imm_packed;
  wire [11:0] _slots_34_io_uop_csr_addr;
  wire [6:0]  _slots_34_io_uop_rob_idx;
  wire [4:0]  _slots_34_io_uop_ldq_idx;
  wire [4:0]  _slots_34_io_uop_stq_idx;
  wire [1:0]  _slots_34_io_uop_rxq_idx;
  wire [6:0]  _slots_34_io_uop_pdst;
  wire [6:0]  _slots_34_io_uop_prs1;
  wire [6:0]  _slots_34_io_uop_prs2;
  wire [6:0]  _slots_34_io_uop_prs3;
  wire [5:0]  _slots_34_io_uop_ppred;
  wire        _slots_34_io_uop_prs1_busy;
  wire        _slots_34_io_uop_prs2_busy;
  wire        _slots_34_io_uop_prs3_busy;
  wire        _slots_34_io_uop_ppred_busy;
  wire [6:0]  _slots_34_io_uop_stale_pdst;
  wire        _slots_34_io_uop_exception;
  wire [63:0] _slots_34_io_uop_exc_cause;
  wire        _slots_34_io_uop_bypassable;
  wire [4:0]  _slots_34_io_uop_mem_cmd;
  wire [1:0]  _slots_34_io_uop_mem_size;
  wire        _slots_34_io_uop_mem_signed;
  wire        _slots_34_io_uop_is_fence;
  wire        _slots_34_io_uop_is_fencei;
  wire        _slots_34_io_uop_is_amo;
  wire        _slots_34_io_uop_uses_ldq;
  wire        _slots_34_io_uop_uses_stq;
  wire        _slots_34_io_uop_is_sys_pc2epc;
  wire        _slots_34_io_uop_is_unique;
  wire        _slots_34_io_uop_flush_on_commit;
  wire        _slots_34_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_34_io_uop_ldst;
  wire [5:0]  _slots_34_io_uop_lrs1;
  wire [5:0]  _slots_34_io_uop_lrs2;
  wire [5:0]  _slots_34_io_uop_lrs3;
  wire        _slots_34_io_uop_ldst_val;
  wire [1:0]  _slots_34_io_uop_dst_rtype;
  wire [1:0]  _slots_34_io_uop_lrs1_rtype;
  wire [1:0]  _slots_34_io_uop_lrs2_rtype;
  wire        _slots_34_io_uop_frs3_en;
  wire        _slots_34_io_uop_fp_val;
  wire        _slots_34_io_uop_fp_single;
  wire        _slots_34_io_uop_xcpt_pf_if;
  wire        _slots_34_io_uop_xcpt_ae_if;
  wire        _slots_34_io_uop_xcpt_ma_if;
  wire        _slots_34_io_uop_bp_debug_if;
  wire        _slots_34_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_34_io_uop_debug_fsrc;
  wire [1:0]  _slots_34_io_uop_debug_tsrc;
  wire        _slots_33_io_valid;
  wire        _slots_33_io_will_be_valid;
  wire        _slots_33_io_request;
  wire [6:0]  _slots_33_io_out_uop_uopc;
  wire [31:0] _slots_33_io_out_uop_inst;
  wire [31:0] _slots_33_io_out_uop_debug_inst;
  wire        _slots_33_io_out_uop_is_rvc;
  wire [39:0] _slots_33_io_out_uop_debug_pc;
  wire [2:0]  _slots_33_io_out_uop_iq_type;
  wire [9:0]  _slots_33_io_out_uop_fu_code;
  wire [1:0]  _slots_33_io_out_uop_iw_state;
  wire        _slots_33_io_out_uop_iw_p1_poisoned;
  wire        _slots_33_io_out_uop_iw_p2_poisoned;
  wire        _slots_33_io_out_uop_is_br;
  wire        _slots_33_io_out_uop_is_jalr;
  wire        _slots_33_io_out_uop_is_jal;
  wire        _slots_33_io_out_uop_is_sfb;
  wire [19:0] _slots_33_io_out_uop_br_mask;
  wire [4:0]  _slots_33_io_out_uop_br_tag;
  wire [5:0]  _slots_33_io_out_uop_ftq_idx;
  wire        _slots_33_io_out_uop_edge_inst;
  wire [5:0]  _slots_33_io_out_uop_pc_lob;
  wire        _slots_33_io_out_uop_taken;
  wire [19:0] _slots_33_io_out_uop_imm_packed;
  wire [11:0] _slots_33_io_out_uop_csr_addr;
  wire [6:0]  _slots_33_io_out_uop_rob_idx;
  wire [4:0]  _slots_33_io_out_uop_ldq_idx;
  wire [4:0]  _slots_33_io_out_uop_stq_idx;
  wire [1:0]  _slots_33_io_out_uop_rxq_idx;
  wire [6:0]  _slots_33_io_out_uop_pdst;
  wire [6:0]  _slots_33_io_out_uop_prs1;
  wire [6:0]  _slots_33_io_out_uop_prs2;
  wire [6:0]  _slots_33_io_out_uop_prs3;
  wire [5:0]  _slots_33_io_out_uop_ppred;
  wire        _slots_33_io_out_uop_prs1_busy;
  wire        _slots_33_io_out_uop_prs2_busy;
  wire        _slots_33_io_out_uop_prs3_busy;
  wire        _slots_33_io_out_uop_ppred_busy;
  wire [6:0]  _slots_33_io_out_uop_stale_pdst;
  wire        _slots_33_io_out_uop_exception;
  wire [63:0] _slots_33_io_out_uop_exc_cause;
  wire        _slots_33_io_out_uop_bypassable;
  wire [4:0]  _slots_33_io_out_uop_mem_cmd;
  wire [1:0]  _slots_33_io_out_uop_mem_size;
  wire        _slots_33_io_out_uop_mem_signed;
  wire        _slots_33_io_out_uop_is_fence;
  wire        _slots_33_io_out_uop_is_fencei;
  wire        _slots_33_io_out_uop_is_amo;
  wire        _slots_33_io_out_uop_uses_ldq;
  wire        _slots_33_io_out_uop_uses_stq;
  wire        _slots_33_io_out_uop_is_sys_pc2epc;
  wire        _slots_33_io_out_uop_is_unique;
  wire        _slots_33_io_out_uop_flush_on_commit;
  wire        _slots_33_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_33_io_out_uop_ldst;
  wire [5:0]  _slots_33_io_out_uop_lrs1;
  wire [5:0]  _slots_33_io_out_uop_lrs2;
  wire [5:0]  _slots_33_io_out_uop_lrs3;
  wire        _slots_33_io_out_uop_ldst_val;
  wire [1:0]  _slots_33_io_out_uop_dst_rtype;
  wire [1:0]  _slots_33_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_33_io_out_uop_lrs2_rtype;
  wire        _slots_33_io_out_uop_frs3_en;
  wire        _slots_33_io_out_uop_fp_val;
  wire        _slots_33_io_out_uop_fp_single;
  wire        _slots_33_io_out_uop_xcpt_pf_if;
  wire        _slots_33_io_out_uop_xcpt_ae_if;
  wire        _slots_33_io_out_uop_xcpt_ma_if;
  wire        _slots_33_io_out_uop_bp_debug_if;
  wire        _slots_33_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_33_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_33_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_33_io_uop_uopc;
  wire [31:0] _slots_33_io_uop_inst;
  wire [31:0] _slots_33_io_uop_debug_inst;
  wire        _slots_33_io_uop_is_rvc;
  wire [39:0] _slots_33_io_uop_debug_pc;
  wire [2:0]  _slots_33_io_uop_iq_type;
  wire [9:0]  _slots_33_io_uop_fu_code;
  wire [1:0]  _slots_33_io_uop_iw_state;
  wire        _slots_33_io_uop_iw_p1_poisoned;
  wire        _slots_33_io_uop_iw_p2_poisoned;
  wire        _slots_33_io_uop_is_br;
  wire        _slots_33_io_uop_is_jalr;
  wire        _slots_33_io_uop_is_jal;
  wire        _slots_33_io_uop_is_sfb;
  wire [19:0] _slots_33_io_uop_br_mask;
  wire [4:0]  _slots_33_io_uop_br_tag;
  wire [5:0]  _slots_33_io_uop_ftq_idx;
  wire        _slots_33_io_uop_edge_inst;
  wire [5:0]  _slots_33_io_uop_pc_lob;
  wire        _slots_33_io_uop_taken;
  wire [19:0] _slots_33_io_uop_imm_packed;
  wire [11:0] _slots_33_io_uop_csr_addr;
  wire [6:0]  _slots_33_io_uop_rob_idx;
  wire [4:0]  _slots_33_io_uop_ldq_idx;
  wire [4:0]  _slots_33_io_uop_stq_idx;
  wire [1:0]  _slots_33_io_uop_rxq_idx;
  wire [6:0]  _slots_33_io_uop_pdst;
  wire [6:0]  _slots_33_io_uop_prs1;
  wire [6:0]  _slots_33_io_uop_prs2;
  wire [6:0]  _slots_33_io_uop_prs3;
  wire [5:0]  _slots_33_io_uop_ppred;
  wire        _slots_33_io_uop_prs1_busy;
  wire        _slots_33_io_uop_prs2_busy;
  wire        _slots_33_io_uop_prs3_busy;
  wire        _slots_33_io_uop_ppred_busy;
  wire [6:0]  _slots_33_io_uop_stale_pdst;
  wire        _slots_33_io_uop_exception;
  wire [63:0] _slots_33_io_uop_exc_cause;
  wire        _slots_33_io_uop_bypassable;
  wire [4:0]  _slots_33_io_uop_mem_cmd;
  wire [1:0]  _slots_33_io_uop_mem_size;
  wire        _slots_33_io_uop_mem_signed;
  wire        _slots_33_io_uop_is_fence;
  wire        _slots_33_io_uop_is_fencei;
  wire        _slots_33_io_uop_is_amo;
  wire        _slots_33_io_uop_uses_ldq;
  wire        _slots_33_io_uop_uses_stq;
  wire        _slots_33_io_uop_is_sys_pc2epc;
  wire        _slots_33_io_uop_is_unique;
  wire        _slots_33_io_uop_flush_on_commit;
  wire        _slots_33_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_33_io_uop_ldst;
  wire [5:0]  _slots_33_io_uop_lrs1;
  wire [5:0]  _slots_33_io_uop_lrs2;
  wire [5:0]  _slots_33_io_uop_lrs3;
  wire        _slots_33_io_uop_ldst_val;
  wire [1:0]  _slots_33_io_uop_dst_rtype;
  wire [1:0]  _slots_33_io_uop_lrs1_rtype;
  wire [1:0]  _slots_33_io_uop_lrs2_rtype;
  wire        _slots_33_io_uop_frs3_en;
  wire        _slots_33_io_uop_fp_val;
  wire        _slots_33_io_uop_fp_single;
  wire        _slots_33_io_uop_xcpt_pf_if;
  wire        _slots_33_io_uop_xcpt_ae_if;
  wire        _slots_33_io_uop_xcpt_ma_if;
  wire        _slots_33_io_uop_bp_debug_if;
  wire        _slots_33_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_33_io_uop_debug_fsrc;
  wire [1:0]  _slots_33_io_uop_debug_tsrc;
  wire        _slots_32_io_valid;
  wire        _slots_32_io_will_be_valid;
  wire        _slots_32_io_request;
  wire [6:0]  _slots_32_io_out_uop_uopc;
  wire [31:0] _slots_32_io_out_uop_inst;
  wire [31:0] _slots_32_io_out_uop_debug_inst;
  wire        _slots_32_io_out_uop_is_rvc;
  wire [39:0] _slots_32_io_out_uop_debug_pc;
  wire [2:0]  _slots_32_io_out_uop_iq_type;
  wire [9:0]  _slots_32_io_out_uop_fu_code;
  wire [1:0]  _slots_32_io_out_uop_iw_state;
  wire        _slots_32_io_out_uop_iw_p1_poisoned;
  wire        _slots_32_io_out_uop_iw_p2_poisoned;
  wire        _slots_32_io_out_uop_is_br;
  wire        _slots_32_io_out_uop_is_jalr;
  wire        _slots_32_io_out_uop_is_jal;
  wire        _slots_32_io_out_uop_is_sfb;
  wire [19:0] _slots_32_io_out_uop_br_mask;
  wire [4:0]  _slots_32_io_out_uop_br_tag;
  wire [5:0]  _slots_32_io_out_uop_ftq_idx;
  wire        _slots_32_io_out_uop_edge_inst;
  wire [5:0]  _slots_32_io_out_uop_pc_lob;
  wire        _slots_32_io_out_uop_taken;
  wire [19:0] _slots_32_io_out_uop_imm_packed;
  wire [11:0] _slots_32_io_out_uop_csr_addr;
  wire [6:0]  _slots_32_io_out_uop_rob_idx;
  wire [4:0]  _slots_32_io_out_uop_ldq_idx;
  wire [4:0]  _slots_32_io_out_uop_stq_idx;
  wire [1:0]  _slots_32_io_out_uop_rxq_idx;
  wire [6:0]  _slots_32_io_out_uop_pdst;
  wire [6:0]  _slots_32_io_out_uop_prs1;
  wire [6:0]  _slots_32_io_out_uop_prs2;
  wire [6:0]  _slots_32_io_out_uop_prs3;
  wire [5:0]  _slots_32_io_out_uop_ppred;
  wire        _slots_32_io_out_uop_prs1_busy;
  wire        _slots_32_io_out_uop_prs2_busy;
  wire        _slots_32_io_out_uop_prs3_busy;
  wire        _slots_32_io_out_uop_ppred_busy;
  wire [6:0]  _slots_32_io_out_uop_stale_pdst;
  wire        _slots_32_io_out_uop_exception;
  wire [63:0] _slots_32_io_out_uop_exc_cause;
  wire        _slots_32_io_out_uop_bypassable;
  wire [4:0]  _slots_32_io_out_uop_mem_cmd;
  wire [1:0]  _slots_32_io_out_uop_mem_size;
  wire        _slots_32_io_out_uop_mem_signed;
  wire        _slots_32_io_out_uop_is_fence;
  wire        _slots_32_io_out_uop_is_fencei;
  wire        _slots_32_io_out_uop_is_amo;
  wire        _slots_32_io_out_uop_uses_ldq;
  wire        _slots_32_io_out_uop_uses_stq;
  wire        _slots_32_io_out_uop_is_sys_pc2epc;
  wire        _slots_32_io_out_uop_is_unique;
  wire        _slots_32_io_out_uop_flush_on_commit;
  wire        _slots_32_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_32_io_out_uop_ldst;
  wire [5:0]  _slots_32_io_out_uop_lrs1;
  wire [5:0]  _slots_32_io_out_uop_lrs2;
  wire [5:0]  _slots_32_io_out_uop_lrs3;
  wire        _slots_32_io_out_uop_ldst_val;
  wire [1:0]  _slots_32_io_out_uop_dst_rtype;
  wire [1:0]  _slots_32_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_32_io_out_uop_lrs2_rtype;
  wire        _slots_32_io_out_uop_frs3_en;
  wire        _slots_32_io_out_uop_fp_val;
  wire        _slots_32_io_out_uop_fp_single;
  wire        _slots_32_io_out_uop_xcpt_pf_if;
  wire        _slots_32_io_out_uop_xcpt_ae_if;
  wire        _slots_32_io_out_uop_xcpt_ma_if;
  wire        _slots_32_io_out_uop_bp_debug_if;
  wire        _slots_32_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_32_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_32_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_32_io_uop_uopc;
  wire [31:0] _slots_32_io_uop_inst;
  wire [31:0] _slots_32_io_uop_debug_inst;
  wire        _slots_32_io_uop_is_rvc;
  wire [39:0] _slots_32_io_uop_debug_pc;
  wire [2:0]  _slots_32_io_uop_iq_type;
  wire [9:0]  _slots_32_io_uop_fu_code;
  wire [1:0]  _slots_32_io_uop_iw_state;
  wire        _slots_32_io_uop_iw_p1_poisoned;
  wire        _slots_32_io_uop_iw_p2_poisoned;
  wire        _slots_32_io_uop_is_br;
  wire        _slots_32_io_uop_is_jalr;
  wire        _slots_32_io_uop_is_jal;
  wire        _slots_32_io_uop_is_sfb;
  wire [19:0] _slots_32_io_uop_br_mask;
  wire [4:0]  _slots_32_io_uop_br_tag;
  wire [5:0]  _slots_32_io_uop_ftq_idx;
  wire        _slots_32_io_uop_edge_inst;
  wire [5:0]  _slots_32_io_uop_pc_lob;
  wire        _slots_32_io_uop_taken;
  wire [19:0] _slots_32_io_uop_imm_packed;
  wire [11:0] _slots_32_io_uop_csr_addr;
  wire [6:0]  _slots_32_io_uop_rob_idx;
  wire [4:0]  _slots_32_io_uop_ldq_idx;
  wire [4:0]  _slots_32_io_uop_stq_idx;
  wire [1:0]  _slots_32_io_uop_rxq_idx;
  wire [6:0]  _slots_32_io_uop_pdst;
  wire [6:0]  _slots_32_io_uop_prs1;
  wire [6:0]  _slots_32_io_uop_prs2;
  wire [6:0]  _slots_32_io_uop_prs3;
  wire [5:0]  _slots_32_io_uop_ppred;
  wire        _slots_32_io_uop_prs1_busy;
  wire        _slots_32_io_uop_prs2_busy;
  wire        _slots_32_io_uop_prs3_busy;
  wire        _slots_32_io_uop_ppred_busy;
  wire [6:0]  _slots_32_io_uop_stale_pdst;
  wire        _slots_32_io_uop_exception;
  wire [63:0] _slots_32_io_uop_exc_cause;
  wire        _slots_32_io_uop_bypassable;
  wire [4:0]  _slots_32_io_uop_mem_cmd;
  wire [1:0]  _slots_32_io_uop_mem_size;
  wire        _slots_32_io_uop_mem_signed;
  wire        _slots_32_io_uop_is_fence;
  wire        _slots_32_io_uop_is_fencei;
  wire        _slots_32_io_uop_is_amo;
  wire        _slots_32_io_uop_uses_ldq;
  wire        _slots_32_io_uop_uses_stq;
  wire        _slots_32_io_uop_is_sys_pc2epc;
  wire        _slots_32_io_uop_is_unique;
  wire        _slots_32_io_uop_flush_on_commit;
  wire        _slots_32_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_32_io_uop_ldst;
  wire [5:0]  _slots_32_io_uop_lrs1;
  wire [5:0]  _slots_32_io_uop_lrs2;
  wire [5:0]  _slots_32_io_uop_lrs3;
  wire        _slots_32_io_uop_ldst_val;
  wire [1:0]  _slots_32_io_uop_dst_rtype;
  wire [1:0]  _slots_32_io_uop_lrs1_rtype;
  wire [1:0]  _slots_32_io_uop_lrs2_rtype;
  wire        _slots_32_io_uop_frs3_en;
  wire        _slots_32_io_uop_fp_val;
  wire        _slots_32_io_uop_fp_single;
  wire        _slots_32_io_uop_xcpt_pf_if;
  wire        _slots_32_io_uop_xcpt_ae_if;
  wire        _slots_32_io_uop_xcpt_ma_if;
  wire        _slots_32_io_uop_bp_debug_if;
  wire        _slots_32_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_32_io_uop_debug_fsrc;
  wire [1:0]  _slots_32_io_uop_debug_tsrc;
  wire        _slots_31_io_valid;
  wire        _slots_31_io_will_be_valid;
  wire        _slots_31_io_request;
  wire [6:0]  _slots_31_io_out_uop_uopc;
  wire [31:0] _slots_31_io_out_uop_inst;
  wire [31:0] _slots_31_io_out_uop_debug_inst;
  wire        _slots_31_io_out_uop_is_rvc;
  wire [39:0] _slots_31_io_out_uop_debug_pc;
  wire [2:0]  _slots_31_io_out_uop_iq_type;
  wire [9:0]  _slots_31_io_out_uop_fu_code;
  wire [1:0]  _slots_31_io_out_uop_iw_state;
  wire        _slots_31_io_out_uop_iw_p1_poisoned;
  wire        _slots_31_io_out_uop_iw_p2_poisoned;
  wire        _slots_31_io_out_uop_is_br;
  wire        _slots_31_io_out_uop_is_jalr;
  wire        _slots_31_io_out_uop_is_jal;
  wire        _slots_31_io_out_uop_is_sfb;
  wire [19:0] _slots_31_io_out_uop_br_mask;
  wire [4:0]  _slots_31_io_out_uop_br_tag;
  wire [5:0]  _slots_31_io_out_uop_ftq_idx;
  wire        _slots_31_io_out_uop_edge_inst;
  wire [5:0]  _slots_31_io_out_uop_pc_lob;
  wire        _slots_31_io_out_uop_taken;
  wire [19:0] _slots_31_io_out_uop_imm_packed;
  wire [11:0] _slots_31_io_out_uop_csr_addr;
  wire [6:0]  _slots_31_io_out_uop_rob_idx;
  wire [4:0]  _slots_31_io_out_uop_ldq_idx;
  wire [4:0]  _slots_31_io_out_uop_stq_idx;
  wire [1:0]  _slots_31_io_out_uop_rxq_idx;
  wire [6:0]  _slots_31_io_out_uop_pdst;
  wire [6:0]  _slots_31_io_out_uop_prs1;
  wire [6:0]  _slots_31_io_out_uop_prs2;
  wire [6:0]  _slots_31_io_out_uop_prs3;
  wire [5:0]  _slots_31_io_out_uop_ppred;
  wire        _slots_31_io_out_uop_prs1_busy;
  wire        _slots_31_io_out_uop_prs2_busy;
  wire        _slots_31_io_out_uop_prs3_busy;
  wire        _slots_31_io_out_uop_ppred_busy;
  wire [6:0]  _slots_31_io_out_uop_stale_pdst;
  wire        _slots_31_io_out_uop_exception;
  wire [63:0] _slots_31_io_out_uop_exc_cause;
  wire        _slots_31_io_out_uop_bypassable;
  wire [4:0]  _slots_31_io_out_uop_mem_cmd;
  wire [1:0]  _slots_31_io_out_uop_mem_size;
  wire        _slots_31_io_out_uop_mem_signed;
  wire        _slots_31_io_out_uop_is_fence;
  wire        _slots_31_io_out_uop_is_fencei;
  wire        _slots_31_io_out_uop_is_amo;
  wire        _slots_31_io_out_uop_uses_ldq;
  wire        _slots_31_io_out_uop_uses_stq;
  wire        _slots_31_io_out_uop_is_sys_pc2epc;
  wire        _slots_31_io_out_uop_is_unique;
  wire        _slots_31_io_out_uop_flush_on_commit;
  wire        _slots_31_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_31_io_out_uop_ldst;
  wire [5:0]  _slots_31_io_out_uop_lrs1;
  wire [5:0]  _slots_31_io_out_uop_lrs2;
  wire [5:0]  _slots_31_io_out_uop_lrs3;
  wire        _slots_31_io_out_uop_ldst_val;
  wire [1:0]  _slots_31_io_out_uop_dst_rtype;
  wire [1:0]  _slots_31_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_31_io_out_uop_lrs2_rtype;
  wire        _slots_31_io_out_uop_frs3_en;
  wire        _slots_31_io_out_uop_fp_val;
  wire        _slots_31_io_out_uop_fp_single;
  wire        _slots_31_io_out_uop_xcpt_pf_if;
  wire        _slots_31_io_out_uop_xcpt_ae_if;
  wire        _slots_31_io_out_uop_xcpt_ma_if;
  wire        _slots_31_io_out_uop_bp_debug_if;
  wire        _slots_31_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_31_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_31_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_31_io_uop_uopc;
  wire [31:0] _slots_31_io_uop_inst;
  wire [31:0] _slots_31_io_uop_debug_inst;
  wire        _slots_31_io_uop_is_rvc;
  wire [39:0] _slots_31_io_uop_debug_pc;
  wire [2:0]  _slots_31_io_uop_iq_type;
  wire [9:0]  _slots_31_io_uop_fu_code;
  wire [1:0]  _slots_31_io_uop_iw_state;
  wire        _slots_31_io_uop_iw_p1_poisoned;
  wire        _slots_31_io_uop_iw_p2_poisoned;
  wire        _slots_31_io_uop_is_br;
  wire        _slots_31_io_uop_is_jalr;
  wire        _slots_31_io_uop_is_jal;
  wire        _slots_31_io_uop_is_sfb;
  wire [19:0] _slots_31_io_uop_br_mask;
  wire [4:0]  _slots_31_io_uop_br_tag;
  wire [5:0]  _slots_31_io_uop_ftq_idx;
  wire        _slots_31_io_uop_edge_inst;
  wire [5:0]  _slots_31_io_uop_pc_lob;
  wire        _slots_31_io_uop_taken;
  wire [19:0] _slots_31_io_uop_imm_packed;
  wire [11:0] _slots_31_io_uop_csr_addr;
  wire [6:0]  _slots_31_io_uop_rob_idx;
  wire [4:0]  _slots_31_io_uop_ldq_idx;
  wire [4:0]  _slots_31_io_uop_stq_idx;
  wire [1:0]  _slots_31_io_uop_rxq_idx;
  wire [6:0]  _slots_31_io_uop_pdst;
  wire [6:0]  _slots_31_io_uop_prs1;
  wire [6:0]  _slots_31_io_uop_prs2;
  wire [6:0]  _slots_31_io_uop_prs3;
  wire [5:0]  _slots_31_io_uop_ppred;
  wire        _slots_31_io_uop_prs1_busy;
  wire        _slots_31_io_uop_prs2_busy;
  wire        _slots_31_io_uop_prs3_busy;
  wire        _slots_31_io_uop_ppred_busy;
  wire [6:0]  _slots_31_io_uop_stale_pdst;
  wire        _slots_31_io_uop_exception;
  wire [63:0] _slots_31_io_uop_exc_cause;
  wire        _slots_31_io_uop_bypassable;
  wire [4:0]  _slots_31_io_uop_mem_cmd;
  wire [1:0]  _slots_31_io_uop_mem_size;
  wire        _slots_31_io_uop_mem_signed;
  wire        _slots_31_io_uop_is_fence;
  wire        _slots_31_io_uop_is_fencei;
  wire        _slots_31_io_uop_is_amo;
  wire        _slots_31_io_uop_uses_ldq;
  wire        _slots_31_io_uop_uses_stq;
  wire        _slots_31_io_uop_is_sys_pc2epc;
  wire        _slots_31_io_uop_is_unique;
  wire        _slots_31_io_uop_flush_on_commit;
  wire        _slots_31_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_31_io_uop_ldst;
  wire [5:0]  _slots_31_io_uop_lrs1;
  wire [5:0]  _slots_31_io_uop_lrs2;
  wire [5:0]  _slots_31_io_uop_lrs3;
  wire        _slots_31_io_uop_ldst_val;
  wire [1:0]  _slots_31_io_uop_dst_rtype;
  wire [1:0]  _slots_31_io_uop_lrs1_rtype;
  wire [1:0]  _slots_31_io_uop_lrs2_rtype;
  wire        _slots_31_io_uop_frs3_en;
  wire        _slots_31_io_uop_fp_val;
  wire        _slots_31_io_uop_fp_single;
  wire        _slots_31_io_uop_xcpt_pf_if;
  wire        _slots_31_io_uop_xcpt_ae_if;
  wire        _slots_31_io_uop_xcpt_ma_if;
  wire        _slots_31_io_uop_bp_debug_if;
  wire        _slots_31_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_31_io_uop_debug_fsrc;
  wire [1:0]  _slots_31_io_uop_debug_tsrc;
  wire        _slots_30_io_valid;
  wire        _slots_30_io_will_be_valid;
  wire        _slots_30_io_request;
  wire [6:0]  _slots_30_io_out_uop_uopc;
  wire [31:0] _slots_30_io_out_uop_inst;
  wire [31:0] _slots_30_io_out_uop_debug_inst;
  wire        _slots_30_io_out_uop_is_rvc;
  wire [39:0] _slots_30_io_out_uop_debug_pc;
  wire [2:0]  _slots_30_io_out_uop_iq_type;
  wire [9:0]  _slots_30_io_out_uop_fu_code;
  wire [1:0]  _slots_30_io_out_uop_iw_state;
  wire        _slots_30_io_out_uop_iw_p1_poisoned;
  wire        _slots_30_io_out_uop_iw_p2_poisoned;
  wire        _slots_30_io_out_uop_is_br;
  wire        _slots_30_io_out_uop_is_jalr;
  wire        _slots_30_io_out_uop_is_jal;
  wire        _slots_30_io_out_uop_is_sfb;
  wire [19:0] _slots_30_io_out_uop_br_mask;
  wire [4:0]  _slots_30_io_out_uop_br_tag;
  wire [5:0]  _slots_30_io_out_uop_ftq_idx;
  wire        _slots_30_io_out_uop_edge_inst;
  wire [5:0]  _slots_30_io_out_uop_pc_lob;
  wire        _slots_30_io_out_uop_taken;
  wire [19:0] _slots_30_io_out_uop_imm_packed;
  wire [11:0] _slots_30_io_out_uop_csr_addr;
  wire [6:0]  _slots_30_io_out_uop_rob_idx;
  wire [4:0]  _slots_30_io_out_uop_ldq_idx;
  wire [4:0]  _slots_30_io_out_uop_stq_idx;
  wire [1:0]  _slots_30_io_out_uop_rxq_idx;
  wire [6:0]  _slots_30_io_out_uop_pdst;
  wire [6:0]  _slots_30_io_out_uop_prs1;
  wire [6:0]  _slots_30_io_out_uop_prs2;
  wire [6:0]  _slots_30_io_out_uop_prs3;
  wire [5:0]  _slots_30_io_out_uop_ppred;
  wire        _slots_30_io_out_uop_prs1_busy;
  wire        _slots_30_io_out_uop_prs2_busy;
  wire        _slots_30_io_out_uop_prs3_busy;
  wire        _slots_30_io_out_uop_ppred_busy;
  wire [6:0]  _slots_30_io_out_uop_stale_pdst;
  wire        _slots_30_io_out_uop_exception;
  wire [63:0] _slots_30_io_out_uop_exc_cause;
  wire        _slots_30_io_out_uop_bypassable;
  wire [4:0]  _slots_30_io_out_uop_mem_cmd;
  wire [1:0]  _slots_30_io_out_uop_mem_size;
  wire        _slots_30_io_out_uop_mem_signed;
  wire        _slots_30_io_out_uop_is_fence;
  wire        _slots_30_io_out_uop_is_fencei;
  wire        _slots_30_io_out_uop_is_amo;
  wire        _slots_30_io_out_uop_uses_ldq;
  wire        _slots_30_io_out_uop_uses_stq;
  wire        _slots_30_io_out_uop_is_sys_pc2epc;
  wire        _slots_30_io_out_uop_is_unique;
  wire        _slots_30_io_out_uop_flush_on_commit;
  wire        _slots_30_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_30_io_out_uop_ldst;
  wire [5:0]  _slots_30_io_out_uop_lrs1;
  wire [5:0]  _slots_30_io_out_uop_lrs2;
  wire [5:0]  _slots_30_io_out_uop_lrs3;
  wire        _slots_30_io_out_uop_ldst_val;
  wire [1:0]  _slots_30_io_out_uop_dst_rtype;
  wire [1:0]  _slots_30_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_30_io_out_uop_lrs2_rtype;
  wire        _slots_30_io_out_uop_frs3_en;
  wire        _slots_30_io_out_uop_fp_val;
  wire        _slots_30_io_out_uop_fp_single;
  wire        _slots_30_io_out_uop_xcpt_pf_if;
  wire        _slots_30_io_out_uop_xcpt_ae_if;
  wire        _slots_30_io_out_uop_xcpt_ma_if;
  wire        _slots_30_io_out_uop_bp_debug_if;
  wire        _slots_30_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_30_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_30_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_30_io_uop_uopc;
  wire [31:0] _slots_30_io_uop_inst;
  wire [31:0] _slots_30_io_uop_debug_inst;
  wire        _slots_30_io_uop_is_rvc;
  wire [39:0] _slots_30_io_uop_debug_pc;
  wire [2:0]  _slots_30_io_uop_iq_type;
  wire [9:0]  _slots_30_io_uop_fu_code;
  wire [1:0]  _slots_30_io_uop_iw_state;
  wire        _slots_30_io_uop_iw_p1_poisoned;
  wire        _slots_30_io_uop_iw_p2_poisoned;
  wire        _slots_30_io_uop_is_br;
  wire        _slots_30_io_uop_is_jalr;
  wire        _slots_30_io_uop_is_jal;
  wire        _slots_30_io_uop_is_sfb;
  wire [19:0] _slots_30_io_uop_br_mask;
  wire [4:0]  _slots_30_io_uop_br_tag;
  wire [5:0]  _slots_30_io_uop_ftq_idx;
  wire        _slots_30_io_uop_edge_inst;
  wire [5:0]  _slots_30_io_uop_pc_lob;
  wire        _slots_30_io_uop_taken;
  wire [19:0] _slots_30_io_uop_imm_packed;
  wire [11:0] _slots_30_io_uop_csr_addr;
  wire [6:0]  _slots_30_io_uop_rob_idx;
  wire [4:0]  _slots_30_io_uop_ldq_idx;
  wire [4:0]  _slots_30_io_uop_stq_idx;
  wire [1:0]  _slots_30_io_uop_rxq_idx;
  wire [6:0]  _slots_30_io_uop_pdst;
  wire [6:0]  _slots_30_io_uop_prs1;
  wire [6:0]  _slots_30_io_uop_prs2;
  wire [6:0]  _slots_30_io_uop_prs3;
  wire [5:0]  _slots_30_io_uop_ppred;
  wire        _slots_30_io_uop_prs1_busy;
  wire        _slots_30_io_uop_prs2_busy;
  wire        _slots_30_io_uop_prs3_busy;
  wire        _slots_30_io_uop_ppred_busy;
  wire [6:0]  _slots_30_io_uop_stale_pdst;
  wire        _slots_30_io_uop_exception;
  wire [63:0] _slots_30_io_uop_exc_cause;
  wire        _slots_30_io_uop_bypassable;
  wire [4:0]  _slots_30_io_uop_mem_cmd;
  wire [1:0]  _slots_30_io_uop_mem_size;
  wire        _slots_30_io_uop_mem_signed;
  wire        _slots_30_io_uop_is_fence;
  wire        _slots_30_io_uop_is_fencei;
  wire        _slots_30_io_uop_is_amo;
  wire        _slots_30_io_uop_uses_ldq;
  wire        _slots_30_io_uop_uses_stq;
  wire        _slots_30_io_uop_is_sys_pc2epc;
  wire        _slots_30_io_uop_is_unique;
  wire        _slots_30_io_uop_flush_on_commit;
  wire        _slots_30_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_30_io_uop_ldst;
  wire [5:0]  _slots_30_io_uop_lrs1;
  wire [5:0]  _slots_30_io_uop_lrs2;
  wire [5:0]  _slots_30_io_uop_lrs3;
  wire        _slots_30_io_uop_ldst_val;
  wire [1:0]  _slots_30_io_uop_dst_rtype;
  wire [1:0]  _slots_30_io_uop_lrs1_rtype;
  wire [1:0]  _slots_30_io_uop_lrs2_rtype;
  wire        _slots_30_io_uop_frs3_en;
  wire        _slots_30_io_uop_fp_val;
  wire        _slots_30_io_uop_fp_single;
  wire        _slots_30_io_uop_xcpt_pf_if;
  wire        _slots_30_io_uop_xcpt_ae_if;
  wire        _slots_30_io_uop_xcpt_ma_if;
  wire        _slots_30_io_uop_bp_debug_if;
  wire        _slots_30_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_30_io_uop_debug_fsrc;
  wire [1:0]  _slots_30_io_uop_debug_tsrc;
  wire        _slots_29_io_valid;
  wire        _slots_29_io_will_be_valid;
  wire        _slots_29_io_request;
  wire [6:0]  _slots_29_io_out_uop_uopc;
  wire [31:0] _slots_29_io_out_uop_inst;
  wire [31:0] _slots_29_io_out_uop_debug_inst;
  wire        _slots_29_io_out_uop_is_rvc;
  wire [39:0] _slots_29_io_out_uop_debug_pc;
  wire [2:0]  _slots_29_io_out_uop_iq_type;
  wire [9:0]  _slots_29_io_out_uop_fu_code;
  wire [1:0]  _slots_29_io_out_uop_iw_state;
  wire        _slots_29_io_out_uop_iw_p1_poisoned;
  wire        _slots_29_io_out_uop_iw_p2_poisoned;
  wire        _slots_29_io_out_uop_is_br;
  wire        _slots_29_io_out_uop_is_jalr;
  wire        _slots_29_io_out_uop_is_jal;
  wire        _slots_29_io_out_uop_is_sfb;
  wire [19:0] _slots_29_io_out_uop_br_mask;
  wire [4:0]  _slots_29_io_out_uop_br_tag;
  wire [5:0]  _slots_29_io_out_uop_ftq_idx;
  wire        _slots_29_io_out_uop_edge_inst;
  wire [5:0]  _slots_29_io_out_uop_pc_lob;
  wire        _slots_29_io_out_uop_taken;
  wire [19:0] _slots_29_io_out_uop_imm_packed;
  wire [11:0] _slots_29_io_out_uop_csr_addr;
  wire [6:0]  _slots_29_io_out_uop_rob_idx;
  wire [4:0]  _slots_29_io_out_uop_ldq_idx;
  wire [4:0]  _slots_29_io_out_uop_stq_idx;
  wire [1:0]  _slots_29_io_out_uop_rxq_idx;
  wire [6:0]  _slots_29_io_out_uop_pdst;
  wire [6:0]  _slots_29_io_out_uop_prs1;
  wire [6:0]  _slots_29_io_out_uop_prs2;
  wire [6:0]  _slots_29_io_out_uop_prs3;
  wire [5:0]  _slots_29_io_out_uop_ppred;
  wire        _slots_29_io_out_uop_prs1_busy;
  wire        _slots_29_io_out_uop_prs2_busy;
  wire        _slots_29_io_out_uop_prs3_busy;
  wire        _slots_29_io_out_uop_ppred_busy;
  wire [6:0]  _slots_29_io_out_uop_stale_pdst;
  wire        _slots_29_io_out_uop_exception;
  wire [63:0] _slots_29_io_out_uop_exc_cause;
  wire        _slots_29_io_out_uop_bypassable;
  wire [4:0]  _slots_29_io_out_uop_mem_cmd;
  wire [1:0]  _slots_29_io_out_uop_mem_size;
  wire        _slots_29_io_out_uop_mem_signed;
  wire        _slots_29_io_out_uop_is_fence;
  wire        _slots_29_io_out_uop_is_fencei;
  wire        _slots_29_io_out_uop_is_amo;
  wire        _slots_29_io_out_uop_uses_ldq;
  wire        _slots_29_io_out_uop_uses_stq;
  wire        _slots_29_io_out_uop_is_sys_pc2epc;
  wire        _slots_29_io_out_uop_is_unique;
  wire        _slots_29_io_out_uop_flush_on_commit;
  wire        _slots_29_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_29_io_out_uop_ldst;
  wire [5:0]  _slots_29_io_out_uop_lrs1;
  wire [5:0]  _slots_29_io_out_uop_lrs2;
  wire [5:0]  _slots_29_io_out_uop_lrs3;
  wire        _slots_29_io_out_uop_ldst_val;
  wire [1:0]  _slots_29_io_out_uop_dst_rtype;
  wire [1:0]  _slots_29_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_29_io_out_uop_lrs2_rtype;
  wire        _slots_29_io_out_uop_frs3_en;
  wire        _slots_29_io_out_uop_fp_val;
  wire        _slots_29_io_out_uop_fp_single;
  wire        _slots_29_io_out_uop_xcpt_pf_if;
  wire        _slots_29_io_out_uop_xcpt_ae_if;
  wire        _slots_29_io_out_uop_xcpt_ma_if;
  wire        _slots_29_io_out_uop_bp_debug_if;
  wire        _slots_29_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_29_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_29_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_29_io_uop_uopc;
  wire [31:0] _slots_29_io_uop_inst;
  wire [31:0] _slots_29_io_uop_debug_inst;
  wire        _slots_29_io_uop_is_rvc;
  wire [39:0] _slots_29_io_uop_debug_pc;
  wire [2:0]  _slots_29_io_uop_iq_type;
  wire [9:0]  _slots_29_io_uop_fu_code;
  wire [1:0]  _slots_29_io_uop_iw_state;
  wire        _slots_29_io_uop_iw_p1_poisoned;
  wire        _slots_29_io_uop_iw_p2_poisoned;
  wire        _slots_29_io_uop_is_br;
  wire        _slots_29_io_uop_is_jalr;
  wire        _slots_29_io_uop_is_jal;
  wire        _slots_29_io_uop_is_sfb;
  wire [19:0] _slots_29_io_uop_br_mask;
  wire [4:0]  _slots_29_io_uop_br_tag;
  wire [5:0]  _slots_29_io_uop_ftq_idx;
  wire        _slots_29_io_uop_edge_inst;
  wire [5:0]  _slots_29_io_uop_pc_lob;
  wire        _slots_29_io_uop_taken;
  wire [19:0] _slots_29_io_uop_imm_packed;
  wire [11:0] _slots_29_io_uop_csr_addr;
  wire [6:0]  _slots_29_io_uop_rob_idx;
  wire [4:0]  _slots_29_io_uop_ldq_idx;
  wire [4:0]  _slots_29_io_uop_stq_idx;
  wire [1:0]  _slots_29_io_uop_rxq_idx;
  wire [6:0]  _slots_29_io_uop_pdst;
  wire [6:0]  _slots_29_io_uop_prs1;
  wire [6:0]  _slots_29_io_uop_prs2;
  wire [6:0]  _slots_29_io_uop_prs3;
  wire [5:0]  _slots_29_io_uop_ppred;
  wire        _slots_29_io_uop_prs1_busy;
  wire        _slots_29_io_uop_prs2_busy;
  wire        _slots_29_io_uop_prs3_busy;
  wire        _slots_29_io_uop_ppred_busy;
  wire [6:0]  _slots_29_io_uop_stale_pdst;
  wire        _slots_29_io_uop_exception;
  wire [63:0] _slots_29_io_uop_exc_cause;
  wire        _slots_29_io_uop_bypassable;
  wire [4:0]  _slots_29_io_uop_mem_cmd;
  wire [1:0]  _slots_29_io_uop_mem_size;
  wire        _slots_29_io_uop_mem_signed;
  wire        _slots_29_io_uop_is_fence;
  wire        _slots_29_io_uop_is_fencei;
  wire        _slots_29_io_uop_is_amo;
  wire        _slots_29_io_uop_uses_ldq;
  wire        _slots_29_io_uop_uses_stq;
  wire        _slots_29_io_uop_is_sys_pc2epc;
  wire        _slots_29_io_uop_is_unique;
  wire        _slots_29_io_uop_flush_on_commit;
  wire        _slots_29_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_29_io_uop_ldst;
  wire [5:0]  _slots_29_io_uop_lrs1;
  wire [5:0]  _slots_29_io_uop_lrs2;
  wire [5:0]  _slots_29_io_uop_lrs3;
  wire        _slots_29_io_uop_ldst_val;
  wire [1:0]  _slots_29_io_uop_dst_rtype;
  wire [1:0]  _slots_29_io_uop_lrs1_rtype;
  wire [1:0]  _slots_29_io_uop_lrs2_rtype;
  wire        _slots_29_io_uop_frs3_en;
  wire        _slots_29_io_uop_fp_val;
  wire        _slots_29_io_uop_fp_single;
  wire        _slots_29_io_uop_xcpt_pf_if;
  wire        _slots_29_io_uop_xcpt_ae_if;
  wire        _slots_29_io_uop_xcpt_ma_if;
  wire        _slots_29_io_uop_bp_debug_if;
  wire        _slots_29_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_29_io_uop_debug_fsrc;
  wire [1:0]  _slots_29_io_uop_debug_tsrc;
  wire        _slots_28_io_valid;
  wire        _slots_28_io_will_be_valid;
  wire        _slots_28_io_request;
  wire [6:0]  _slots_28_io_out_uop_uopc;
  wire [31:0] _slots_28_io_out_uop_inst;
  wire [31:0] _slots_28_io_out_uop_debug_inst;
  wire        _slots_28_io_out_uop_is_rvc;
  wire [39:0] _slots_28_io_out_uop_debug_pc;
  wire [2:0]  _slots_28_io_out_uop_iq_type;
  wire [9:0]  _slots_28_io_out_uop_fu_code;
  wire [1:0]  _slots_28_io_out_uop_iw_state;
  wire        _slots_28_io_out_uop_iw_p1_poisoned;
  wire        _slots_28_io_out_uop_iw_p2_poisoned;
  wire        _slots_28_io_out_uop_is_br;
  wire        _slots_28_io_out_uop_is_jalr;
  wire        _slots_28_io_out_uop_is_jal;
  wire        _slots_28_io_out_uop_is_sfb;
  wire [19:0] _slots_28_io_out_uop_br_mask;
  wire [4:0]  _slots_28_io_out_uop_br_tag;
  wire [5:0]  _slots_28_io_out_uop_ftq_idx;
  wire        _slots_28_io_out_uop_edge_inst;
  wire [5:0]  _slots_28_io_out_uop_pc_lob;
  wire        _slots_28_io_out_uop_taken;
  wire [19:0] _slots_28_io_out_uop_imm_packed;
  wire [11:0] _slots_28_io_out_uop_csr_addr;
  wire [6:0]  _slots_28_io_out_uop_rob_idx;
  wire [4:0]  _slots_28_io_out_uop_ldq_idx;
  wire [4:0]  _slots_28_io_out_uop_stq_idx;
  wire [1:0]  _slots_28_io_out_uop_rxq_idx;
  wire [6:0]  _slots_28_io_out_uop_pdst;
  wire [6:0]  _slots_28_io_out_uop_prs1;
  wire [6:0]  _slots_28_io_out_uop_prs2;
  wire [6:0]  _slots_28_io_out_uop_prs3;
  wire [5:0]  _slots_28_io_out_uop_ppred;
  wire        _slots_28_io_out_uop_prs1_busy;
  wire        _slots_28_io_out_uop_prs2_busy;
  wire        _slots_28_io_out_uop_prs3_busy;
  wire        _slots_28_io_out_uop_ppred_busy;
  wire [6:0]  _slots_28_io_out_uop_stale_pdst;
  wire        _slots_28_io_out_uop_exception;
  wire [63:0] _slots_28_io_out_uop_exc_cause;
  wire        _slots_28_io_out_uop_bypassable;
  wire [4:0]  _slots_28_io_out_uop_mem_cmd;
  wire [1:0]  _slots_28_io_out_uop_mem_size;
  wire        _slots_28_io_out_uop_mem_signed;
  wire        _slots_28_io_out_uop_is_fence;
  wire        _slots_28_io_out_uop_is_fencei;
  wire        _slots_28_io_out_uop_is_amo;
  wire        _slots_28_io_out_uop_uses_ldq;
  wire        _slots_28_io_out_uop_uses_stq;
  wire        _slots_28_io_out_uop_is_sys_pc2epc;
  wire        _slots_28_io_out_uop_is_unique;
  wire        _slots_28_io_out_uop_flush_on_commit;
  wire        _slots_28_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_28_io_out_uop_ldst;
  wire [5:0]  _slots_28_io_out_uop_lrs1;
  wire [5:0]  _slots_28_io_out_uop_lrs2;
  wire [5:0]  _slots_28_io_out_uop_lrs3;
  wire        _slots_28_io_out_uop_ldst_val;
  wire [1:0]  _slots_28_io_out_uop_dst_rtype;
  wire [1:0]  _slots_28_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_28_io_out_uop_lrs2_rtype;
  wire        _slots_28_io_out_uop_frs3_en;
  wire        _slots_28_io_out_uop_fp_val;
  wire        _slots_28_io_out_uop_fp_single;
  wire        _slots_28_io_out_uop_xcpt_pf_if;
  wire        _slots_28_io_out_uop_xcpt_ae_if;
  wire        _slots_28_io_out_uop_xcpt_ma_if;
  wire        _slots_28_io_out_uop_bp_debug_if;
  wire        _slots_28_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_28_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_28_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_28_io_uop_uopc;
  wire [31:0] _slots_28_io_uop_inst;
  wire [31:0] _slots_28_io_uop_debug_inst;
  wire        _slots_28_io_uop_is_rvc;
  wire [39:0] _slots_28_io_uop_debug_pc;
  wire [2:0]  _slots_28_io_uop_iq_type;
  wire [9:0]  _slots_28_io_uop_fu_code;
  wire [1:0]  _slots_28_io_uop_iw_state;
  wire        _slots_28_io_uop_iw_p1_poisoned;
  wire        _slots_28_io_uop_iw_p2_poisoned;
  wire        _slots_28_io_uop_is_br;
  wire        _slots_28_io_uop_is_jalr;
  wire        _slots_28_io_uop_is_jal;
  wire        _slots_28_io_uop_is_sfb;
  wire [19:0] _slots_28_io_uop_br_mask;
  wire [4:0]  _slots_28_io_uop_br_tag;
  wire [5:0]  _slots_28_io_uop_ftq_idx;
  wire        _slots_28_io_uop_edge_inst;
  wire [5:0]  _slots_28_io_uop_pc_lob;
  wire        _slots_28_io_uop_taken;
  wire [19:0] _slots_28_io_uop_imm_packed;
  wire [11:0] _slots_28_io_uop_csr_addr;
  wire [6:0]  _slots_28_io_uop_rob_idx;
  wire [4:0]  _slots_28_io_uop_ldq_idx;
  wire [4:0]  _slots_28_io_uop_stq_idx;
  wire [1:0]  _slots_28_io_uop_rxq_idx;
  wire [6:0]  _slots_28_io_uop_pdst;
  wire [6:0]  _slots_28_io_uop_prs1;
  wire [6:0]  _slots_28_io_uop_prs2;
  wire [6:0]  _slots_28_io_uop_prs3;
  wire [5:0]  _slots_28_io_uop_ppred;
  wire        _slots_28_io_uop_prs1_busy;
  wire        _slots_28_io_uop_prs2_busy;
  wire        _slots_28_io_uop_prs3_busy;
  wire        _slots_28_io_uop_ppred_busy;
  wire [6:0]  _slots_28_io_uop_stale_pdst;
  wire        _slots_28_io_uop_exception;
  wire [63:0] _slots_28_io_uop_exc_cause;
  wire        _slots_28_io_uop_bypassable;
  wire [4:0]  _slots_28_io_uop_mem_cmd;
  wire [1:0]  _slots_28_io_uop_mem_size;
  wire        _slots_28_io_uop_mem_signed;
  wire        _slots_28_io_uop_is_fence;
  wire        _slots_28_io_uop_is_fencei;
  wire        _slots_28_io_uop_is_amo;
  wire        _slots_28_io_uop_uses_ldq;
  wire        _slots_28_io_uop_uses_stq;
  wire        _slots_28_io_uop_is_sys_pc2epc;
  wire        _slots_28_io_uop_is_unique;
  wire        _slots_28_io_uop_flush_on_commit;
  wire        _slots_28_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_28_io_uop_ldst;
  wire [5:0]  _slots_28_io_uop_lrs1;
  wire [5:0]  _slots_28_io_uop_lrs2;
  wire [5:0]  _slots_28_io_uop_lrs3;
  wire        _slots_28_io_uop_ldst_val;
  wire [1:0]  _slots_28_io_uop_dst_rtype;
  wire [1:0]  _slots_28_io_uop_lrs1_rtype;
  wire [1:0]  _slots_28_io_uop_lrs2_rtype;
  wire        _slots_28_io_uop_frs3_en;
  wire        _slots_28_io_uop_fp_val;
  wire        _slots_28_io_uop_fp_single;
  wire        _slots_28_io_uop_xcpt_pf_if;
  wire        _slots_28_io_uop_xcpt_ae_if;
  wire        _slots_28_io_uop_xcpt_ma_if;
  wire        _slots_28_io_uop_bp_debug_if;
  wire        _slots_28_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_28_io_uop_debug_fsrc;
  wire [1:0]  _slots_28_io_uop_debug_tsrc;
  wire        _slots_27_io_valid;
  wire        _slots_27_io_will_be_valid;
  wire        _slots_27_io_request;
  wire [6:0]  _slots_27_io_out_uop_uopc;
  wire [31:0] _slots_27_io_out_uop_inst;
  wire [31:0] _slots_27_io_out_uop_debug_inst;
  wire        _slots_27_io_out_uop_is_rvc;
  wire [39:0] _slots_27_io_out_uop_debug_pc;
  wire [2:0]  _slots_27_io_out_uop_iq_type;
  wire [9:0]  _slots_27_io_out_uop_fu_code;
  wire [1:0]  _slots_27_io_out_uop_iw_state;
  wire        _slots_27_io_out_uop_iw_p1_poisoned;
  wire        _slots_27_io_out_uop_iw_p2_poisoned;
  wire        _slots_27_io_out_uop_is_br;
  wire        _slots_27_io_out_uop_is_jalr;
  wire        _slots_27_io_out_uop_is_jal;
  wire        _slots_27_io_out_uop_is_sfb;
  wire [19:0] _slots_27_io_out_uop_br_mask;
  wire [4:0]  _slots_27_io_out_uop_br_tag;
  wire [5:0]  _slots_27_io_out_uop_ftq_idx;
  wire        _slots_27_io_out_uop_edge_inst;
  wire [5:0]  _slots_27_io_out_uop_pc_lob;
  wire        _slots_27_io_out_uop_taken;
  wire [19:0] _slots_27_io_out_uop_imm_packed;
  wire [11:0] _slots_27_io_out_uop_csr_addr;
  wire [6:0]  _slots_27_io_out_uop_rob_idx;
  wire [4:0]  _slots_27_io_out_uop_ldq_idx;
  wire [4:0]  _slots_27_io_out_uop_stq_idx;
  wire [1:0]  _slots_27_io_out_uop_rxq_idx;
  wire [6:0]  _slots_27_io_out_uop_pdst;
  wire [6:0]  _slots_27_io_out_uop_prs1;
  wire [6:0]  _slots_27_io_out_uop_prs2;
  wire [6:0]  _slots_27_io_out_uop_prs3;
  wire [5:0]  _slots_27_io_out_uop_ppred;
  wire        _slots_27_io_out_uop_prs1_busy;
  wire        _slots_27_io_out_uop_prs2_busy;
  wire        _slots_27_io_out_uop_prs3_busy;
  wire        _slots_27_io_out_uop_ppred_busy;
  wire [6:0]  _slots_27_io_out_uop_stale_pdst;
  wire        _slots_27_io_out_uop_exception;
  wire [63:0] _slots_27_io_out_uop_exc_cause;
  wire        _slots_27_io_out_uop_bypassable;
  wire [4:0]  _slots_27_io_out_uop_mem_cmd;
  wire [1:0]  _slots_27_io_out_uop_mem_size;
  wire        _slots_27_io_out_uop_mem_signed;
  wire        _slots_27_io_out_uop_is_fence;
  wire        _slots_27_io_out_uop_is_fencei;
  wire        _slots_27_io_out_uop_is_amo;
  wire        _slots_27_io_out_uop_uses_ldq;
  wire        _slots_27_io_out_uop_uses_stq;
  wire        _slots_27_io_out_uop_is_sys_pc2epc;
  wire        _slots_27_io_out_uop_is_unique;
  wire        _slots_27_io_out_uop_flush_on_commit;
  wire        _slots_27_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_27_io_out_uop_ldst;
  wire [5:0]  _slots_27_io_out_uop_lrs1;
  wire [5:0]  _slots_27_io_out_uop_lrs2;
  wire [5:0]  _slots_27_io_out_uop_lrs3;
  wire        _slots_27_io_out_uop_ldst_val;
  wire [1:0]  _slots_27_io_out_uop_dst_rtype;
  wire [1:0]  _slots_27_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_27_io_out_uop_lrs2_rtype;
  wire        _slots_27_io_out_uop_frs3_en;
  wire        _slots_27_io_out_uop_fp_val;
  wire        _slots_27_io_out_uop_fp_single;
  wire        _slots_27_io_out_uop_xcpt_pf_if;
  wire        _slots_27_io_out_uop_xcpt_ae_if;
  wire        _slots_27_io_out_uop_xcpt_ma_if;
  wire        _slots_27_io_out_uop_bp_debug_if;
  wire        _slots_27_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_27_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_27_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_27_io_uop_uopc;
  wire [31:0] _slots_27_io_uop_inst;
  wire [31:0] _slots_27_io_uop_debug_inst;
  wire        _slots_27_io_uop_is_rvc;
  wire [39:0] _slots_27_io_uop_debug_pc;
  wire [2:0]  _slots_27_io_uop_iq_type;
  wire [9:0]  _slots_27_io_uop_fu_code;
  wire [1:0]  _slots_27_io_uop_iw_state;
  wire        _slots_27_io_uop_iw_p1_poisoned;
  wire        _slots_27_io_uop_iw_p2_poisoned;
  wire        _slots_27_io_uop_is_br;
  wire        _slots_27_io_uop_is_jalr;
  wire        _slots_27_io_uop_is_jal;
  wire        _slots_27_io_uop_is_sfb;
  wire [19:0] _slots_27_io_uop_br_mask;
  wire [4:0]  _slots_27_io_uop_br_tag;
  wire [5:0]  _slots_27_io_uop_ftq_idx;
  wire        _slots_27_io_uop_edge_inst;
  wire [5:0]  _slots_27_io_uop_pc_lob;
  wire        _slots_27_io_uop_taken;
  wire [19:0] _slots_27_io_uop_imm_packed;
  wire [11:0] _slots_27_io_uop_csr_addr;
  wire [6:0]  _slots_27_io_uop_rob_idx;
  wire [4:0]  _slots_27_io_uop_ldq_idx;
  wire [4:0]  _slots_27_io_uop_stq_idx;
  wire [1:0]  _slots_27_io_uop_rxq_idx;
  wire [6:0]  _slots_27_io_uop_pdst;
  wire [6:0]  _slots_27_io_uop_prs1;
  wire [6:0]  _slots_27_io_uop_prs2;
  wire [6:0]  _slots_27_io_uop_prs3;
  wire [5:0]  _slots_27_io_uop_ppred;
  wire        _slots_27_io_uop_prs1_busy;
  wire        _slots_27_io_uop_prs2_busy;
  wire        _slots_27_io_uop_prs3_busy;
  wire        _slots_27_io_uop_ppred_busy;
  wire [6:0]  _slots_27_io_uop_stale_pdst;
  wire        _slots_27_io_uop_exception;
  wire [63:0] _slots_27_io_uop_exc_cause;
  wire        _slots_27_io_uop_bypassable;
  wire [4:0]  _slots_27_io_uop_mem_cmd;
  wire [1:0]  _slots_27_io_uop_mem_size;
  wire        _slots_27_io_uop_mem_signed;
  wire        _slots_27_io_uop_is_fence;
  wire        _slots_27_io_uop_is_fencei;
  wire        _slots_27_io_uop_is_amo;
  wire        _slots_27_io_uop_uses_ldq;
  wire        _slots_27_io_uop_uses_stq;
  wire        _slots_27_io_uop_is_sys_pc2epc;
  wire        _slots_27_io_uop_is_unique;
  wire        _slots_27_io_uop_flush_on_commit;
  wire        _slots_27_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_27_io_uop_ldst;
  wire [5:0]  _slots_27_io_uop_lrs1;
  wire [5:0]  _slots_27_io_uop_lrs2;
  wire [5:0]  _slots_27_io_uop_lrs3;
  wire        _slots_27_io_uop_ldst_val;
  wire [1:0]  _slots_27_io_uop_dst_rtype;
  wire [1:0]  _slots_27_io_uop_lrs1_rtype;
  wire [1:0]  _slots_27_io_uop_lrs2_rtype;
  wire        _slots_27_io_uop_frs3_en;
  wire        _slots_27_io_uop_fp_val;
  wire        _slots_27_io_uop_fp_single;
  wire        _slots_27_io_uop_xcpt_pf_if;
  wire        _slots_27_io_uop_xcpt_ae_if;
  wire        _slots_27_io_uop_xcpt_ma_if;
  wire        _slots_27_io_uop_bp_debug_if;
  wire        _slots_27_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_27_io_uop_debug_fsrc;
  wire [1:0]  _slots_27_io_uop_debug_tsrc;
  wire        _slots_26_io_valid;
  wire        _slots_26_io_will_be_valid;
  wire        _slots_26_io_request;
  wire [6:0]  _slots_26_io_out_uop_uopc;
  wire [31:0] _slots_26_io_out_uop_inst;
  wire [31:0] _slots_26_io_out_uop_debug_inst;
  wire        _slots_26_io_out_uop_is_rvc;
  wire [39:0] _slots_26_io_out_uop_debug_pc;
  wire [2:0]  _slots_26_io_out_uop_iq_type;
  wire [9:0]  _slots_26_io_out_uop_fu_code;
  wire [1:0]  _slots_26_io_out_uop_iw_state;
  wire        _slots_26_io_out_uop_iw_p1_poisoned;
  wire        _slots_26_io_out_uop_iw_p2_poisoned;
  wire        _slots_26_io_out_uop_is_br;
  wire        _slots_26_io_out_uop_is_jalr;
  wire        _slots_26_io_out_uop_is_jal;
  wire        _slots_26_io_out_uop_is_sfb;
  wire [19:0] _slots_26_io_out_uop_br_mask;
  wire [4:0]  _slots_26_io_out_uop_br_tag;
  wire [5:0]  _slots_26_io_out_uop_ftq_idx;
  wire        _slots_26_io_out_uop_edge_inst;
  wire [5:0]  _slots_26_io_out_uop_pc_lob;
  wire        _slots_26_io_out_uop_taken;
  wire [19:0] _slots_26_io_out_uop_imm_packed;
  wire [11:0] _slots_26_io_out_uop_csr_addr;
  wire [6:0]  _slots_26_io_out_uop_rob_idx;
  wire [4:0]  _slots_26_io_out_uop_ldq_idx;
  wire [4:0]  _slots_26_io_out_uop_stq_idx;
  wire [1:0]  _slots_26_io_out_uop_rxq_idx;
  wire [6:0]  _slots_26_io_out_uop_pdst;
  wire [6:0]  _slots_26_io_out_uop_prs1;
  wire [6:0]  _slots_26_io_out_uop_prs2;
  wire [6:0]  _slots_26_io_out_uop_prs3;
  wire [5:0]  _slots_26_io_out_uop_ppred;
  wire        _slots_26_io_out_uop_prs1_busy;
  wire        _slots_26_io_out_uop_prs2_busy;
  wire        _slots_26_io_out_uop_prs3_busy;
  wire        _slots_26_io_out_uop_ppred_busy;
  wire [6:0]  _slots_26_io_out_uop_stale_pdst;
  wire        _slots_26_io_out_uop_exception;
  wire [63:0] _slots_26_io_out_uop_exc_cause;
  wire        _slots_26_io_out_uop_bypassable;
  wire [4:0]  _slots_26_io_out_uop_mem_cmd;
  wire [1:0]  _slots_26_io_out_uop_mem_size;
  wire        _slots_26_io_out_uop_mem_signed;
  wire        _slots_26_io_out_uop_is_fence;
  wire        _slots_26_io_out_uop_is_fencei;
  wire        _slots_26_io_out_uop_is_amo;
  wire        _slots_26_io_out_uop_uses_ldq;
  wire        _slots_26_io_out_uop_uses_stq;
  wire        _slots_26_io_out_uop_is_sys_pc2epc;
  wire        _slots_26_io_out_uop_is_unique;
  wire        _slots_26_io_out_uop_flush_on_commit;
  wire        _slots_26_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_26_io_out_uop_ldst;
  wire [5:0]  _slots_26_io_out_uop_lrs1;
  wire [5:0]  _slots_26_io_out_uop_lrs2;
  wire [5:0]  _slots_26_io_out_uop_lrs3;
  wire        _slots_26_io_out_uop_ldst_val;
  wire [1:0]  _slots_26_io_out_uop_dst_rtype;
  wire [1:0]  _slots_26_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_26_io_out_uop_lrs2_rtype;
  wire        _slots_26_io_out_uop_frs3_en;
  wire        _slots_26_io_out_uop_fp_val;
  wire        _slots_26_io_out_uop_fp_single;
  wire        _slots_26_io_out_uop_xcpt_pf_if;
  wire        _slots_26_io_out_uop_xcpt_ae_if;
  wire        _slots_26_io_out_uop_xcpt_ma_if;
  wire        _slots_26_io_out_uop_bp_debug_if;
  wire        _slots_26_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_26_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_26_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_26_io_uop_uopc;
  wire [31:0] _slots_26_io_uop_inst;
  wire [31:0] _slots_26_io_uop_debug_inst;
  wire        _slots_26_io_uop_is_rvc;
  wire [39:0] _slots_26_io_uop_debug_pc;
  wire [2:0]  _slots_26_io_uop_iq_type;
  wire [9:0]  _slots_26_io_uop_fu_code;
  wire [1:0]  _slots_26_io_uop_iw_state;
  wire        _slots_26_io_uop_iw_p1_poisoned;
  wire        _slots_26_io_uop_iw_p2_poisoned;
  wire        _slots_26_io_uop_is_br;
  wire        _slots_26_io_uop_is_jalr;
  wire        _slots_26_io_uop_is_jal;
  wire        _slots_26_io_uop_is_sfb;
  wire [19:0] _slots_26_io_uop_br_mask;
  wire [4:0]  _slots_26_io_uop_br_tag;
  wire [5:0]  _slots_26_io_uop_ftq_idx;
  wire        _slots_26_io_uop_edge_inst;
  wire [5:0]  _slots_26_io_uop_pc_lob;
  wire        _slots_26_io_uop_taken;
  wire [19:0] _slots_26_io_uop_imm_packed;
  wire [11:0] _slots_26_io_uop_csr_addr;
  wire [6:0]  _slots_26_io_uop_rob_idx;
  wire [4:0]  _slots_26_io_uop_ldq_idx;
  wire [4:0]  _slots_26_io_uop_stq_idx;
  wire [1:0]  _slots_26_io_uop_rxq_idx;
  wire [6:0]  _slots_26_io_uop_pdst;
  wire [6:0]  _slots_26_io_uop_prs1;
  wire [6:0]  _slots_26_io_uop_prs2;
  wire [6:0]  _slots_26_io_uop_prs3;
  wire [5:0]  _slots_26_io_uop_ppred;
  wire        _slots_26_io_uop_prs1_busy;
  wire        _slots_26_io_uop_prs2_busy;
  wire        _slots_26_io_uop_prs3_busy;
  wire        _slots_26_io_uop_ppred_busy;
  wire [6:0]  _slots_26_io_uop_stale_pdst;
  wire        _slots_26_io_uop_exception;
  wire [63:0] _slots_26_io_uop_exc_cause;
  wire        _slots_26_io_uop_bypassable;
  wire [4:0]  _slots_26_io_uop_mem_cmd;
  wire [1:0]  _slots_26_io_uop_mem_size;
  wire        _slots_26_io_uop_mem_signed;
  wire        _slots_26_io_uop_is_fence;
  wire        _slots_26_io_uop_is_fencei;
  wire        _slots_26_io_uop_is_amo;
  wire        _slots_26_io_uop_uses_ldq;
  wire        _slots_26_io_uop_uses_stq;
  wire        _slots_26_io_uop_is_sys_pc2epc;
  wire        _slots_26_io_uop_is_unique;
  wire        _slots_26_io_uop_flush_on_commit;
  wire        _slots_26_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_26_io_uop_ldst;
  wire [5:0]  _slots_26_io_uop_lrs1;
  wire [5:0]  _slots_26_io_uop_lrs2;
  wire [5:0]  _slots_26_io_uop_lrs3;
  wire        _slots_26_io_uop_ldst_val;
  wire [1:0]  _slots_26_io_uop_dst_rtype;
  wire [1:0]  _slots_26_io_uop_lrs1_rtype;
  wire [1:0]  _slots_26_io_uop_lrs2_rtype;
  wire        _slots_26_io_uop_frs3_en;
  wire        _slots_26_io_uop_fp_val;
  wire        _slots_26_io_uop_fp_single;
  wire        _slots_26_io_uop_xcpt_pf_if;
  wire        _slots_26_io_uop_xcpt_ae_if;
  wire        _slots_26_io_uop_xcpt_ma_if;
  wire        _slots_26_io_uop_bp_debug_if;
  wire        _slots_26_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_26_io_uop_debug_fsrc;
  wire [1:0]  _slots_26_io_uop_debug_tsrc;
  wire        _slots_25_io_valid;
  wire        _slots_25_io_will_be_valid;
  wire        _slots_25_io_request;
  wire [6:0]  _slots_25_io_out_uop_uopc;
  wire [31:0] _slots_25_io_out_uop_inst;
  wire [31:0] _slots_25_io_out_uop_debug_inst;
  wire        _slots_25_io_out_uop_is_rvc;
  wire [39:0] _slots_25_io_out_uop_debug_pc;
  wire [2:0]  _slots_25_io_out_uop_iq_type;
  wire [9:0]  _slots_25_io_out_uop_fu_code;
  wire [1:0]  _slots_25_io_out_uop_iw_state;
  wire        _slots_25_io_out_uop_iw_p1_poisoned;
  wire        _slots_25_io_out_uop_iw_p2_poisoned;
  wire        _slots_25_io_out_uop_is_br;
  wire        _slots_25_io_out_uop_is_jalr;
  wire        _slots_25_io_out_uop_is_jal;
  wire        _slots_25_io_out_uop_is_sfb;
  wire [19:0] _slots_25_io_out_uop_br_mask;
  wire [4:0]  _slots_25_io_out_uop_br_tag;
  wire [5:0]  _slots_25_io_out_uop_ftq_idx;
  wire        _slots_25_io_out_uop_edge_inst;
  wire [5:0]  _slots_25_io_out_uop_pc_lob;
  wire        _slots_25_io_out_uop_taken;
  wire [19:0] _slots_25_io_out_uop_imm_packed;
  wire [11:0] _slots_25_io_out_uop_csr_addr;
  wire [6:0]  _slots_25_io_out_uop_rob_idx;
  wire [4:0]  _slots_25_io_out_uop_ldq_idx;
  wire [4:0]  _slots_25_io_out_uop_stq_idx;
  wire [1:0]  _slots_25_io_out_uop_rxq_idx;
  wire [6:0]  _slots_25_io_out_uop_pdst;
  wire [6:0]  _slots_25_io_out_uop_prs1;
  wire [6:0]  _slots_25_io_out_uop_prs2;
  wire [6:0]  _slots_25_io_out_uop_prs3;
  wire [5:0]  _slots_25_io_out_uop_ppred;
  wire        _slots_25_io_out_uop_prs1_busy;
  wire        _slots_25_io_out_uop_prs2_busy;
  wire        _slots_25_io_out_uop_prs3_busy;
  wire        _slots_25_io_out_uop_ppred_busy;
  wire [6:0]  _slots_25_io_out_uop_stale_pdst;
  wire        _slots_25_io_out_uop_exception;
  wire [63:0] _slots_25_io_out_uop_exc_cause;
  wire        _slots_25_io_out_uop_bypassable;
  wire [4:0]  _slots_25_io_out_uop_mem_cmd;
  wire [1:0]  _slots_25_io_out_uop_mem_size;
  wire        _slots_25_io_out_uop_mem_signed;
  wire        _slots_25_io_out_uop_is_fence;
  wire        _slots_25_io_out_uop_is_fencei;
  wire        _slots_25_io_out_uop_is_amo;
  wire        _slots_25_io_out_uop_uses_ldq;
  wire        _slots_25_io_out_uop_uses_stq;
  wire        _slots_25_io_out_uop_is_sys_pc2epc;
  wire        _slots_25_io_out_uop_is_unique;
  wire        _slots_25_io_out_uop_flush_on_commit;
  wire        _slots_25_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_25_io_out_uop_ldst;
  wire [5:0]  _slots_25_io_out_uop_lrs1;
  wire [5:0]  _slots_25_io_out_uop_lrs2;
  wire [5:0]  _slots_25_io_out_uop_lrs3;
  wire        _slots_25_io_out_uop_ldst_val;
  wire [1:0]  _slots_25_io_out_uop_dst_rtype;
  wire [1:0]  _slots_25_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_25_io_out_uop_lrs2_rtype;
  wire        _slots_25_io_out_uop_frs3_en;
  wire        _slots_25_io_out_uop_fp_val;
  wire        _slots_25_io_out_uop_fp_single;
  wire        _slots_25_io_out_uop_xcpt_pf_if;
  wire        _slots_25_io_out_uop_xcpt_ae_if;
  wire        _slots_25_io_out_uop_xcpt_ma_if;
  wire        _slots_25_io_out_uop_bp_debug_if;
  wire        _slots_25_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_25_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_25_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_25_io_uop_uopc;
  wire [31:0] _slots_25_io_uop_inst;
  wire [31:0] _slots_25_io_uop_debug_inst;
  wire        _slots_25_io_uop_is_rvc;
  wire [39:0] _slots_25_io_uop_debug_pc;
  wire [2:0]  _slots_25_io_uop_iq_type;
  wire [9:0]  _slots_25_io_uop_fu_code;
  wire [1:0]  _slots_25_io_uop_iw_state;
  wire        _slots_25_io_uop_iw_p1_poisoned;
  wire        _slots_25_io_uop_iw_p2_poisoned;
  wire        _slots_25_io_uop_is_br;
  wire        _slots_25_io_uop_is_jalr;
  wire        _slots_25_io_uop_is_jal;
  wire        _slots_25_io_uop_is_sfb;
  wire [19:0] _slots_25_io_uop_br_mask;
  wire [4:0]  _slots_25_io_uop_br_tag;
  wire [5:0]  _slots_25_io_uop_ftq_idx;
  wire        _slots_25_io_uop_edge_inst;
  wire [5:0]  _slots_25_io_uop_pc_lob;
  wire        _slots_25_io_uop_taken;
  wire [19:0] _slots_25_io_uop_imm_packed;
  wire [11:0] _slots_25_io_uop_csr_addr;
  wire [6:0]  _slots_25_io_uop_rob_idx;
  wire [4:0]  _slots_25_io_uop_ldq_idx;
  wire [4:0]  _slots_25_io_uop_stq_idx;
  wire [1:0]  _slots_25_io_uop_rxq_idx;
  wire [6:0]  _slots_25_io_uop_pdst;
  wire [6:0]  _slots_25_io_uop_prs1;
  wire [6:0]  _slots_25_io_uop_prs2;
  wire [6:0]  _slots_25_io_uop_prs3;
  wire [5:0]  _slots_25_io_uop_ppred;
  wire        _slots_25_io_uop_prs1_busy;
  wire        _slots_25_io_uop_prs2_busy;
  wire        _slots_25_io_uop_prs3_busy;
  wire        _slots_25_io_uop_ppred_busy;
  wire [6:0]  _slots_25_io_uop_stale_pdst;
  wire        _slots_25_io_uop_exception;
  wire [63:0] _slots_25_io_uop_exc_cause;
  wire        _slots_25_io_uop_bypassable;
  wire [4:0]  _slots_25_io_uop_mem_cmd;
  wire [1:0]  _slots_25_io_uop_mem_size;
  wire        _slots_25_io_uop_mem_signed;
  wire        _slots_25_io_uop_is_fence;
  wire        _slots_25_io_uop_is_fencei;
  wire        _slots_25_io_uop_is_amo;
  wire        _slots_25_io_uop_uses_ldq;
  wire        _slots_25_io_uop_uses_stq;
  wire        _slots_25_io_uop_is_sys_pc2epc;
  wire        _slots_25_io_uop_is_unique;
  wire        _slots_25_io_uop_flush_on_commit;
  wire        _slots_25_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_25_io_uop_ldst;
  wire [5:0]  _slots_25_io_uop_lrs1;
  wire [5:0]  _slots_25_io_uop_lrs2;
  wire [5:0]  _slots_25_io_uop_lrs3;
  wire        _slots_25_io_uop_ldst_val;
  wire [1:0]  _slots_25_io_uop_dst_rtype;
  wire [1:0]  _slots_25_io_uop_lrs1_rtype;
  wire [1:0]  _slots_25_io_uop_lrs2_rtype;
  wire        _slots_25_io_uop_frs3_en;
  wire        _slots_25_io_uop_fp_val;
  wire        _slots_25_io_uop_fp_single;
  wire        _slots_25_io_uop_xcpt_pf_if;
  wire        _slots_25_io_uop_xcpt_ae_if;
  wire        _slots_25_io_uop_xcpt_ma_if;
  wire        _slots_25_io_uop_bp_debug_if;
  wire        _slots_25_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_25_io_uop_debug_fsrc;
  wire [1:0]  _slots_25_io_uop_debug_tsrc;
  wire        _slots_24_io_valid;
  wire        _slots_24_io_will_be_valid;
  wire        _slots_24_io_request;
  wire [6:0]  _slots_24_io_out_uop_uopc;
  wire [31:0] _slots_24_io_out_uop_inst;
  wire [31:0] _slots_24_io_out_uop_debug_inst;
  wire        _slots_24_io_out_uop_is_rvc;
  wire [39:0] _slots_24_io_out_uop_debug_pc;
  wire [2:0]  _slots_24_io_out_uop_iq_type;
  wire [9:0]  _slots_24_io_out_uop_fu_code;
  wire [1:0]  _slots_24_io_out_uop_iw_state;
  wire        _slots_24_io_out_uop_iw_p1_poisoned;
  wire        _slots_24_io_out_uop_iw_p2_poisoned;
  wire        _slots_24_io_out_uop_is_br;
  wire        _slots_24_io_out_uop_is_jalr;
  wire        _slots_24_io_out_uop_is_jal;
  wire        _slots_24_io_out_uop_is_sfb;
  wire [19:0] _slots_24_io_out_uop_br_mask;
  wire [4:0]  _slots_24_io_out_uop_br_tag;
  wire [5:0]  _slots_24_io_out_uop_ftq_idx;
  wire        _slots_24_io_out_uop_edge_inst;
  wire [5:0]  _slots_24_io_out_uop_pc_lob;
  wire        _slots_24_io_out_uop_taken;
  wire [19:0] _slots_24_io_out_uop_imm_packed;
  wire [11:0] _slots_24_io_out_uop_csr_addr;
  wire [6:0]  _slots_24_io_out_uop_rob_idx;
  wire [4:0]  _slots_24_io_out_uop_ldq_idx;
  wire [4:0]  _slots_24_io_out_uop_stq_idx;
  wire [1:0]  _slots_24_io_out_uop_rxq_idx;
  wire [6:0]  _slots_24_io_out_uop_pdst;
  wire [6:0]  _slots_24_io_out_uop_prs1;
  wire [6:0]  _slots_24_io_out_uop_prs2;
  wire [6:0]  _slots_24_io_out_uop_prs3;
  wire [5:0]  _slots_24_io_out_uop_ppred;
  wire        _slots_24_io_out_uop_prs1_busy;
  wire        _slots_24_io_out_uop_prs2_busy;
  wire        _slots_24_io_out_uop_prs3_busy;
  wire        _slots_24_io_out_uop_ppred_busy;
  wire [6:0]  _slots_24_io_out_uop_stale_pdst;
  wire        _slots_24_io_out_uop_exception;
  wire [63:0] _slots_24_io_out_uop_exc_cause;
  wire        _slots_24_io_out_uop_bypassable;
  wire [4:0]  _slots_24_io_out_uop_mem_cmd;
  wire [1:0]  _slots_24_io_out_uop_mem_size;
  wire        _slots_24_io_out_uop_mem_signed;
  wire        _slots_24_io_out_uop_is_fence;
  wire        _slots_24_io_out_uop_is_fencei;
  wire        _slots_24_io_out_uop_is_amo;
  wire        _slots_24_io_out_uop_uses_ldq;
  wire        _slots_24_io_out_uop_uses_stq;
  wire        _slots_24_io_out_uop_is_sys_pc2epc;
  wire        _slots_24_io_out_uop_is_unique;
  wire        _slots_24_io_out_uop_flush_on_commit;
  wire        _slots_24_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_24_io_out_uop_ldst;
  wire [5:0]  _slots_24_io_out_uop_lrs1;
  wire [5:0]  _slots_24_io_out_uop_lrs2;
  wire [5:0]  _slots_24_io_out_uop_lrs3;
  wire        _slots_24_io_out_uop_ldst_val;
  wire [1:0]  _slots_24_io_out_uop_dst_rtype;
  wire [1:0]  _slots_24_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_24_io_out_uop_lrs2_rtype;
  wire        _slots_24_io_out_uop_frs3_en;
  wire        _slots_24_io_out_uop_fp_val;
  wire        _slots_24_io_out_uop_fp_single;
  wire        _slots_24_io_out_uop_xcpt_pf_if;
  wire        _slots_24_io_out_uop_xcpt_ae_if;
  wire        _slots_24_io_out_uop_xcpt_ma_if;
  wire        _slots_24_io_out_uop_bp_debug_if;
  wire        _slots_24_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_24_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_24_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_24_io_uop_uopc;
  wire [31:0] _slots_24_io_uop_inst;
  wire [31:0] _slots_24_io_uop_debug_inst;
  wire        _slots_24_io_uop_is_rvc;
  wire [39:0] _slots_24_io_uop_debug_pc;
  wire [2:0]  _slots_24_io_uop_iq_type;
  wire [9:0]  _slots_24_io_uop_fu_code;
  wire [1:0]  _slots_24_io_uop_iw_state;
  wire        _slots_24_io_uop_iw_p1_poisoned;
  wire        _slots_24_io_uop_iw_p2_poisoned;
  wire        _slots_24_io_uop_is_br;
  wire        _slots_24_io_uop_is_jalr;
  wire        _slots_24_io_uop_is_jal;
  wire        _slots_24_io_uop_is_sfb;
  wire [19:0] _slots_24_io_uop_br_mask;
  wire [4:0]  _slots_24_io_uop_br_tag;
  wire [5:0]  _slots_24_io_uop_ftq_idx;
  wire        _slots_24_io_uop_edge_inst;
  wire [5:0]  _slots_24_io_uop_pc_lob;
  wire        _slots_24_io_uop_taken;
  wire [19:0] _slots_24_io_uop_imm_packed;
  wire [11:0] _slots_24_io_uop_csr_addr;
  wire [6:0]  _slots_24_io_uop_rob_idx;
  wire [4:0]  _slots_24_io_uop_ldq_idx;
  wire [4:0]  _slots_24_io_uop_stq_idx;
  wire [1:0]  _slots_24_io_uop_rxq_idx;
  wire [6:0]  _slots_24_io_uop_pdst;
  wire [6:0]  _slots_24_io_uop_prs1;
  wire [6:0]  _slots_24_io_uop_prs2;
  wire [6:0]  _slots_24_io_uop_prs3;
  wire [5:0]  _slots_24_io_uop_ppred;
  wire        _slots_24_io_uop_prs1_busy;
  wire        _slots_24_io_uop_prs2_busy;
  wire        _slots_24_io_uop_prs3_busy;
  wire        _slots_24_io_uop_ppred_busy;
  wire [6:0]  _slots_24_io_uop_stale_pdst;
  wire        _slots_24_io_uop_exception;
  wire [63:0] _slots_24_io_uop_exc_cause;
  wire        _slots_24_io_uop_bypassable;
  wire [4:0]  _slots_24_io_uop_mem_cmd;
  wire [1:0]  _slots_24_io_uop_mem_size;
  wire        _slots_24_io_uop_mem_signed;
  wire        _slots_24_io_uop_is_fence;
  wire        _slots_24_io_uop_is_fencei;
  wire        _slots_24_io_uop_is_amo;
  wire        _slots_24_io_uop_uses_ldq;
  wire        _slots_24_io_uop_uses_stq;
  wire        _slots_24_io_uop_is_sys_pc2epc;
  wire        _slots_24_io_uop_is_unique;
  wire        _slots_24_io_uop_flush_on_commit;
  wire        _slots_24_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_24_io_uop_ldst;
  wire [5:0]  _slots_24_io_uop_lrs1;
  wire [5:0]  _slots_24_io_uop_lrs2;
  wire [5:0]  _slots_24_io_uop_lrs3;
  wire        _slots_24_io_uop_ldst_val;
  wire [1:0]  _slots_24_io_uop_dst_rtype;
  wire [1:0]  _slots_24_io_uop_lrs1_rtype;
  wire [1:0]  _slots_24_io_uop_lrs2_rtype;
  wire        _slots_24_io_uop_frs3_en;
  wire        _slots_24_io_uop_fp_val;
  wire        _slots_24_io_uop_fp_single;
  wire        _slots_24_io_uop_xcpt_pf_if;
  wire        _slots_24_io_uop_xcpt_ae_if;
  wire        _slots_24_io_uop_xcpt_ma_if;
  wire        _slots_24_io_uop_bp_debug_if;
  wire        _slots_24_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_24_io_uop_debug_fsrc;
  wire [1:0]  _slots_24_io_uop_debug_tsrc;
  wire        _slots_23_io_valid;
  wire        _slots_23_io_will_be_valid;
  wire        _slots_23_io_request;
  wire [6:0]  _slots_23_io_out_uop_uopc;
  wire [31:0] _slots_23_io_out_uop_inst;
  wire [31:0] _slots_23_io_out_uop_debug_inst;
  wire        _slots_23_io_out_uop_is_rvc;
  wire [39:0] _slots_23_io_out_uop_debug_pc;
  wire [2:0]  _slots_23_io_out_uop_iq_type;
  wire [9:0]  _slots_23_io_out_uop_fu_code;
  wire [1:0]  _slots_23_io_out_uop_iw_state;
  wire        _slots_23_io_out_uop_iw_p1_poisoned;
  wire        _slots_23_io_out_uop_iw_p2_poisoned;
  wire        _slots_23_io_out_uop_is_br;
  wire        _slots_23_io_out_uop_is_jalr;
  wire        _slots_23_io_out_uop_is_jal;
  wire        _slots_23_io_out_uop_is_sfb;
  wire [19:0] _slots_23_io_out_uop_br_mask;
  wire [4:0]  _slots_23_io_out_uop_br_tag;
  wire [5:0]  _slots_23_io_out_uop_ftq_idx;
  wire        _slots_23_io_out_uop_edge_inst;
  wire [5:0]  _slots_23_io_out_uop_pc_lob;
  wire        _slots_23_io_out_uop_taken;
  wire [19:0] _slots_23_io_out_uop_imm_packed;
  wire [11:0] _slots_23_io_out_uop_csr_addr;
  wire [6:0]  _slots_23_io_out_uop_rob_idx;
  wire [4:0]  _slots_23_io_out_uop_ldq_idx;
  wire [4:0]  _slots_23_io_out_uop_stq_idx;
  wire [1:0]  _slots_23_io_out_uop_rxq_idx;
  wire [6:0]  _slots_23_io_out_uop_pdst;
  wire [6:0]  _slots_23_io_out_uop_prs1;
  wire [6:0]  _slots_23_io_out_uop_prs2;
  wire [6:0]  _slots_23_io_out_uop_prs3;
  wire [5:0]  _slots_23_io_out_uop_ppred;
  wire        _slots_23_io_out_uop_prs1_busy;
  wire        _slots_23_io_out_uop_prs2_busy;
  wire        _slots_23_io_out_uop_prs3_busy;
  wire        _slots_23_io_out_uop_ppred_busy;
  wire [6:0]  _slots_23_io_out_uop_stale_pdst;
  wire        _slots_23_io_out_uop_exception;
  wire [63:0] _slots_23_io_out_uop_exc_cause;
  wire        _slots_23_io_out_uop_bypassable;
  wire [4:0]  _slots_23_io_out_uop_mem_cmd;
  wire [1:0]  _slots_23_io_out_uop_mem_size;
  wire        _slots_23_io_out_uop_mem_signed;
  wire        _slots_23_io_out_uop_is_fence;
  wire        _slots_23_io_out_uop_is_fencei;
  wire        _slots_23_io_out_uop_is_amo;
  wire        _slots_23_io_out_uop_uses_ldq;
  wire        _slots_23_io_out_uop_uses_stq;
  wire        _slots_23_io_out_uop_is_sys_pc2epc;
  wire        _slots_23_io_out_uop_is_unique;
  wire        _slots_23_io_out_uop_flush_on_commit;
  wire        _slots_23_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_23_io_out_uop_ldst;
  wire [5:0]  _slots_23_io_out_uop_lrs1;
  wire [5:0]  _slots_23_io_out_uop_lrs2;
  wire [5:0]  _slots_23_io_out_uop_lrs3;
  wire        _slots_23_io_out_uop_ldst_val;
  wire [1:0]  _slots_23_io_out_uop_dst_rtype;
  wire [1:0]  _slots_23_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_23_io_out_uop_lrs2_rtype;
  wire        _slots_23_io_out_uop_frs3_en;
  wire        _slots_23_io_out_uop_fp_val;
  wire        _slots_23_io_out_uop_fp_single;
  wire        _slots_23_io_out_uop_xcpt_pf_if;
  wire        _slots_23_io_out_uop_xcpt_ae_if;
  wire        _slots_23_io_out_uop_xcpt_ma_if;
  wire        _slots_23_io_out_uop_bp_debug_if;
  wire        _slots_23_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_23_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_23_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_23_io_uop_uopc;
  wire [31:0] _slots_23_io_uop_inst;
  wire [31:0] _slots_23_io_uop_debug_inst;
  wire        _slots_23_io_uop_is_rvc;
  wire [39:0] _slots_23_io_uop_debug_pc;
  wire [2:0]  _slots_23_io_uop_iq_type;
  wire [9:0]  _slots_23_io_uop_fu_code;
  wire [1:0]  _slots_23_io_uop_iw_state;
  wire        _slots_23_io_uop_iw_p1_poisoned;
  wire        _slots_23_io_uop_iw_p2_poisoned;
  wire        _slots_23_io_uop_is_br;
  wire        _slots_23_io_uop_is_jalr;
  wire        _slots_23_io_uop_is_jal;
  wire        _slots_23_io_uop_is_sfb;
  wire [19:0] _slots_23_io_uop_br_mask;
  wire [4:0]  _slots_23_io_uop_br_tag;
  wire [5:0]  _slots_23_io_uop_ftq_idx;
  wire        _slots_23_io_uop_edge_inst;
  wire [5:0]  _slots_23_io_uop_pc_lob;
  wire        _slots_23_io_uop_taken;
  wire [19:0] _slots_23_io_uop_imm_packed;
  wire [11:0] _slots_23_io_uop_csr_addr;
  wire [6:0]  _slots_23_io_uop_rob_idx;
  wire [4:0]  _slots_23_io_uop_ldq_idx;
  wire [4:0]  _slots_23_io_uop_stq_idx;
  wire [1:0]  _slots_23_io_uop_rxq_idx;
  wire [6:0]  _slots_23_io_uop_pdst;
  wire [6:0]  _slots_23_io_uop_prs1;
  wire [6:0]  _slots_23_io_uop_prs2;
  wire [6:0]  _slots_23_io_uop_prs3;
  wire [5:0]  _slots_23_io_uop_ppred;
  wire        _slots_23_io_uop_prs1_busy;
  wire        _slots_23_io_uop_prs2_busy;
  wire        _slots_23_io_uop_prs3_busy;
  wire        _slots_23_io_uop_ppred_busy;
  wire [6:0]  _slots_23_io_uop_stale_pdst;
  wire        _slots_23_io_uop_exception;
  wire [63:0] _slots_23_io_uop_exc_cause;
  wire        _slots_23_io_uop_bypassable;
  wire [4:0]  _slots_23_io_uop_mem_cmd;
  wire [1:0]  _slots_23_io_uop_mem_size;
  wire        _slots_23_io_uop_mem_signed;
  wire        _slots_23_io_uop_is_fence;
  wire        _slots_23_io_uop_is_fencei;
  wire        _slots_23_io_uop_is_amo;
  wire        _slots_23_io_uop_uses_ldq;
  wire        _slots_23_io_uop_uses_stq;
  wire        _slots_23_io_uop_is_sys_pc2epc;
  wire        _slots_23_io_uop_is_unique;
  wire        _slots_23_io_uop_flush_on_commit;
  wire        _slots_23_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_23_io_uop_ldst;
  wire [5:0]  _slots_23_io_uop_lrs1;
  wire [5:0]  _slots_23_io_uop_lrs2;
  wire [5:0]  _slots_23_io_uop_lrs3;
  wire        _slots_23_io_uop_ldst_val;
  wire [1:0]  _slots_23_io_uop_dst_rtype;
  wire [1:0]  _slots_23_io_uop_lrs1_rtype;
  wire [1:0]  _slots_23_io_uop_lrs2_rtype;
  wire        _slots_23_io_uop_frs3_en;
  wire        _slots_23_io_uop_fp_val;
  wire        _slots_23_io_uop_fp_single;
  wire        _slots_23_io_uop_xcpt_pf_if;
  wire        _slots_23_io_uop_xcpt_ae_if;
  wire        _slots_23_io_uop_xcpt_ma_if;
  wire        _slots_23_io_uop_bp_debug_if;
  wire        _slots_23_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_23_io_uop_debug_fsrc;
  wire [1:0]  _slots_23_io_uop_debug_tsrc;
  wire        _slots_22_io_valid;
  wire        _slots_22_io_will_be_valid;
  wire        _slots_22_io_request;
  wire [6:0]  _slots_22_io_out_uop_uopc;
  wire [31:0] _slots_22_io_out_uop_inst;
  wire [31:0] _slots_22_io_out_uop_debug_inst;
  wire        _slots_22_io_out_uop_is_rvc;
  wire [39:0] _slots_22_io_out_uop_debug_pc;
  wire [2:0]  _slots_22_io_out_uop_iq_type;
  wire [9:0]  _slots_22_io_out_uop_fu_code;
  wire [1:0]  _slots_22_io_out_uop_iw_state;
  wire        _slots_22_io_out_uop_iw_p1_poisoned;
  wire        _slots_22_io_out_uop_iw_p2_poisoned;
  wire        _slots_22_io_out_uop_is_br;
  wire        _slots_22_io_out_uop_is_jalr;
  wire        _slots_22_io_out_uop_is_jal;
  wire        _slots_22_io_out_uop_is_sfb;
  wire [19:0] _slots_22_io_out_uop_br_mask;
  wire [4:0]  _slots_22_io_out_uop_br_tag;
  wire [5:0]  _slots_22_io_out_uop_ftq_idx;
  wire        _slots_22_io_out_uop_edge_inst;
  wire [5:0]  _slots_22_io_out_uop_pc_lob;
  wire        _slots_22_io_out_uop_taken;
  wire [19:0] _slots_22_io_out_uop_imm_packed;
  wire [11:0] _slots_22_io_out_uop_csr_addr;
  wire [6:0]  _slots_22_io_out_uop_rob_idx;
  wire [4:0]  _slots_22_io_out_uop_ldq_idx;
  wire [4:0]  _slots_22_io_out_uop_stq_idx;
  wire [1:0]  _slots_22_io_out_uop_rxq_idx;
  wire [6:0]  _slots_22_io_out_uop_pdst;
  wire [6:0]  _slots_22_io_out_uop_prs1;
  wire [6:0]  _slots_22_io_out_uop_prs2;
  wire [6:0]  _slots_22_io_out_uop_prs3;
  wire [5:0]  _slots_22_io_out_uop_ppred;
  wire        _slots_22_io_out_uop_prs1_busy;
  wire        _slots_22_io_out_uop_prs2_busy;
  wire        _slots_22_io_out_uop_prs3_busy;
  wire        _slots_22_io_out_uop_ppred_busy;
  wire [6:0]  _slots_22_io_out_uop_stale_pdst;
  wire        _slots_22_io_out_uop_exception;
  wire [63:0] _slots_22_io_out_uop_exc_cause;
  wire        _slots_22_io_out_uop_bypassable;
  wire [4:0]  _slots_22_io_out_uop_mem_cmd;
  wire [1:0]  _slots_22_io_out_uop_mem_size;
  wire        _slots_22_io_out_uop_mem_signed;
  wire        _slots_22_io_out_uop_is_fence;
  wire        _slots_22_io_out_uop_is_fencei;
  wire        _slots_22_io_out_uop_is_amo;
  wire        _slots_22_io_out_uop_uses_ldq;
  wire        _slots_22_io_out_uop_uses_stq;
  wire        _slots_22_io_out_uop_is_sys_pc2epc;
  wire        _slots_22_io_out_uop_is_unique;
  wire        _slots_22_io_out_uop_flush_on_commit;
  wire        _slots_22_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_22_io_out_uop_ldst;
  wire [5:0]  _slots_22_io_out_uop_lrs1;
  wire [5:0]  _slots_22_io_out_uop_lrs2;
  wire [5:0]  _slots_22_io_out_uop_lrs3;
  wire        _slots_22_io_out_uop_ldst_val;
  wire [1:0]  _slots_22_io_out_uop_dst_rtype;
  wire [1:0]  _slots_22_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_22_io_out_uop_lrs2_rtype;
  wire        _slots_22_io_out_uop_frs3_en;
  wire        _slots_22_io_out_uop_fp_val;
  wire        _slots_22_io_out_uop_fp_single;
  wire        _slots_22_io_out_uop_xcpt_pf_if;
  wire        _slots_22_io_out_uop_xcpt_ae_if;
  wire        _slots_22_io_out_uop_xcpt_ma_if;
  wire        _slots_22_io_out_uop_bp_debug_if;
  wire        _slots_22_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_22_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_22_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_22_io_uop_uopc;
  wire [31:0] _slots_22_io_uop_inst;
  wire [31:0] _slots_22_io_uop_debug_inst;
  wire        _slots_22_io_uop_is_rvc;
  wire [39:0] _slots_22_io_uop_debug_pc;
  wire [2:0]  _slots_22_io_uop_iq_type;
  wire [9:0]  _slots_22_io_uop_fu_code;
  wire [1:0]  _slots_22_io_uop_iw_state;
  wire        _slots_22_io_uop_iw_p1_poisoned;
  wire        _slots_22_io_uop_iw_p2_poisoned;
  wire        _slots_22_io_uop_is_br;
  wire        _slots_22_io_uop_is_jalr;
  wire        _slots_22_io_uop_is_jal;
  wire        _slots_22_io_uop_is_sfb;
  wire [19:0] _slots_22_io_uop_br_mask;
  wire [4:0]  _slots_22_io_uop_br_tag;
  wire [5:0]  _slots_22_io_uop_ftq_idx;
  wire        _slots_22_io_uop_edge_inst;
  wire [5:0]  _slots_22_io_uop_pc_lob;
  wire        _slots_22_io_uop_taken;
  wire [19:0] _slots_22_io_uop_imm_packed;
  wire [11:0] _slots_22_io_uop_csr_addr;
  wire [6:0]  _slots_22_io_uop_rob_idx;
  wire [4:0]  _slots_22_io_uop_ldq_idx;
  wire [4:0]  _slots_22_io_uop_stq_idx;
  wire [1:0]  _slots_22_io_uop_rxq_idx;
  wire [6:0]  _slots_22_io_uop_pdst;
  wire [6:0]  _slots_22_io_uop_prs1;
  wire [6:0]  _slots_22_io_uop_prs2;
  wire [6:0]  _slots_22_io_uop_prs3;
  wire [5:0]  _slots_22_io_uop_ppred;
  wire        _slots_22_io_uop_prs1_busy;
  wire        _slots_22_io_uop_prs2_busy;
  wire        _slots_22_io_uop_prs3_busy;
  wire        _slots_22_io_uop_ppred_busy;
  wire [6:0]  _slots_22_io_uop_stale_pdst;
  wire        _slots_22_io_uop_exception;
  wire [63:0] _slots_22_io_uop_exc_cause;
  wire        _slots_22_io_uop_bypassable;
  wire [4:0]  _slots_22_io_uop_mem_cmd;
  wire [1:0]  _slots_22_io_uop_mem_size;
  wire        _slots_22_io_uop_mem_signed;
  wire        _slots_22_io_uop_is_fence;
  wire        _slots_22_io_uop_is_fencei;
  wire        _slots_22_io_uop_is_amo;
  wire        _slots_22_io_uop_uses_ldq;
  wire        _slots_22_io_uop_uses_stq;
  wire        _slots_22_io_uop_is_sys_pc2epc;
  wire        _slots_22_io_uop_is_unique;
  wire        _slots_22_io_uop_flush_on_commit;
  wire        _slots_22_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_22_io_uop_ldst;
  wire [5:0]  _slots_22_io_uop_lrs1;
  wire [5:0]  _slots_22_io_uop_lrs2;
  wire [5:0]  _slots_22_io_uop_lrs3;
  wire        _slots_22_io_uop_ldst_val;
  wire [1:0]  _slots_22_io_uop_dst_rtype;
  wire [1:0]  _slots_22_io_uop_lrs1_rtype;
  wire [1:0]  _slots_22_io_uop_lrs2_rtype;
  wire        _slots_22_io_uop_frs3_en;
  wire        _slots_22_io_uop_fp_val;
  wire        _slots_22_io_uop_fp_single;
  wire        _slots_22_io_uop_xcpt_pf_if;
  wire        _slots_22_io_uop_xcpt_ae_if;
  wire        _slots_22_io_uop_xcpt_ma_if;
  wire        _slots_22_io_uop_bp_debug_if;
  wire        _slots_22_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_22_io_uop_debug_fsrc;
  wire [1:0]  _slots_22_io_uop_debug_tsrc;
  wire        _slots_21_io_valid;
  wire        _slots_21_io_will_be_valid;
  wire        _slots_21_io_request;
  wire [6:0]  _slots_21_io_out_uop_uopc;
  wire [31:0] _slots_21_io_out_uop_inst;
  wire [31:0] _slots_21_io_out_uop_debug_inst;
  wire        _slots_21_io_out_uop_is_rvc;
  wire [39:0] _slots_21_io_out_uop_debug_pc;
  wire [2:0]  _slots_21_io_out_uop_iq_type;
  wire [9:0]  _slots_21_io_out_uop_fu_code;
  wire [1:0]  _slots_21_io_out_uop_iw_state;
  wire        _slots_21_io_out_uop_iw_p1_poisoned;
  wire        _slots_21_io_out_uop_iw_p2_poisoned;
  wire        _slots_21_io_out_uop_is_br;
  wire        _slots_21_io_out_uop_is_jalr;
  wire        _slots_21_io_out_uop_is_jal;
  wire        _slots_21_io_out_uop_is_sfb;
  wire [19:0] _slots_21_io_out_uop_br_mask;
  wire [4:0]  _slots_21_io_out_uop_br_tag;
  wire [5:0]  _slots_21_io_out_uop_ftq_idx;
  wire        _slots_21_io_out_uop_edge_inst;
  wire [5:0]  _slots_21_io_out_uop_pc_lob;
  wire        _slots_21_io_out_uop_taken;
  wire [19:0] _slots_21_io_out_uop_imm_packed;
  wire [11:0] _slots_21_io_out_uop_csr_addr;
  wire [6:0]  _slots_21_io_out_uop_rob_idx;
  wire [4:0]  _slots_21_io_out_uop_ldq_idx;
  wire [4:0]  _slots_21_io_out_uop_stq_idx;
  wire [1:0]  _slots_21_io_out_uop_rxq_idx;
  wire [6:0]  _slots_21_io_out_uop_pdst;
  wire [6:0]  _slots_21_io_out_uop_prs1;
  wire [6:0]  _slots_21_io_out_uop_prs2;
  wire [6:0]  _slots_21_io_out_uop_prs3;
  wire [5:0]  _slots_21_io_out_uop_ppred;
  wire        _slots_21_io_out_uop_prs1_busy;
  wire        _slots_21_io_out_uop_prs2_busy;
  wire        _slots_21_io_out_uop_prs3_busy;
  wire        _slots_21_io_out_uop_ppred_busy;
  wire [6:0]  _slots_21_io_out_uop_stale_pdst;
  wire        _slots_21_io_out_uop_exception;
  wire [63:0] _slots_21_io_out_uop_exc_cause;
  wire        _slots_21_io_out_uop_bypassable;
  wire [4:0]  _slots_21_io_out_uop_mem_cmd;
  wire [1:0]  _slots_21_io_out_uop_mem_size;
  wire        _slots_21_io_out_uop_mem_signed;
  wire        _slots_21_io_out_uop_is_fence;
  wire        _slots_21_io_out_uop_is_fencei;
  wire        _slots_21_io_out_uop_is_amo;
  wire        _slots_21_io_out_uop_uses_ldq;
  wire        _slots_21_io_out_uop_uses_stq;
  wire        _slots_21_io_out_uop_is_sys_pc2epc;
  wire        _slots_21_io_out_uop_is_unique;
  wire        _slots_21_io_out_uop_flush_on_commit;
  wire        _slots_21_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_21_io_out_uop_ldst;
  wire [5:0]  _slots_21_io_out_uop_lrs1;
  wire [5:0]  _slots_21_io_out_uop_lrs2;
  wire [5:0]  _slots_21_io_out_uop_lrs3;
  wire        _slots_21_io_out_uop_ldst_val;
  wire [1:0]  _slots_21_io_out_uop_dst_rtype;
  wire [1:0]  _slots_21_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_21_io_out_uop_lrs2_rtype;
  wire        _slots_21_io_out_uop_frs3_en;
  wire        _slots_21_io_out_uop_fp_val;
  wire        _slots_21_io_out_uop_fp_single;
  wire        _slots_21_io_out_uop_xcpt_pf_if;
  wire        _slots_21_io_out_uop_xcpt_ae_if;
  wire        _slots_21_io_out_uop_xcpt_ma_if;
  wire        _slots_21_io_out_uop_bp_debug_if;
  wire        _slots_21_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_21_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_21_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_21_io_uop_uopc;
  wire [31:0] _slots_21_io_uop_inst;
  wire [31:0] _slots_21_io_uop_debug_inst;
  wire        _slots_21_io_uop_is_rvc;
  wire [39:0] _slots_21_io_uop_debug_pc;
  wire [2:0]  _slots_21_io_uop_iq_type;
  wire [9:0]  _slots_21_io_uop_fu_code;
  wire [1:0]  _slots_21_io_uop_iw_state;
  wire        _slots_21_io_uop_iw_p1_poisoned;
  wire        _slots_21_io_uop_iw_p2_poisoned;
  wire        _slots_21_io_uop_is_br;
  wire        _slots_21_io_uop_is_jalr;
  wire        _slots_21_io_uop_is_jal;
  wire        _slots_21_io_uop_is_sfb;
  wire [19:0] _slots_21_io_uop_br_mask;
  wire [4:0]  _slots_21_io_uop_br_tag;
  wire [5:0]  _slots_21_io_uop_ftq_idx;
  wire        _slots_21_io_uop_edge_inst;
  wire [5:0]  _slots_21_io_uop_pc_lob;
  wire        _slots_21_io_uop_taken;
  wire [19:0] _slots_21_io_uop_imm_packed;
  wire [11:0] _slots_21_io_uop_csr_addr;
  wire [6:0]  _slots_21_io_uop_rob_idx;
  wire [4:0]  _slots_21_io_uop_ldq_idx;
  wire [4:0]  _slots_21_io_uop_stq_idx;
  wire [1:0]  _slots_21_io_uop_rxq_idx;
  wire [6:0]  _slots_21_io_uop_pdst;
  wire [6:0]  _slots_21_io_uop_prs1;
  wire [6:0]  _slots_21_io_uop_prs2;
  wire [6:0]  _slots_21_io_uop_prs3;
  wire [5:0]  _slots_21_io_uop_ppred;
  wire        _slots_21_io_uop_prs1_busy;
  wire        _slots_21_io_uop_prs2_busy;
  wire        _slots_21_io_uop_prs3_busy;
  wire        _slots_21_io_uop_ppred_busy;
  wire [6:0]  _slots_21_io_uop_stale_pdst;
  wire        _slots_21_io_uop_exception;
  wire [63:0] _slots_21_io_uop_exc_cause;
  wire        _slots_21_io_uop_bypassable;
  wire [4:0]  _slots_21_io_uop_mem_cmd;
  wire [1:0]  _slots_21_io_uop_mem_size;
  wire        _slots_21_io_uop_mem_signed;
  wire        _slots_21_io_uop_is_fence;
  wire        _slots_21_io_uop_is_fencei;
  wire        _slots_21_io_uop_is_amo;
  wire        _slots_21_io_uop_uses_ldq;
  wire        _slots_21_io_uop_uses_stq;
  wire        _slots_21_io_uop_is_sys_pc2epc;
  wire        _slots_21_io_uop_is_unique;
  wire        _slots_21_io_uop_flush_on_commit;
  wire        _slots_21_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_21_io_uop_ldst;
  wire [5:0]  _slots_21_io_uop_lrs1;
  wire [5:0]  _slots_21_io_uop_lrs2;
  wire [5:0]  _slots_21_io_uop_lrs3;
  wire        _slots_21_io_uop_ldst_val;
  wire [1:0]  _slots_21_io_uop_dst_rtype;
  wire [1:0]  _slots_21_io_uop_lrs1_rtype;
  wire [1:0]  _slots_21_io_uop_lrs2_rtype;
  wire        _slots_21_io_uop_frs3_en;
  wire        _slots_21_io_uop_fp_val;
  wire        _slots_21_io_uop_fp_single;
  wire        _slots_21_io_uop_xcpt_pf_if;
  wire        _slots_21_io_uop_xcpt_ae_if;
  wire        _slots_21_io_uop_xcpt_ma_if;
  wire        _slots_21_io_uop_bp_debug_if;
  wire        _slots_21_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_21_io_uop_debug_fsrc;
  wire [1:0]  _slots_21_io_uop_debug_tsrc;
  wire        _slots_20_io_valid;
  wire        _slots_20_io_will_be_valid;
  wire        _slots_20_io_request;
  wire [6:0]  _slots_20_io_out_uop_uopc;
  wire [31:0] _slots_20_io_out_uop_inst;
  wire [31:0] _slots_20_io_out_uop_debug_inst;
  wire        _slots_20_io_out_uop_is_rvc;
  wire [39:0] _slots_20_io_out_uop_debug_pc;
  wire [2:0]  _slots_20_io_out_uop_iq_type;
  wire [9:0]  _slots_20_io_out_uop_fu_code;
  wire [1:0]  _slots_20_io_out_uop_iw_state;
  wire        _slots_20_io_out_uop_iw_p1_poisoned;
  wire        _slots_20_io_out_uop_iw_p2_poisoned;
  wire        _slots_20_io_out_uop_is_br;
  wire        _slots_20_io_out_uop_is_jalr;
  wire        _slots_20_io_out_uop_is_jal;
  wire        _slots_20_io_out_uop_is_sfb;
  wire [19:0] _slots_20_io_out_uop_br_mask;
  wire [4:0]  _slots_20_io_out_uop_br_tag;
  wire [5:0]  _slots_20_io_out_uop_ftq_idx;
  wire        _slots_20_io_out_uop_edge_inst;
  wire [5:0]  _slots_20_io_out_uop_pc_lob;
  wire        _slots_20_io_out_uop_taken;
  wire [19:0] _slots_20_io_out_uop_imm_packed;
  wire [11:0] _slots_20_io_out_uop_csr_addr;
  wire [6:0]  _slots_20_io_out_uop_rob_idx;
  wire [4:0]  _slots_20_io_out_uop_ldq_idx;
  wire [4:0]  _slots_20_io_out_uop_stq_idx;
  wire [1:0]  _slots_20_io_out_uop_rxq_idx;
  wire [6:0]  _slots_20_io_out_uop_pdst;
  wire [6:0]  _slots_20_io_out_uop_prs1;
  wire [6:0]  _slots_20_io_out_uop_prs2;
  wire [6:0]  _slots_20_io_out_uop_prs3;
  wire [5:0]  _slots_20_io_out_uop_ppred;
  wire        _slots_20_io_out_uop_prs1_busy;
  wire        _slots_20_io_out_uop_prs2_busy;
  wire        _slots_20_io_out_uop_prs3_busy;
  wire        _slots_20_io_out_uop_ppred_busy;
  wire [6:0]  _slots_20_io_out_uop_stale_pdst;
  wire        _slots_20_io_out_uop_exception;
  wire [63:0] _slots_20_io_out_uop_exc_cause;
  wire        _slots_20_io_out_uop_bypassable;
  wire [4:0]  _slots_20_io_out_uop_mem_cmd;
  wire [1:0]  _slots_20_io_out_uop_mem_size;
  wire        _slots_20_io_out_uop_mem_signed;
  wire        _slots_20_io_out_uop_is_fence;
  wire        _slots_20_io_out_uop_is_fencei;
  wire        _slots_20_io_out_uop_is_amo;
  wire        _slots_20_io_out_uop_uses_ldq;
  wire        _slots_20_io_out_uop_uses_stq;
  wire        _slots_20_io_out_uop_is_sys_pc2epc;
  wire        _slots_20_io_out_uop_is_unique;
  wire        _slots_20_io_out_uop_flush_on_commit;
  wire        _slots_20_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_20_io_out_uop_ldst;
  wire [5:0]  _slots_20_io_out_uop_lrs1;
  wire [5:0]  _slots_20_io_out_uop_lrs2;
  wire [5:0]  _slots_20_io_out_uop_lrs3;
  wire        _slots_20_io_out_uop_ldst_val;
  wire [1:0]  _slots_20_io_out_uop_dst_rtype;
  wire [1:0]  _slots_20_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_20_io_out_uop_lrs2_rtype;
  wire        _slots_20_io_out_uop_frs3_en;
  wire        _slots_20_io_out_uop_fp_val;
  wire        _slots_20_io_out_uop_fp_single;
  wire        _slots_20_io_out_uop_xcpt_pf_if;
  wire        _slots_20_io_out_uop_xcpt_ae_if;
  wire        _slots_20_io_out_uop_xcpt_ma_if;
  wire        _slots_20_io_out_uop_bp_debug_if;
  wire        _slots_20_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_20_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_20_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_20_io_uop_uopc;
  wire [31:0] _slots_20_io_uop_inst;
  wire [31:0] _slots_20_io_uop_debug_inst;
  wire        _slots_20_io_uop_is_rvc;
  wire [39:0] _slots_20_io_uop_debug_pc;
  wire [2:0]  _slots_20_io_uop_iq_type;
  wire [9:0]  _slots_20_io_uop_fu_code;
  wire [1:0]  _slots_20_io_uop_iw_state;
  wire        _slots_20_io_uop_iw_p1_poisoned;
  wire        _slots_20_io_uop_iw_p2_poisoned;
  wire        _slots_20_io_uop_is_br;
  wire        _slots_20_io_uop_is_jalr;
  wire        _slots_20_io_uop_is_jal;
  wire        _slots_20_io_uop_is_sfb;
  wire [19:0] _slots_20_io_uop_br_mask;
  wire [4:0]  _slots_20_io_uop_br_tag;
  wire [5:0]  _slots_20_io_uop_ftq_idx;
  wire        _slots_20_io_uop_edge_inst;
  wire [5:0]  _slots_20_io_uop_pc_lob;
  wire        _slots_20_io_uop_taken;
  wire [19:0] _slots_20_io_uop_imm_packed;
  wire [11:0] _slots_20_io_uop_csr_addr;
  wire [6:0]  _slots_20_io_uop_rob_idx;
  wire [4:0]  _slots_20_io_uop_ldq_idx;
  wire [4:0]  _slots_20_io_uop_stq_idx;
  wire [1:0]  _slots_20_io_uop_rxq_idx;
  wire [6:0]  _slots_20_io_uop_pdst;
  wire [6:0]  _slots_20_io_uop_prs1;
  wire [6:0]  _slots_20_io_uop_prs2;
  wire [6:0]  _slots_20_io_uop_prs3;
  wire [5:0]  _slots_20_io_uop_ppred;
  wire        _slots_20_io_uop_prs1_busy;
  wire        _slots_20_io_uop_prs2_busy;
  wire        _slots_20_io_uop_prs3_busy;
  wire        _slots_20_io_uop_ppred_busy;
  wire [6:0]  _slots_20_io_uop_stale_pdst;
  wire        _slots_20_io_uop_exception;
  wire [63:0] _slots_20_io_uop_exc_cause;
  wire        _slots_20_io_uop_bypassable;
  wire [4:0]  _slots_20_io_uop_mem_cmd;
  wire [1:0]  _slots_20_io_uop_mem_size;
  wire        _slots_20_io_uop_mem_signed;
  wire        _slots_20_io_uop_is_fence;
  wire        _slots_20_io_uop_is_fencei;
  wire        _slots_20_io_uop_is_amo;
  wire        _slots_20_io_uop_uses_ldq;
  wire        _slots_20_io_uop_uses_stq;
  wire        _slots_20_io_uop_is_sys_pc2epc;
  wire        _slots_20_io_uop_is_unique;
  wire        _slots_20_io_uop_flush_on_commit;
  wire        _slots_20_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_20_io_uop_ldst;
  wire [5:0]  _slots_20_io_uop_lrs1;
  wire [5:0]  _slots_20_io_uop_lrs2;
  wire [5:0]  _slots_20_io_uop_lrs3;
  wire        _slots_20_io_uop_ldst_val;
  wire [1:0]  _slots_20_io_uop_dst_rtype;
  wire [1:0]  _slots_20_io_uop_lrs1_rtype;
  wire [1:0]  _slots_20_io_uop_lrs2_rtype;
  wire        _slots_20_io_uop_frs3_en;
  wire        _slots_20_io_uop_fp_val;
  wire        _slots_20_io_uop_fp_single;
  wire        _slots_20_io_uop_xcpt_pf_if;
  wire        _slots_20_io_uop_xcpt_ae_if;
  wire        _slots_20_io_uop_xcpt_ma_if;
  wire        _slots_20_io_uop_bp_debug_if;
  wire        _slots_20_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_20_io_uop_debug_fsrc;
  wire [1:0]  _slots_20_io_uop_debug_tsrc;
  wire        _slots_19_io_valid;
  wire        _slots_19_io_will_be_valid;
  wire        _slots_19_io_request;
  wire [6:0]  _slots_19_io_out_uop_uopc;
  wire [31:0] _slots_19_io_out_uop_inst;
  wire [31:0] _slots_19_io_out_uop_debug_inst;
  wire        _slots_19_io_out_uop_is_rvc;
  wire [39:0] _slots_19_io_out_uop_debug_pc;
  wire [2:0]  _slots_19_io_out_uop_iq_type;
  wire [9:0]  _slots_19_io_out_uop_fu_code;
  wire [1:0]  _slots_19_io_out_uop_iw_state;
  wire        _slots_19_io_out_uop_iw_p1_poisoned;
  wire        _slots_19_io_out_uop_iw_p2_poisoned;
  wire        _slots_19_io_out_uop_is_br;
  wire        _slots_19_io_out_uop_is_jalr;
  wire        _slots_19_io_out_uop_is_jal;
  wire        _slots_19_io_out_uop_is_sfb;
  wire [19:0] _slots_19_io_out_uop_br_mask;
  wire [4:0]  _slots_19_io_out_uop_br_tag;
  wire [5:0]  _slots_19_io_out_uop_ftq_idx;
  wire        _slots_19_io_out_uop_edge_inst;
  wire [5:0]  _slots_19_io_out_uop_pc_lob;
  wire        _slots_19_io_out_uop_taken;
  wire [19:0] _slots_19_io_out_uop_imm_packed;
  wire [11:0] _slots_19_io_out_uop_csr_addr;
  wire [6:0]  _slots_19_io_out_uop_rob_idx;
  wire [4:0]  _slots_19_io_out_uop_ldq_idx;
  wire [4:0]  _slots_19_io_out_uop_stq_idx;
  wire [1:0]  _slots_19_io_out_uop_rxq_idx;
  wire [6:0]  _slots_19_io_out_uop_pdst;
  wire [6:0]  _slots_19_io_out_uop_prs1;
  wire [6:0]  _slots_19_io_out_uop_prs2;
  wire [6:0]  _slots_19_io_out_uop_prs3;
  wire [5:0]  _slots_19_io_out_uop_ppred;
  wire        _slots_19_io_out_uop_prs1_busy;
  wire        _slots_19_io_out_uop_prs2_busy;
  wire        _slots_19_io_out_uop_prs3_busy;
  wire        _slots_19_io_out_uop_ppred_busy;
  wire [6:0]  _slots_19_io_out_uop_stale_pdst;
  wire        _slots_19_io_out_uop_exception;
  wire [63:0] _slots_19_io_out_uop_exc_cause;
  wire        _slots_19_io_out_uop_bypassable;
  wire [4:0]  _slots_19_io_out_uop_mem_cmd;
  wire [1:0]  _slots_19_io_out_uop_mem_size;
  wire        _slots_19_io_out_uop_mem_signed;
  wire        _slots_19_io_out_uop_is_fence;
  wire        _slots_19_io_out_uop_is_fencei;
  wire        _slots_19_io_out_uop_is_amo;
  wire        _slots_19_io_out_uop_uses_ldq;
  wire        _slots_19_io_out_uop_uses_stq;
  wire        _slots_19_io_out_uop_is_sys_pc2epc;
  wire        _slots_19_io_out_uop_is_unique;
  wire        _slots_19_io_out_uop_flush_on_commit;
  wire        _slots_19_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_19_io_out_uop_ldst;
  wire [5:0]  _slots_19_io_out_uop_lrs1;
  wire [5:0]  _slots_19_io_out_uop_lrs2;
  wire [5:0]  _slots_19_io_out_uop_lrs3;
  wire        _slots_19_io_out_uop_ldst_val;
  wire [1:0]  _slots_19_io_out_uop_dst_rtype;
  wire [1:0]  _slots_19_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_19_io_out_uop_lrs2_rtype;
  wire        _slots_19_io_out_uop_frs3_en;
  wire        _slots_19_io_out_uop_fp_val;
  wire        _slots_19_io_out_uop_fp_single;
  wire        _slots_19_io_out_uop_xcpt_pf_if;
  wire        _slots_19_io_out_uop_xcpt_ae_if;
  wire        _slots_19_io_out_uop_xcpt_ma_if;
  wire        _slots_19_io_out_uop_bp_debug_if;
  wire        _slots_19_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_19_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_19_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_19_io_uop_uopc;
  wire [31:0] _slots_19_io_uop_inst;
  wire [31:0] _slots_19_io_uop_debug_inst;
  wire        _slots_19_io_uop_is_rvc;
  wire [39:0] _slots_19_io_uop_debug_pc;
  wire [2:0]  _slots_19_io_uop_iq_type;
  wire [9:0]  _slots_19_io_uop_fu_code;
  wire [1:0]  _slots_19_io_uop_iw_state;
  wire        _slots_19_io_uop_iw_p1_poisoned;
  wire        _slots_19_io_uop_iw_p2_poisoned;
  wire        _slots_19_io_uop_is_br;
  wire        _slots_19_io_uop_is_jalr;
  wire        _slots_19_io_uop_is_jal;
  wire        _slots_19_io_uop_is_sfb;
  wire [19:0] _slots_19_io_uop_br_mask;
  wire [4:0]  _slots_19_io_uop_br_tag;
  wire [5:0]  _slots_19_io_uop_ftq_idx;
  wire        _slots_19_io_uop_edge_inst;
  wire [5:0]  _slots_19_io_uop_pc_lob;
  wire        _slots_19_io_uop_taken;
  wire [19:0] _slots_19_io_uop_imm_packed;
  wire [11:0] _slots_19_io_uop_csr_addr;
  wire [6:0]  _slots_19_io_uop_rob_idx;
  wire [4:0]  _slots_19_io_uop_ldq_idx;
  wire [4:0]  _slots_19_io_uop_stq_idx;
  wire [1:0]  _slots_19_io_uop_rxq_idx;
  wire [6:0]  _slots_19_io_uop_pdst;
  wire [6:0]  _slots_19_io_uop_prs1;
  wire [6:0]  _slots_19_io_uop_prs2;
  wire [6:0]  _slots_19_io_uop_prs3;
  wire [5:0]  _slots_19_io_uop_ppred;
  wire        _slots_19_io_uop_prs1_busy;
  wire        _slots_19_io_uop_prs2_busy;
  wire        _slots_19_io_uop_prs3_busy;
  wire        _slots_19_io_uop_ppred_busy;
  wire [6:0]  _slots_19_io_uop_stale_pdst;
  wire        _slots_19_io_uop_exception;
  wire [63:0] _slots_19_io_uop_exc_cause;
  wire        _slots_19_io_uop_bypassable;
  wire [4:0]  _slots_19_io_uop_mem_cmd;
  wire [1:0]  _slots_19_io_uop_mem_size;
  wire        _slots_19_io_uop_mem_signed;
  wire        _slots_19_io_uop_is_fence;
  wire        _slots_19_io_uop_is_fencei;
  wire        _slots_19_io_uop_is_amo;
  wire        _slots_19_io_uop_uses_ldq;
  wire        _slots_19_io_uop_uses_stq;
  wire        _slots_19_io_uop_is_sys_pc2epc;
  wire        _slots_19_io_uop_is_unique;
  wire        _slots_19_io_uop_flush_on_commit;
  wire        _slots_19_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_19_io_uop_ldst;
  wire [5:0]  _slots_19_io_uop_lrs1;
  wire [5:0]  _slots_19_io_uop_lrs2;
  wire [5:0]  _slots_19_io_uop_lrs3;
  wire        _slots_19_io_uop_ldst_val;
  wire [1:0]  _slots_19_io_uop_dst_rtype;
  wire [1:0]  _slots_19_io_uop_lrs1_rtype;
  wire [1:0]  _slots_19_io_uop_lrs2_rtype;
  wire        _slots_19_io_uop_frs3_en;
  wire        _slots_19_io_uop_fp_val;
  wire        _slots_19_io_uop_fp_single;
  wire        _slots_19_io_uop_xcpt_pf_if;
  wire        _slots_19_io_uop_xcpt_ae_if;
  wire        _slots_19_io_uop_xcpt_ma_if;
  wire        _slots_19_io_uop_bp_debug_if;
  wire        _slots_19_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_19_io_uop_debug_fsrc;
  wire [1:0]  _slots_19_io_uop_debug_tsrc;
  wire        _slots_18_io_valid;
  wire        _slots_18_io_will_be_valid;
  wire        _slots_18_io_request;
  wire [6:0]  _slots_18_io_out_uop_uopc;
  wire [31:0] _slots_18_io_out_uop_inst;
  wire [31:0] _slots_18_io_out_uop_debug_inst;
  wire        _slots_18_io_out_uop_is_rvc;
  wire [39:0] _slots_18_io_out_uop_debug_pc;
  wire [2:0]  _slots_18_io_out_uop_iq_type;
  wire [9:0]  _slots_18_io_out_uop_fu_code;
  wire [1:0]  _slots_18_io_out_uop_iw_state;
  wire        _slots_18_io_out_uop_iw_p1_poisoned;
  wire        _slots_18_io_out_uop_iw_p2_poisoned;
  wire        _slots_18_io_out_uop_is_br;
  wire        _slots_18_io_out_uop_is_jalr;
  wire        _slots_18_io_out_uop_is_jal;
  wire        _slots_18_io_out_uop_is_sfb;
  wire [19:0] _slots_18_io_out_uop_br_mask;
  wire [4:0]  _slots_18_io_out_uop_br_tag;
  wire [5:0]  _slots_18_io_out_uop_ftq_idx;
  wire        _slots_18_io_out_uop_edge_inst;
  wire [5:0]  _slots_18_io_out_uop_pc_lob;
  wire        _slots_18_io_out_uop_taken;
  wire [19:0] _slots_18_io_out_uop_imm_packed;
  wire [11:0] _slots_18_io_out_uop_csr_addr;
  wire [6:0]  _slots_18_io_out_uop_rob_idx;
  wire [4:0]  _slots_18_io_out_uop_ldq_idx;
  wire [4:0]  _slots_18_io_out_uop_stq_idx;
  wire [1:0]  _slots_18_io_out_uop_rxq_idx;
  wire [6:0]  _slots_18_io_out_uop_pdst;
  wire [6:0]  _slots_18_io_out_uop_prs1;
  wire [6:0]  _slots_18_io_out_uop_prs2;
  wire [6:0]  _slots_18_io_out_uop_prs3;
  wire [5:0]  _slots_18_io_out_uop_ppred;
  wire        _slots_18_io_out_uop_prs1_busy;
  wire        _slots_18_io_out_uop_prs2_busy;
  wire        _slots_18_io_out_uop_prs3_busy;
  wire        _slots_18_io_out_uop_ppred_busy;
  wire [6:0]  _slots_18_io_out_uop_stale_pdst;
  wire        _slots_18_io_out_uop_exception;
  wire [63:0] _slots_18_io_out_uop_exc_cause;
  wire        _slots_18_io_out_uop_bypassable;
  wire [4:0]  _slots_18_io_out_uop_mem_cmd;
  wire [1:0]  _slots_18_io_out_uop_mem_size;
  wire        _slots_18_io_out_uop_mem_signed;
  wire        _slots_18_io_out_uop_is_fence;
  wire        _slots_18_io_out_uop_is_fencei;
  wire        _slots_18_io_out_uop_is_amo;
  wire        _slots_18_io_out_uop_uses_ldq;
  wire        _slots_18_io_out_uop_uses_stq;
  wire        _slots_18_io_out_uop_is_sys_pc2epc;
  wire        _slots_18_io_out_uop_is_unique;
  wire        _slots_18_io_out_uop_flush_on_commit;
  wire        _slots_18_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_18_io_out_uop_ldst;
  wire [5:0]  _slots_18_io_out_uop_lrs1;
  wire [5:0]  _slots_18_io_out_uop_lrs2;
  wire [5:0]  _slots_18_io_out_uop_lrs3;
  wire        _slots_18_io_out_uop_ldst_val;
  wire [1:0]  _slots_18_io_out_uop_dst_rtype;
  wire [1:0]  _slots_18_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_18_io_out_uop_lrs2_rtype;
  wire        _slots_18_io_out_uop_frs3_en;
  wire        _slots_18_io_out_uop_fp_val;
  wire        _slots_18_io_out_uop_fp_single;
  wire        _slots_18_io_out_uop_xcpt_pf_if;
  wire        _slots_18_io_out_uop_xcpt_ae_if;
  wire        _slots_18_io_out_uop_xcpt_ma_if;
  wire        _slots_18_io_out_uop_bp_debug_if;
  wire        _slots_18_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_18_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_18_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_18_io_uop_uopc;
  wire [31:0] _slots_18_io_uop_inst;
  wire [31:0] _slots_18_io_uop_debug_inst;
  wire        _slots_18_io_uop_is_rvc;
  wire [39:0] _slots_18_io_uop_debug_pc;
  wire [2:0]  _slots_18_io_uop_iq_type;
  wire [9:0]  _slots_18_io_uop_fu_code;
  wire [1:0]  _slots_18_io_uop_iw_state;
  wire        _slots_18_io_uop_iw_p1_poisoned;
  wire        _slots_18_io_uop_iw_p2_poisoned;
  wire        _slots_18_io_uop_is_br;
  wire        _slots_18_io_uop_is_jalr;
  wire        _slots_18_io_uop_is_jal;
  wire        _slots_18_io_uop_is_sfb;
  wire [19:0] _slots_18_io_uop_br_mask;
  wire [4:0]  _slots_18_io_uop_br_tag;
  wire [5:0]  _slots_18_io_uop_ftq_idx;
  wire        _slots_18_io_uop_edge_inst;
  wire [5:0]  _slots_18_io_uop_pc_lob;
  wire        _slots_18_io_uop_taken;
  wire [19:0] _slots_18_io_uop_imm_packed;
  wire [11:0] _slots_18_io_uop_csr_addr;
  wire [6:0]  _slots_18_io_uop_rob_idx;
  wire [4:0]  _slots_18_io_uop_ldq_idx;
  wire [4:0]  _slots_18_io_uop_stq_idx;
  wire [1:0]  _slots_18_io_uop_rxq_idx;
  wire [6:0]  _slots_18_io_uop_pdst;
  wire [6:0]  _slots_18_io_uop_prs1;
  wire [6:0]  _slots_18_io_uop_prs2;
  wire [6:0]  _slots_18_io_uop_prs3;
  wire [5:0]  _slots_18_io_uop_ppred;
  wire        _slots_18_io_uop_prs1_busy;
  wire        _slots_18_io_uop_prs2_busy;
  wire        _slots_18_io_uop_prs3_busy;
  wire        _slots_18_io_uop_ppred_busy;
  wire [6:0]  _slots_18_io_uop_stale_pdst;
  wire        _slots_18_io_uop_exception;
  wire [63:0] _slots_18_io_uop_exc_cause;
  wire        _slots_18_io_uop_bypassable;
  wire [4:0]  _slots_18_io_uop_mem_cmd;
  wire [1:0]  _slots_18_io_uop_mem_size;
  wire        _slots_18_io_uop_mem_signed;
  wire        _slots_18_io_uop_is_fence;
  wire        _slots_18_io_uop_is_fencei;
  wire        _slots_18_io_uop_is_amo;
  wire        _slots_18_io_uop_uses_ldq;
  wire        _slots_18_io_uop_uses_stq;
  wire        _slots_18_io_uop_is_sys_pc2epc;
  wire        _slots_18_io_uop_is_unique;
  wire        _slots_18_io_uop_flush_on_commit;
  wire        _slots_18_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_18_io_uop_ldst;
  wire [5:0]  _slots_18_io_uop_lrs1;
  wire [5:0]  _slots_18_io_uop_lrs2;
  wire [5:0]  _slots_18_io_uop_lrs3;
  wire        _slots_18_io_uop_ldst_val;
  wire [1:0]  _slots_18_io_uop_dst_rtype;
  wire [1:0]  _slots_18_io_uop_lrs1_rtype;
  wire [1:0]  _slots_18_io_uop_lrs2_rtype;
  wire        _slots_18_io_uop_frs3_en;
  wire        _slots_18_io_uop_fp_val;
  wire        _slots_18_io_uop_fp_single;
  wire        _slots_18_io_uop_xcpt_pf_if;
  wire        _slots_18_io_uop_xcpt_ae_if;
  wire        _slots_18_io_uop_xcpt_ma_if;
  wire        _slots_18_io_uop_bp_debug_if;
  wire        _slots_18_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_18_io_uop_debug_fsrc;
  wire [1:0]  _slots_18_io_uop_debug_tsrc;
  wire        _slots_17_io_valid;
  wire        _slots_17_io_will_be_valid;
  wire        _slots_17_io_request;
  wire [6:0]  _slots_17_io_out_uop_uopc;
  wire [31:0] _slots_17_io_out_uop_inst;
  wire [31:0] _slots_17_io_out_uop_debug_inst;
  wire        _slots_17_io_out_uop_is_rvc;
  wire [39:0] _slots_17_io_out_uop_debug_pc;
  wire [2:0]  _slots_17_io_out_uop_iq_type;
  wire [9:0]  _slots_17_io_out_uop_fu_code;
  wire [1:0]  _slots_17_io_out_uop_iw_state;
  wire        _slots_17_io_out_uop_iw_p1_poisoned;
  wire        _slots_17_io_out_uop_iw_p2_poisoned;
  wire        _slots_17_io_out_uop_is_br;
  wire        _slots_17_io_out_uop_is_jalr;
  wire        _slots_17_io_out_uop_is_jal;
  wire        _slots_17_io_out_uop_is_sfb;
  wire [19:0] _slots_17_io_out_uop_br_mask;
  wire [4:0]  _slots_17_io_out_uop_br_tag;
  wire [5:0]  _slots_17_io_out_uop_ftq_idx;
  wire        _slots_17_io_out_uop_edge_inst;
  wire [5:0]  _slots_17_io_out_uop_pc_lob;
  wire        _slots_17_io_out_uop_taken;
  wire [19:0] _slots_17_io_out_uop_imm_packed;
  wire [11:0] _slots_17_io_out_uop_csr_addr;
  wire [6:0]  _slots_17_io_out_uop_rob_idx;
  wire [4:0]  _slots_17_io_out_uop_ldq_idx;
  wire [4:0]  _slots_17_io_out_uop_stq_idx;
  wire [1:0]  _slots_17_io_out_uop_rxq_idx;
  wire [6:0]  _slots_17_io_out_uop_pdst;
  wire [6:0]  _slots_17_io_out_uop_prs1;
  wire [6:0]  _slots_17_io_out_uop_prs2;
  wire [6:0]  _slots_17_io_out_uop_prs3;
  wire [5:0]  _slots_17_io_out_uop_ppred;
  wire        _slots_17_io_out_uop_prs1_busy;
  wire        _slots_17_io_out_uop_prs2_busy;
  wire        _slots_17_io_out_uop_prs3_busy;
  wire        _slots_17_io_out_uop_ppred_busy;
  wire [6:0]  _slots_17_io_out_uop_stale_pdst;
  wire        _slots_17_io_out_uop_exception;
  wire [63:0] _slots_17_io_out_uop_exc_cause;
  wire        _slots_17_io_out_uop_bypassable;
  wire [4:0]  _slots_17_io_out_uop_mem_cmd;
  wire [1:0]  _slots_17_io_out_uop_mem_size;
  wire        _slots_17_io_out_uop_mem_signed;
  wire        _slots_17_io_out_uop_is_fence;
  wire        _slots_17_io_out_uop_is_fencei;
  wire        _slots_17_io_out_uop_is_amo;
  wire        _slots_17_io_out_uop_uses_ldq;
  wire        _slots_17_io_out_uop_uses_stq;
  wire        _slots_17_io_out_uop_is_sys_pc2epc;
  wire        _slots_17_io_out_uop_is_unique;
  wire        _slots_17_io_out_uop_flush_on_commit;
  wire        _slots_17_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_17_io_out_uop_ldst;
  wire [5:0]  _slots_17_io_out_uop_lrs1;
  wire [5:0]  _slots_17_io_out_uop_lrs2;
  wire [5:0]  _slots_17_io_out_uop_lrs3;
  wire        _slots_17_io_out_uop_ldst_val;
  wire [1:0]  _slots_17_io_out_uop_dst_rtype;
  wire [1:0]  _slots_17_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_17_io_out_uop_lrs2_rtype;
  wire        _slots_17_io_out_uop_frs3_en;
  wire        _slots_17_io_out_uop_fp_val;
  wire        _slots_17_io_out_uop_fp_single;
  wire        _slots_17_io_out_uop_xcpt_pf_if;
  wire        _slots_17_io_out_uop_xcpt_ae_if;
  wire        _slots_17_io_out_uop_xcpt_ma_if;
  wire        _slots_17_io_out_uop_bp_debug_if;
  wire        _slots_17_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_17_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_17_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_17_io_uop_uopc;
  wire [31:0] _slots_17_io_uop_inst;
  wire [31:0] _slots_17_io_uop_debug_inst;
  wire        _slots_17_io_uop_is_rvc;
  wire [39:0] _slots_17_io_uop_debug_pc;
  wire [2:0]  _slots_17_io_uop_iq_type;
  wire [9:0]  _slots_17_io_uop_fu_code;
  wire [1:0]  _slots_17_io_uop_iw_state;
  wire        _slots_17_io_uop_iw_p1_poisoned;
  wire        _slots_17_io_uop_iw_p2_poisoned;
  wire        _slots_17_io_uop_is_br;
  wire        _slots_17_io_uop_is_jalr;
  wire        _slots_17_io_uop_is_jal;
  wire        _slots_17_io_uop_is_sfb;
  wire [19:0] _slots_17_io_uop_br_mask;
  wire [4:0]  _slots_17_io_uop_br_tag;
  wire [5:0]  _slots_17_io_uop_ftq_idx;
  wire        _slots_17_io_uop_edge_inst;
  wire [5:0]  _slots_17_io_uop_pc_lob;
  wire        _slots_17_io_uop_taken;
  wire [19:0] _slots_17_io_uop_imm_packed;
  wire [11:0] _slots_17_io_uop_csr_addr;
  wire [6:0]  _slots_17_io_uop_rob_idx;
  wire [4:0]  _slots_17_io_uop_ldq_idx;
  wire [4:0]  _slots_17_io_uop_stq_idx;
  wire [1:0]  _slots_17_io_uop_rxq_idx;
  wire [6:0]  _slots_17_io_uop_pdst;
  wire [6:0]  _slots_17_io_uop_prs1;
  wire [6:0]  _slots_17_io_uop_prs2;
  wire [6:0]  _slots_17_io_uop_prs3;
  wire [5:0]  _slots_17_io_uop_ppred;
  wire        _slots_17_io_uop_prs1_busy;
  wire        _slots_17_io_uop_prs2_busy;
  wire        _slots_17_io_uop_prs3_busy;
  wire        _slots_17_io_uop_ppred_busy;
  wire [6:0]  _slots_17_io_uop_stale_pdst;
  wire        _slots_17_io_uop_exception;
  wire [63:0] _slots_17_io_uop_exc_cause;
  wire        _slots_17_io_uop_bypassable;
  wire [4:0]  _slots_17_io_uop_mem_cmd;
  wire [1:0]  _slots_17_io_uop_mem_size;
  wire        _slots_17_io_uop_mem_signed;
  wire        _slots_17_io_uop_is_fence;
  wire        _slots_17_io_uop_is_fencei;
  wire        _slots_17_io_uop_is_amo;
  wire        _slots_17_io_uop_uses_ldq;
  wire        _slots_17_io_uop_uses_stq;
  wire        _slots_17_io_uop_is_sys_pc2epc;
  wire        _slots_17_io_uop_is_unique;
  wire        _slots_17_io_uop_flush_on_commit;
  wire        _slots_17_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_17_io_uop_ldst;
  wire [5:0]  _slots_17_io_uop_lrs1;
  wire [5:0]  _slots_17_io_uop_lrs2;
  wire [5:0]  _slots_17_io_uop_lrs3;
  wire        _slots_17_io_uop_ldst_val;
  wire [1:0]  _slots_17_io_uop_dst_rtype;
  wire [1:0]  _slots_17_io_uop_lrs1_rtype;
  wire [1:0]  _slots_17_io_uop_lrs2_rtype;
  wire        _slots_17_io_uop_frs3_en;
  wire        _slots_17_io_uop_fp_val;
  wire        _slots_17_io_uop_fp_single;
  wire        _slots_17_io_uop_xcpt_pf_if;
  wire        _slots_17_io_uop_xcpt_ae_if;
  wire        _slots_17_io_uop_xcpt_ma_if;
  wire        _slots_17_io_uop_bp_debug_if;
  wire        _slots_17_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_17_io_uop_debug_fsrc;
  wire [1:0]  _slots_17_io_uop_debug_tsrc;
  wire        _slots_16_io_valid;
  wire        _slots_16_io_will_be_valid;
  wire        _slots_16_io_request;
  wire [6:0]  _slots_16_io_out_uop_uopc;
  wire [31:0] _slots_16_io_out_uop_inst;
  wire [31:0] _slots_16_io_out_uop_debug_inst;
  wire        _slots_16_io_out_uop_is_rvc;
  wire [39:0] _slots_16_io_out_uop_debug_pc;
  wire [2:0]  _slots_16_io_out_uop_iq_type;
  wire [9:0]  _slots_16_io_out_uop_fu_code;
  wire [1:0]  _slots_16_io_out_uop_iw_state;
  wire        _slots_16_io_out_uop_iw_p1_poisoned;
  wire        _slots_16_io_out_uop_iw_p2_poisoned;
  wire        _slots_16_io_out_uop_is_br;
  wire        _slots_16_io_out_uop_is_jalr;
  wire        _slots_16_io_out_uop_is_jal;
  wire        _slots_16_io_out_uop_is_sfb;
  wire [19:0] _slots_16_io_out_uop_br_mask;
  wire [4:0]  _slots_16_io_out_uop_br_tag;
  wire [5:0]  _slots_16_io_out_uop_ftq_idx;
  wire        _slots_16_io_out_uop_edge_inst;
  wire [5:0]  _slots_16_io_out_uop_pc_lob;
  wire        _slots_16_io_out_uop_taken;
  wire [19:0] _slots_16_io_out_uop_imm_packed;
  wire [11:0] _slots_16_io_out_uop_csr_addr;
  wire [6:0]  _slots_16_io_out_uop_rob_idx;
  wire [4:0]  _slots_16_io_out_uop_ldq_idx;
  wire [4:0]  _slots_16_io_out_uop_stq_idx;
  wire [1:0]  _slots_16_io_out_uop_rxq_idx;
  wire [6:0]  _slots_16_io_out_uop_pdst;
  wire [6:0]  _slots_16_io_out_uop_prs1;
  wire [6:0]  _slots_16_io_out_uop_prs2;
  wire [6:0]  _slots_16_io_out_uop_prs3;
  wire [5:0]  _slots_16_io_out_uop_ppred;
  wire        _slots_16_io_out_uop_prs1_busy;
  wire        _slots_16_io_out_uop_prs2_busy;
  wire        _slots_16_io_out_uop_prs3_busy;
  wire        _slots_16_io_out_uop_ppred_busy;
  wire [6:0]  _slots_16_io_out_uop_stale_pdst;
  wire        _slots_16_io_out_uop_exception;
  wire [63:0] _slots_16_io_out_uop_exc_cause;
  wire        _slots_16_io_out_uop_bypassable;
  wire [4:0]  _slots_16_io_out_uop_mem_cmd;
  wire [1:0]  _slots_16_io_out_uop_mem_size;
  wire        _slots_16_io_out_uop_mem_signed;
  wire        _slots_16_io_out_uop_is_fence;
  wire        _slots_16_io_out_uop_is_fencei;
  wire        _slots_16_io_out_uop_is_amo;
  wire        _slots_16_io_out_uop_uses_ldq;
  wire        _slots_16_io_out_uop_uses_stq;
  wire        _slots_16_io_out_uop_is_sys_pc2epc;
  wire        _slots_16_io_out_uop_is_unique;
  wire        _slots_16_io_out_uop_flush_on_commit;
  wire        _slots_16_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_16_io_out_uop_ldst;
  wire [5:0]  _slots_16_io_out_uop_lrs1;
  wire [5:0]  _slots_16_io_out_uop_lrs2;
  wire [5:0]  _slots_16_io_out_uop_lrs3;
  wire        _slots_16_io_out_uop_ldst_val;
  wire [1:0]  _slots_16_io_out_uop_dst_rtype;
  wire [1:0]  _slots_16_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_16_io_out_uop_lrs2_rtype;
  wire        _slots_16_io_out_uop_frs3_en;
  wire        _slots_16_io_out_uop_fp_val;
  wire        _slots_16_io_out_uop_fp_single;
  wire        _slots_16_io_out_uop_xcpt_pf_if;
  wire        _slots_16_io_out_uop_xcpt_ae_if;
  wire        _slots_16_io_out_uop_xcpt_ma_if;
  wire        _slots_16_io_out_uop_bp_debug_if;
  wire        _slots_16_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_16_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_16_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_16_io_uop_uopc;
  wire [31:0] _slots_16_io_uop_inst;
  wire [31:0] _slots_16_io_uop_debug_inst;
  wire        _slots_16_io_uop_is_rvc;
  wire [39:0] _slots_16_io_uop_debug_pc;
  wire [2:0]  _slots_16_io_uop_iq_type;
  wire [9:0]  _slots_16_io_uop_fu_code;
  wire [1:0]  _slots_16_io_uop_iw_state;
  wire        _slots_16_io_uop_iw_p1_poisoned;
  wire        _slots_16_io_uop_iw_p2_poisoned;
  wire        _slots_16_io_uop_is_br;
  wire        _slots_16_io_uop_is_jalr;
  wire        _slots_16_io_uop_is_jal;
  wire        _slots_16_io_uop_is_sfb;
  wire [19:0] _slots_16_io_uop_br_mask;
  wire [4:0]  _slots_16_io_uop_br_tag;
  wire [5:0]  _slots_16_io_uop_ftq_idx;
  wire        _slots_16_io_uop_edge_inst;
  wire [5:0]  _slots_16_io_uop_pc_lob;
  wire        _slots_16_io_uop_taken;
  wire [19:0] _slots_16_io_uop_imm_packed;
  wire [11:0] _slots_16_io_uop_csr_addr;
  wire [6:0]  _slots_16_io_uop_rob_idx;
  wire [4:0]  _slots_16_io_uop_ldq_idx;
  wire [4:0]  _slots_16_io_uop_stq_idx;
  wire [1:0]  _slots_16_io_uop_rxq_idx;
  wire [6:0]  _slots_16_io_uop_pdst;
  wire [6:0]  _slots_16_io_uop_prs1;
  wire [6:0]  _slots_16_io_uop_prs2;
  wire [6:0]  _slots_16_io_uop_prs3;
  wire [5:0]  _slots_16_io_uop_ppred;
  wire        _slots_16_io_uop_prs1_busy;
  wire        _slots_16_io_uop_prs2_busy;
  wire        _slots_16_io_uop_prs3_busy;
  wire        _slots_16_io_uop_ppred_busy;
  wire [6:0]  _slots_16_io_uop_stale_pdst;
  wire        _slots_16_io_uop_exception;
  wire [63:0] _slots_16_io_uop_exc_cause;
  wire        _slots_16_io_uop_bypassable;
  wire [4:0]  _slots_16_io_uop_mem_cmd;
  wire [1:0]  _slots_16_io_uop_mem_size;
  wire        _slots_16_io_uop_mem_signed;
  wire        _slots_16_io_uop_is_fence;
  wire        _slots_16_io_uop_is_fencei;
  wire        _slots_16_io_uop_is_amo;
  wire        _slots_16_io_uop_uses_ldq;
  wire        _slots_16_io_uop_uses_stq;
  wire        _slots_16_io_uop_is_sys_pc2epc;
  wire        _slots_16_io_uop_is_unique;
  wire        _slots_16_io_uop_flush_on_commit;
  wire        _slots_16_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_16_io_uop_ldst;
  wire [5:0]  _slots_16_io_uop_lrs1;
  wire [5:0]  _slots_16_io_uop_lrs2;
  wire [5:0]  _slots_16_io_uop_lrs3;
  wire        _slots_16_io_uop_ldst_val;
  wire [1:0]  _slots_16_io_uop_dst_rtype;
  wire [1:0]  _slots_16_io_uop_lrs1_rtype;
  wire [1:0]  _slots_16_io_uop_lrs2_rtype;
  wire        _slots_16_io_uop_frs3_en;
  wire        _slots_16_io_uop_fp_val;
  wire        _slots_16_io_uop_fp_single;
  wire        _slots_16_io_uop_xcpt_pf_if;
  wire        _slots_16_io_uop_xcpt_ae_if;
  wire        _slots_16_io_uop_xcpt_ma_if;
  wire        _slots_16_io_uop_bp_debug_if;
  wire        _slots_16_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_16_io_uop_debug_fsrc;
  wire [1:0]  _slots_16_io_uop_debug_tsrc;
  wire        _slots_15_io_valid;
  wire        _slots_15_io_will_be_valid;
  wire        _slots_15_io_request;
  wire [6:0]  _slots_15_io_out_uop_uopc;
  wire [31:0] _slots_15_io_out_uop_inst;
  wire [31:0] _slots_15_io_out_uop_debug_inst;
  wire        _slots_15_io_out_uop_is_rvc;
  wire [39:0] _slots_15_io_out_uop_debug_pc;
  wire [2:0]  _slots_15_io_out_uop_iq_type;
  wire [9:0]  _slots_15_io_out_uop_fu_code;
  wire [1:0]  _slots_15_io_out_uop_iw_state;
  wire        _slots_15_io_out_uop_iw_p1_poisoned;
  wire        _slots_15_io_out_uop_iw_p2_poisoned;
  wire        _slots_15_io_out_uop_is_br;
  wire        _slots_15_io_out_uop_is_jalr;
  wire        _slots_15_io_out_uop_is_jal;
  wire        _slots_15_io_out_uop_is_sfb;
  wire [19:0] _slots_15_io_out_uop_br_mask;
  wire [4:0]  _slots_15_io_out_uop_br_tag;
  wire [5:0]  _slots_15_io_out_uop_ftq_idx;
  wire        _slots_15_io_out_uop_edge_inst;
  wire [5:0]  _slots_15_io_out_uop_pc_lob;
  wire        _slots_15_io_out_uop_taken;
  wire [19:0] _slots_15_io_out_uop_imm_packed;
  wire [11:0] _slots_15_io_out_uop_csr_addr;
  wire [6:0]  _slots_15_io_out_uop_rob_idx;
  wire [4:0]  _slots_15_io_out_uop_ldq_idx;
  wire [4:0]  _slots_15_io_out_uop_stq_idx;
  wire [1:0]  _slots_15_io_out_uop_rxq_idx;
  wire [6:0]  _slots_15_io_out_uop_pdst;
  wire [6:0]  _slots_15_io_out_uop_prs1;
  wire [6:0]  _slots_15_io_out_uop_prs2;
  wire [6:0]  _slots_15_io_out_uop_prs3;
  wire [5:0]  _slots_15_io_out_uop_ppred;
  wire        _slots_15_io_out_uop_prs1_busy;
  wire        _slots_15_io_out_uop_prs2_busy;
  wire        _slots_15_io_out_uop_prs3_busy;
  wire        _slots_15_io_out_uop_ppred_busy;
  wire [6:0]  _slots_15_io_out_uop_stale_pdst;
  wire        _slots_15_io_out_uop_exception;
  wire [63:0] _slots_15_io_out_uop_exc_cause;
  wire        _slots_15_io_out_uop_bypassable;
  wire [4:0]  _slots_15_io_out_uop_mem_cmd;
  wire [1:0]  _slots_15_io_out_uop_mem_size;
  wire        _slots_15_io_out_uop_mem_signed;
  wire        _slots_15_io_out_uop_is_fence;
  wire        _slots_15_io_out_uop_is_fencei;
  wire        _slots_15_io_out_uop_is_amo;
  wire        _slots_15_io_out_uop_uses_ldq;
  wire        _slots_15_io_out_uop_uses_stq;
  wire        _slots_15_io_out_uop_is_sys_pc2epc;
  wire        _slots_15_io_out_uop_is_unique;
  wire        _slots_15_io_out_uop_flush_on_commit;
  wire        _slots_15_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_15_io_out_uop_ldst;
  wire [5:0]  _slots_15_io_out_uop_lrs1;
  wire [5:0]  _slots_15_io_out_uop_lrs2;
  wire [5:0]  _slots_15_io_out_uop_lrs3;
  wire        _slots_15_io_out_uop_ldst_val;
  wire [1:0]  _slots_15_io_out_uop_dst_rtype;
  wire [1:0]  _slots_15_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_15_io_out_uop_lrs2_rtype;
  wire        _slots_15_io_out_uop_frs3_en;
  wire        _slots_15_io_out_uop_fp_val;
  wire        _slots_15_io_out_uop_fp_single;
  wire        _slots_15_io_out_uop_xcpt_pf_if;
  wire        _slots_15_io_out_uop_xcpt_ae_if;
  wire        _slots_15_io_out_uop_xcpt_ma_if;
  wire        _slots_15_io_out_uop_bp_debug_if;
  wire        _slots_15_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_15_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_15_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_15_io_uop_uopc;
  wire [31:0] _slots_15_io_uop_inst;
  wire [31:0] _slots_15_io_uop_debug_inst;
  wire        _slots_15_io_uop_is_rvc;
  wire [39:0] _slots_15_io_uop_debug_pc;
  wire [2:0]  _slots_15_io_uop_iq_type;
  wire [9:0]  _slots_15_io_uop_fu_code;
  wire [1:0]  _slots_15_io_uop_iw_state;
  wire        _slots_15_io_uop_iw_p1_poisoned;
  wire        _slots_15_io_uop_iw_p2_poisoned;
  wire        _slots_15_io_uop_is_br;
  wire        _slots_15_io_uop_is_jalr;
  wire        _slots_15_io_uop_is_jal;
  wire        _slots_15_io_uop_is_sfb;
  wire [19:0] _slots_15_io_uop_br_mask;
  wire [4:0]  _slots_15_io_uop_br_tag;
  wire [5:0]  _slots_15_io_uop_ftq_idx;
  wire        _slots_15_io_uop_edge_inst;
  wire [5:0]  _slots_15_io_uop_pc_lob;
  wire        _slots_15_io_uop_taken;
  wire [19:0] _slots_15_io_uop_imm_packed;
  wire [11:0] _slots_15_io_uop_csr_addr;
  wire [6:0]  _slots_15_io_uop_rob_idx;
  wire [4:0]  _slots_15_io_uop_ldq_idx;
  wire [4:0]  _slots_15_io_uop_stq_idx;
  wire [1:0]  _slots_15_io_uop_rxq_idx;
  wire [6:0]  _slots_15_io_uop_pdst;
  wire [6:0]  _slots_15_io_uop_prs1;
  wire [6:0]  _slots_15_io_uop_prs2;
  wire [6:0]  _slots_15_io_uop_prs3;
  wire [5:0]  _slots_15_io_uop_ppred;
  wire        _slots_15_io_uop_prs1_busy;
  wire        _slots_15_io_uop_prs2_busy;
  wire        _slots_15_io_uop_prs3_busy;
  wire        _slots_15_io_uop_ppred_busy;
  wire [6:0]  _slots_15_io_uop_stale_pdst;
  wire        _slots_15_io_uop_exception;
  wire [63:0] _slots_15_io_uop_exc_cause;
  wire        _slots_15_io_uop_bypassable;
  wire [4:0]  _slots_15_io_uop_mem_cmd;
  wire [1:0]  _slots_15_io_uop_mem_size;
  wire        _slots_15_io_uop_mem_signed;
  wire        _slots_15_io_uop_is_fence;
  wire        _slots_15_io_uop_is_fencei;
  wire        _slots_15_io_uop_is_amo;
  wire        _slots_15_io_uop_uses_ldq;
  wire        _slots_15_io_uop_uses_stq;
  wire        _slots_15_io_uop_is_sys_pc2epc;
  wire        _slots_15_io_uop_is_unique;
  wire        _slots_15_io_uop_flush_on_commit;
  wire        _slots_15_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_15_io_uop_ldst;
  wire [5:0]  _slots_15_io_uop_lrs1;
  wire [5:0]  _slots_15_io_uop_lrs2;
  wire [5:0]  _slots_15_io_uop_lrs3;
  wire        _slots_15_io_uop_ldst_val;
  wire [1:0]  _slots_15_io_uop_dst_rtype;
  wire [1:0]  _slots_15_io_uop_lrs1_rtype;
  wire [1:0]  _slots_15_io_uop_lrs2_rtype;
  wire        _slots_15_io_uop_frs3_en;
  wire        _slots_15_io_uop_fp_val;
  wire        _slots_15_io_uop_fp_single;
  wire        _slots_15_io_uop_xcpt_pf_if;
  wire        _slots_15_io_uop_xcpt_ae_if;
  wire        _slots_15_io_uop_xcpt_ma_if;
  wire        _slots_15_io_uop_bp_debug_if;
  wire        _slots_15_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_15_io_uop_debug_fsrc;
  wire [1:0]  _slots_15_io_uop_debug_tsrc;
  wire        _slots_14_io_valid;
  wire        _slots_14_io_will_be_valid;
  wire        _slots_14_io_request;
  wire [6:0]  _slots_14_io_out_uop_uopc;
  wire [31:0] _slots_14_io_out_uop_inst;
  wire [31:0] _slots_14_io_out_uop_debug_inst;
  wire        _slots_14_io_out_uop_is_rvc;
  wire [39:0] _slots_14_io_out_uop_debug_pc;
  wire [2:0]  _slots_14_io_out_uop_iq_type;
  wire [9:0]  _slots_14_io_out_uop_fu_code;
  wire [1:0]  _slots_14_io_out_uop_iw_state;
  wire        _slots_14_io_out_uop_iw_p1_poisoned;
  wire        _slots_14_io_out_uop_iw_p2_poisoned;
  wire        _slots_14_io_out_uop_is_br;
  wire        _slots_14_io_out_uop_is_jalr;
  wire        _slots_14_io_out_uop_is_jal;
  wire        _slots_14_io_out_uop_is_sfb;
  wire [19:0] _slots_14_io_out_uop_br_mask;
  wire [4:0]  _slots_14_io_out_uop_br_tag;
  wire [5:0]  _slots_14_io_out_uop_ftq_idx;
  wire        _slots_14_io_out_uop_edge_inst;
  wire [5:0]  _slots_14_io_out_uop_pc_lob;
  wire        _slots_14_io_out_uop_taken;
  wire [19:0] _slots_14_io_out_uop_imm_packed;
  wire [11:0] _slots_14_io_out_uop_csr_addr;
  wire [6:0]  _slots_14_io_out_uop_rob_idx;
  wire [4:0]  _slots_14_io_out_uop_ldq_idx;
  wire [4:0]  _slots_14_io_out_uop_stq_idx;
  wire [1:0]  _slots_14_io_out_uop_rxq_idx;
  wire [6:0]  _slots_14_io_out_uop_pdst;
  wire [6:0]  _slots_14_io_out_uop_prs1;
  wire [6:0]  _slots_14_io_out_uop_prs2;
  wire [6:0]  _slots_14_io_out_uop_prs3;
  wire [5:0]  _slots_14_io_out_uop_ppred;
  wire        _slots_14_io_out_uop_prs1_busy;
  wire        _slots_14_io_out_uop_prs2_busy;
  wire        _slots_14_io_out_uop_prs3_busy;
  wire        _slots_14_io_out_uop_ppred_busy;
  wire [6:0]  _slots_14_io_out_uop_stale_pdst;
  wire        _slots_14_io_out_uop_exception;
  wire [63:0] _slots_14_io_out_uop_exc_cause;
  wire        _slots_14_io_out_uop_bypassable;
  wire [4:0]  _slots_14_io_out_uop_mem_cmd;
  wire [1:0]  _slots_14_io_out_uop_mem_size;
  wire        _slots_14_io_out_uop_mem_signed;
  wire        _slots_14_io_out_uop_is_fence;
  wire        _slots_14_io_out_uop_is_fencei;
  wire        _slots_14_io_out_uop_is_amo;
  wire        _slots_14_io_out_uop_uses_ldq;
  wire        _slots_14_io_out_uop_uses_stq;
  wire        _slots_14_io_out_uop_is_sys_pc2epc;
  wire        _slots_14_io_out_uop_is_unique;
  wire        _slots_14_io_out_uop_flush_on_commit;
  wire        _slots_14_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_14_io_out_uop_ldst;
  wire [5:0]  _slots_14_io_out_uop_lrs1;
  wire [5:0]  _slots_14_io_out_uop_lrs2;
  wire [5:0]  _slots_14_io_out_uop_lrs3;
  wire        _slots_14_io_out_uop_ldst_val;
  wire [1:0]  _slots_14_io_out_uop_dst_rtype;
  wire [1:0]  _slots_14_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_14_io_out_uop_lrs2_rtype;
  wire        _slots_14_io_out_uop_frs3_en;
  wire        _slots_14_io_out_uop_fp_val;
  wire        _slots_14_io_out_uop_fp_single;
  wire        _slots_14_io_out_uop_xcpt_pf_if;
  wire        _slots_14_io_out_uop_xcpt_ae_if;
  wire        _slots_14_io_out_uop_xcpt_ma_if;
  wire        _slots_14_io_out_uop_bp_debug_if;
  wire        _slots_14_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_14_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_14_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_14_io_uop_uopc;
  wire [31:0] _slots_14_io_uop_inst;
  wire [31:0] _slots_14_io_uop_debug_inst;
  wire        _slots_14_io_uop_is_rvc;
  wire [39:0] _slots_14_io_uop_debug_pc;
  wire [2:0]  _slots_14_io_uop_iq_type;
  wire [9:0]  _slots_14_io_uop_fu_code;
  wire [1:0]  _slots_14_io_uop_iw_state;
  wire        _slots_14_io_uop_iw_p1_poisoned;
  wire        _slots_14_io_uop_iw_p2_poisoned;
  wire        _slots_14_io_uop_is_br;
  wire        _slots_14_io_uop_is_jalr;
  wire        _slots_14_io_uop_is_jal;
  wire        _slots_14_io_uop_is_sfb;
  wire [19:0] _slots_14_io_uop_br_mask;
  wire [4:0]  _slots_14_io_uop_br_tag;
  wire [5:0]  _slots_14_io_uop_ftq_idx;
  wire        _slots_14_io_uop_edge_inst;
  wire [5:0]  _slots_14_io_uop_pc_lob;
  wire        _slots_14_io_uop_taken;
  wire [19:0] _slots_14_io_uop_imm_packed;
  wire [11:0] _slots_14_io_uop_csr_addr;
  wire [6:0]  _slots_14_io_uop_rob_idx;
  wire [4:0]  _slots_14_io_uop_ldq_idx;
  wire [4:0]  _slots_14_io_uop_stq_idx;
  wire [1:0]  _slots_14_io_uop_rxq_idx;
  wire [6:0]  _slots_14_io_uop_pdst;
  wire [6:0]  _slots_14_io_uop_prs1;
  wire [6:0]  _slots_14_io_uop_prs2;
  wire [6:0]  _slots_14_io_uop_prs3;
  wire [5:0]  _slots_14_io_uop_ppred;
  wire        _slots_14_io_uop_prs1_busy;
  wire        _slots_14_io_uop_prs2_busy;
  wire        _slots_14_io_uop_prs3_busy;
  wire        _slots_14_io_uop_ppred_busy;
  wire [6:0]  _slots_14_io_uop_stale_pdst;
  wire        _slots_14_io_uop_exception;
  wire [63:0] _slots_14_io_uop_exc_cause;
  wire        _slots_14_io_uop_bypassable;
  wire [4:0]  _slots_14_io_uop_mem_cmd;
  wire [1:0]  _slots_14_io_uop_mem_size;
  wire        _slots_14_io_uop_mem_signed;
  wire        _slots_14_io_uop_is_fence;
  wire        _slots_14_io_uop_is_fencei;
  wire        _slots_14_io_uop_is_amo;
  wire        _slots_14_io_uop_uses_ldq;
  wire        _slots_14_io_uop_uses_stq;
  wire        _slots_14_io_uop_is_sys_pc2epc;
  wire        _slots_14_io_uop_is_unique;
  wire        _slots_14_io_uop_flush_on_commit;
  wire        _slots_14_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_14_io_uop_ldst;
  wire [5:0]  _slots_14_io_uop_lrs1;
  wire [5:0]  _slots_14_io_uop_lrs2;
  wire [5:0]  _slots_14_io_uop_lrs3;
  wire        _slots_14_io_uop_ldst_val;
  wire [1:0]  _slots_14_io_uop_dst_rtype;
  wire [1:0]  _slots_14_io_uop_lrs1_rtype;
  wire [1:0]  _slots_14_io_uop_lrs2_rtype;
  wire        _slots_14_io_uop_frs3_en;
  wire        _slots_14_io_uop_fp_val;
  wire        _slots_14_io_uop_fp_single;
  wire        _slots_14_io_uop_xcpt_pf_if;
  wire        _slots_14_io_uop_xcpt_ae_if;
  wire        _slots_14_io_uop_xcpt_ma_if;
  wire        _slots_14_io_uop_bp_debug_if;
  wire        _slots_14_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_14_io_uop_debug_fsrc;
  wire [1:0]  _slots_14_io_uop_debug_tsrc;
  wire        _slots_13_io_valid;
  wire        _slots_13_io_will_be_valid;
  wire        _slots_13_io_request;
  wire [6:0]  _slots_13_io_out_uop_uopc;
  wire [31:0] _slots_13_io_out_uop_inst;
  wire [31:0] _slots_13_io_out_uop_debug_inst;
  wire        _slots_13_io_out_uop_is_rvc;
  wire [39:0] _slots_13_io_out_uop_debug_pc;
  wire [2:0]  _slots_13_io_out_uop_iq_type;
  wire [9:0]  _slots_13_io_out_uop_fu_code;
  wire [1:0]  _slots_13_io_out_uop_iw_state;
  wire        _slots_13_io_out_uop_iw_p1_poisoned;
  wire        _slots_13_io_out_uop_iw_p2_poisoned;
  wire        _slots_13_io_out_uop_is_br;
  wire        _slots_13_io_out_uop_is_jalr;
  wire        _slots_13_io_out_uop_is_jal;
  wire        _slots_13_io_out_uop_is_sfb;
  wire [19:0] _slots_13_io_out_uop_br_mask;
  wire [4:0]  _slots_13_io_out_uop_br_tag;
  wire [5:0]  _slots_13_io_out_uop_ftq_idx;
  wire        _slots_13_io_out_uop_edge_inst;
  wire [5:0]  _slots_13_io_out_uop_pc_lob;
  wire        _slots_13_io_out_uop_taken;
  wire [19:0] _slots_13_io_out_uop_imm_packed;
  wire [11:0] _slots_13_io_out_uop_csr_addr;
  wire [6:0]  _slots_13_io_out_uop_rob_idx;
  wire [4:0]  _slots_13_io_out_uop_ldq_idx;
  wire [4:0]  _slots_13_io_out_uop_stq_idx;
  wire [1:0]  _slots_13_io_out_uop_rxq_idx;
  wire [6:0]  _slots_13_io_out_uop_pdst;
  wire [6:0]  _slots_13_io_out_uop_prs1;
  wire [6:0]  _slots_13_io_out_uop_prs2;
  wire [6:0]  _slots_13_io_out_uop_prs3;
  wire [5:0]  _slots_13_io_out_uop_ppred;
  wire        _slots_13_io_out_uop_prs1_busy;
  wire        _slots_13_io_out_uop_prs2_busy;
  wire        _slots_13_io_out_uop_prs3_busy;
  wire        _slots_13_io_out_uop_ppred_busy;
  wire [6:0]  _slots_13_io_out_uop_stale_pdst;
  wire        _slots_13_io_out_uop_exception;
  wire [63:0] _slots_13_io_out_uop_exc_cause;
  wire        _slots_13_io_out_uop_bypassable;
  wire [4:0]  _slots_13_io_out_uop_mem_cmd;
  wire [1:0]  _slots_13_io_out_uop_mem_size;
  wire        _slots_13_io_out_uop_mem_signed;
  wire        _slots_13_io_out_uop_is_fence;
  wire        _slots_13_io_out_uop_is_fencei;
  wire        _slots_13_io_out_uop_is_amo;
  wire        _slots_13_io_out_uop_uses_ldq;
  wire        _slots_13_io_out_uop_uses_stq;
  wire        _slots_13_io_out_uop_is_sys_pc2epc;
  wire        _slots_13_io_out_uop_is_unique;
  wire        _slots_13_io_out_uop_flush_on_commit;
  wire        _slots_13_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_13_io_out_uop_ldst;
  wire [5:0]  _slots_13_io_out_uop_lrs1;
  wire [5:0]  _slots_13_io_out_uop_lrs2;
  wire [5:0]  _slots_13_io_out_uop_lrs3;
  wire        _slots_13_io_out_uop_ldst_val;
  wire [1:0]  _slots_13_io_out_uop_dst_rtype;
  wire [1:0]  _slots_13_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_13_io_out_uop_lrs2_rtype;
  wire        _slots_13_io_out_uop_frs3_en;
  wire        _slots_13_io_out_uop_fp_val;
  wire        _slots_13_io_out_uop_fp_single;
  wire        _slots_13_io_out_uop_xcpt_pf_if;
  wire        _slots_13_io_out_uop_xcpt_ae_if;
  wire        _slots_13_io_out_uop_xcpt_ma_if;
  wire        _slots_13_io_out_uop_bp_debug_if;
  wire        _slots_13_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_13_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_13_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_13_io_uop_uopc;
  wire [31:0] _slots_13_io_uop_inst;
  wire [31:0] _slots_13_io_uop_debug_inst;
  wire        _slots_13_io_uop_is_rvc;
  wire [39:0] _slots_13_io_uop_debug_pc;
  wire [2:0]  _slots_13_io_uop_iq_type;
  wire [9:0]  _slots_13_io_uop_fu_code;
  wire [1:0]  _slots_13_io_uop_iw_state;
  wire        _slots_13_io_uop_iw_p1_poisoned;
  wire        _slots_13_io_uop_iw_p2_poisoned;
  wire        _slots_13_io_uop_is_br;
  wire        _slots_13_io_uop_is_jalr;
  wire        _slots_13_io_uop_is_jal;
  wire        _slots_13_io_uop_is_sfb;
  wire [19:0] _slots_13_io_uop_br_mask;
  wire [4:0]  _slots_13_io_uop_br_tag;
  wire [5:0]  _slots_13_io_uop_ftq_idx;
  wire        _slots_13_io_uop_edge_inst;
  wire [5:0]  _slots_13_io_uop_pc_lob;
  wire        _slots_13_io_uop_taken;
  wire [19:0] _slots_13_io_uop_imm_packed;
  wire [11:0] _slots_13_io_uop_csr_addr;
  wire [6:0]  _slots_13_io_uop_rob_idx;
  wire [4:0]  _slots_13_io_uop_ldq_idx;
  wire [4:0]  _slots_13_io_uop_stq_idx;
  wire [1:0]  _slots_13_io_uop_rxq_idx;
  wire [6:0]  _slots_13_io_uop_pdst;
  wire [6:0]  _slots_13_io_uop_prs1;
  wire [6:0]  _slots_13_io_uop_prs2;
  wire [6:0]  _slots_13_io_uop_prs3;
  wire [5:0]  _slots_13_io_uop_ppred;
  wire        _slots_13_io_uop_prs1_busy;
  wire        _slots_13_io_uop_prs2_busy;
  wire        _slots_13_io_uop_prs3_busy;
  wire        _slots_13_io_uop_ppred_busy;
  wire [6:0]  _slots_13_io_uop_stale_pdst;
  wire        _slots_13_io_uop_exception;
  wire [63:0] _slots_13_io_uop_exc_cause;
  wire        _slots_13_io_uop_bypassable;
  wire [4:0]  _slots_13_io_uop_mem_cmd;
  wire [1:0]  _slots_13_io_uop_mem_size;
  wire        _slots_13_io_uop_mem_signed;
  wire        _slots_13_io_uop_is_fence;
  wire        _slots_13_io_uop_is_fencei;
  wire        _slots_13_io_uop_is_amo;
  wire        _slots_13_io_uop_uses_ldq;
  wire        _slots_13_io_uop_uses_stq;
  wire        _slots_13_io_uop_is_sys_pc2epc;
  wire        _slots_13_io_uop_is_unique;
  wire        _slots_13_io_uop_flush_on_commit;
  wire        _slots_13_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_13_io_uop_ldst;
  wire [5:0]  _slots_13_io_uop_lrs1;
  wire [5:0]  _slots_13_io_uop_lrs2;
  wire [5:0]  _slots_13_io_uop_lrs3;
  wire        _slots_13_io_uop_ldst_val;
  wire [1:0]  _slots_13_io_uop_dst_rtype;
  wire [1:0]  _slots_13_io_uop_lrs1_rtype;
  wire [1:0]  _slots_13_io_uop_lrs2_rtype;
  wire        _slots_13_io_uop_frs3_en;
  wire        _slots_13_io_uop_fp_val;
  wire        _slots_13_io_uop_fp_single;
  wire        _slots_13_io_uop_xcpt_pf_if;
  wire        _slots_13_io_uop_xcpt_ae_if;
  wire        _slots_13_io_uop_xcpt_ma_if;
  wire        _slots_13_io_uop_bp_debug_if;
  wire        _slots_13_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_13_io_uop_debug_fsrc;
  wire [1:0]  _slots_13_io_uop_debug_tsrc;
  wire        _slots_12_io_valid;
  wire        _slots_12_io_will_be_valid;
  wire        _slots_12_io_request;
  wire [6:0]  _slots_12_io_out_uop_uopc;
  wire [31:0] _slots_12_io_out_uop_inst;
  wire [31:0] _slots_12_io_out_uop_debug_inst;
  wire        _slots_12_io_out_uop_is_rvc;
  wire [39:0] _slots_12_io_out_uop_debug_pc;
  wire [2:0]  _slots_12_io_out_uop_iq_type;
  wire [9:0]  _slots_12_io_out_uop_fu_code;
  wire [1:0]  _slots_12_io_out_uop_iw_state;
  wire        _slots_12_io_out_uop_iw_p1_poisoned;
  wire        _slots_12_io_out_uop_iw_p2_poisoned;
  wire        _slots_12_io_out_uop_is_br;
  wire        _slots_12_io_out_uop_is_jalr;
  wire        _slots_12_io_out_uop_is_jal;
  wire        _slots_12_io_out_uop_is_sfb;
  wire [19:0] _slots_12_io_out_uop_br_mask;
  wire [4:0]  _slots_12_io_out_uop_br_tag;
  wire [5:0]  _slots_12_io_out_uop_ftq_idx;
  wire        _slots_12_io_out_uop_edge_inst;
  wire [5:0]  _slots_12_io_out_uop_pc_lob;
  wire        _slots_12_io_out_uop_taken;
  wire [19:0] _slots_12_io_out_uop_imm_packed;
  wire [11:0] _slots_12_io_out_uop_csr_addr;
  wire [6:0]  _slots_12_io_out_uop_rob_idx;
  wire [4:0]  _slots_12_io_out_uop_ldq_idx;
  wire [4:0]  _slots_12_io_out_uop_stq_idx;
  wire [1:0]  _slots_12_io_out_uop_rxq_idx;
  wire [6:0]  _slots_12_io_out_uop_pdst;
  wire [6:0]  _slots_12_io_out_uop_prs1;
  wire [6:0]  _slots_12_io_out_uop_prs2;
  wire [6:0]  _slots_12_io_out_uop_prs3;
  wire [5:0]  _slots_12_io_out_uop_ppred;
  wire        _slots_12_io_out_uop_prs1_busy;
  wire        _slots_12_io_out_uop_prs2_busy;
  wire        _slots_12_io_out_uop_prs3_busy;
  wire        _slots_12_io_out_uop_ppred_busy;
  wire [6:0]  _slots_12_io_out_uop_stale_pdst;
  wire        _slots_12_io_out_uop_exception;
  wire [63:0] _slots_12_io_out_uop_exc_cause;
  wire        _slots_12_io_out_uop_bypassable;
  wire [4:0]  _slots_12_io_out_uop_mem_cmd;
  wire [1:0]  _slots_12_io_out_uop_mem_size;
  wire        _slots_12_io_out_uop_mem_signed;
  wire        _slots_12_io_out_uop_is_fence;
  wire        _slots_12_io_out_uop_is_fencei;
  wire        _slots_12_io_out_uop_is_amo;
  wire        _slots_12_io_out_uop_uses_ldq;
  wire        _slots_12_io_out_uop_uses_stq;
  wire        _slots_12_io_out_uop_is_sys_pc2epc;
  wire        _slots_12_io_out_uop_is_unique;
  wire        _slots_12_io_out_uop_flush_on_commit;
  wire        _slots_12_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_12_io_out_uop_ldst;
  wire [5:0]  _slots_12_io_out_uop_lrs1;
  wire [5:0]  _slots_12_io_out_uop_lrs2;
  wire [5:0]  _slots_12_io_out_uop_lrs3;
  wire        _slots_12_io_out_uop_ldst_val;
  wire [1:0]  _slots_12_io_out_uop_dst_rtype;
  wire [1:0]  _slots_12_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_12_io_out_uop_lrs2_rtype;
  wire        _slots_12_io_out_uop_frs3_en;
  wire        _slots_12_io_out_uop_fp_val;
  wire        _slots_12_io_out_uop_fp_single;
  wire        _slots_12_io_out_uop_xcpt_pf_if;
  wire        _slots_12_io_out_uop_xcpt_ae_if;
  wire        _slots_12_io_out_uop_xcpt_ma_if;
  wire        _slots_12_io_out_uop_bp_debug_if;
  wire        _slots_12_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_12_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_12_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_12_io_uop_uopc;
  wire [31:0] _slots_12_io_uop_inst;
  wire [31:0] _slots_12_io_uop_debug_inst;
  wire        _slots_12_io_uop_is_rvc;
  wire [39:0] _slots_12_io_uop_debug_pc;
  wire [2:0]  _slots_12_io_uop_iq_type;
  wire [9:0]  _slots_12_io_uop_fu_code;
  wire [1:0]  _slots_12_io_uop_iw_state;
  wire        _slots_12_io_uop_iw_p1_poisoned;
  wire        _slots_12_io_uop_iw_p2_poisoned;
  wire        _slots_12_io_uop_is_br;
  wire        _slots_12_io_uop_is_jalr;
  wire        _slots_12_io_uop_is_jal;
  wire        _slots_12_io_uop_is_sfb;
  wire [19:0] _slots_12_io_uop_br_mask;
  wire [4:0]  _slots_12_io_uop_br_tag;
  wire [5:0]  _slots_12_io_uop_ftq_idx;
  wire        _slots_12_io_uop_edge_inst;
  wire [5:0]  _slots_12_io_uop_pc_lob;
  wire        _slots_12_io_uop_taken;
  wire [19:0] _slots_12_io_uop_imm_packed;
  wire [11:0] _slots_12_io_uop_csr_addr;
  wire [6:0]  _slots_12_io_uop_rob_idx;
  wire [4:0]  _slots_12_io_uop_ldq_idx;
  wire [4:0]  _slots_12_io_uop_stq_idx;
  wire [1:0]  _slots_12_io_uop_rxq_idx;
  wire [6:0]  _slots_12_io_uop_pdst;
  wire [6:0]  _slots_12_io_uop_prs1;
  wire [6:0]  _slots_12_io_uop_prs2;
  wire [6:0]  _slots_12_io_uop_prs3;
  wire [5:0]  _slots_12_io_uop_ppred;
  wire        _slots_12_io_uop_prs1_busy;
  wire        _slots_12_io_uop_prs2_busy;
  wire        _slots_12_io_uop_prs3_busy;
  wire        _slots_12_io_uop_ppred_busy;
  wire [6:0]  _slots_12_io_uop_stale_pdst;
  wire        _slots_12_io_uop_exception;
  wire [63:0] _slots_12_io_uop_exc_cause;
  wire        _slots_12_io_uop_bypassable;
  wire [4:0]  _slots_12_io_uop_mem_cmd;
  wire [1:0]  _slots_12_io_uop_mem_size;
  wire        _slots_12_io_uop_mem_signed;
  wire        _slots_12_io_uop_is_fence;
  wire        _slots_12_io_uop_is_fencei;
  wire        _slots_12_io_uop_is_amo;
  wire        _slots_12_io_uop_uses_ldq;
  wire        _slots_12_io_uop_uses_stq;
  wire        _slots_12_io_uop_is_sys_pc2epc;
  wire        _slots_12_io_uop_is_unique;
  wire        _slots_12_io_uop_flush_on_commit;
  wire        _slots_12_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_12_io_uop_ldst;
  wire [5:0]  _slots_12_io_uop_lrs1;
  wire [5:0]  _slots_12_io_uop_lrs2;
  wire [5:0]  _slots_12_io_uop_lrs3;
  wire        _slots_12_io_uop_ldst_val;
  wire [1:0]  _slots_12_io_uop_dst_rtype;
  wire [1:0]  _slots_12_io_uop_lrs1_rtype;
  wire [1:0]  _slots_12_io_uop_lrs2_rtype;
  wire        _slots_12_io_uop_frs3_en;
  wire        _slots_12_io_uop_fp_val;
  wire        _slots_12_io_uop_fp_single;
  wire        _slots_12_io_uop_xcpt_pf_if;
  wire        _slots_12_io_uop_xcpt_ae_if;
  wire        _slots_12_io_uop_xcpt_ma_if;
  wire        _slots_12_io_uop_bp_debug_if;
  wire        _slots_12_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_12_io_uop_debug_fsrc;
  wire [1:0]  _slots_12_io_uop_debug_tsrc;
  wire        _slots_11_io_valid;
  wire        _slots_11_io_will_be_valid;
  wire        _slots_11_io_request;
  wire [6:0]  _slots_11_io_out_uop_uopc;
  wire [31:0] _slots_11_io_out_uop_inst;
  wire [31:0] _slots_11_io_out_uop_debug_inst;
  wire        _slots_11_io_out_uop_is_rvc;
  wire [39:0] _slots_11_io_out_uop_debug_pc;
  wire [2:0]  _slots_11_io_out_uop_iq_type;
  wire [9:0]  _slots_11_io_out_uop_fu_code;
  wire [1:0]  _slots_11_io_out_uop_iw_state;
  wire        _slots_11_io_out_uop_iw_p1_poisoned;
  wire        _slots_11_io_out_uop_iw_p2_poisoned;
  wire        _slots_11_io_out_uop_is_br;
  wire        _slots_11_io_out_uop_is_jalr;
  wire        _slots_11_io_out_uop_is_jal;
  wire        _slots_11_io_out_uop_is_sfb;
  wire [19:0] _slots_11_io_out_uop_br_mask;
  wire [4:0]  _slots_11_io_out_uop_br_tag;
  wire [5:0]  _slots_11_io_out_uop_ftq_idx;
  wire        _slots_11_io_out_uop_edge_inst;
  wire [5:0]  _slots_11_io_out_uop_pc_lob;
  wire        _slots_11_io_out_uop_taken;
  wire [19:0] _slots_11_io_out_uop_imm_packed;
  wire [11:0] _slots_11_io_out_uop_csr_addr;
  wire [6:0]  _slots_11_io_out_uop_rob_idx;
  wire [4:0]  _slots_11_io_out_uop_ldq_idx;
  wire [4:0]  _slots_11_io_out_uop_stq_idx;
  wire [1:0]  _slots_11_io_out_uop_rxq_idx;
  wire [6:0]  _slots_11_io_out_uop_pdst;
  wire [6:0]  _slots_11_io_out_uop_prs1;
  wire [6:0]  _slots_11_io_out_uop_prs2;
  wire [6:0]  _slots_11_io_out_uop_prs3;
  wire [5:0]  _slots_11_io_out_uop_ppred;
  wire        _slots_11_io_out_uop_prs1_busy;
  wire        _slots_11_io_out_uop_prs2_busy;
  wire        _slots_11_io_out_uop_prs3_busy;
  wire        _slots_11_io_out_uop_ppred_busy;
  wire [6:0]  _slots_11_io_out_uop_stale_pdst;
  wire        _slots_11_io_out_uop_exception;
  wire [63:0] _slots_11_io_out_uop_exc_cause;
  wire        _slots_11_io_out_uop_bypassable;
  wire [4:0]  _slots_11_io_out_uop_mem_cmd;
  wire [1:0]  _slots_11_io_out_uop_mem_size;
  wire        _slots_11_io_out_uop_mem_signed;
  wire        _slots_11_io_out_uop_is_fence;
  wire        _slots_11_io_out_uop_is_fencei;
  wire        _slots_11_io_out_uop_is_amo;
  wire        _slots_11_io_out_uop_uses_ldq;
  wire        _slots_11_io_out_uop_uses_stq;
  wire        _slots_11_io_out_uop_is_sys_pc2epc;
  wire        _slots_11_io_out_uop_is_unique;
  wire        _slots_11_io_out_uop_flush_on_commit;
  wire        _slots_11_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_11_io_out_uop_ldst;
  wire [5:0]  _slots_11_io_out_uop_lrs1;
  wire [5:0]  _slots_11_io_out_uop_lrs2;
  wire [5:0]  _slots_11_io_out_uop_lrs3;
  wire        _slots_11_io_out_uop_ldst_val;
  wire [1:0]  _slots_11_io_out_uop_dst_rtype;
  wire [1:0]  _slots_11_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_11_io_out_uop_lrs2_rtype;
  wire        _slots_11_io_out_uop_frs3_en;
  wire        _slots_11_io_out_uop_fp_val;
  wire        _slots_11_io_out_uop_fp_single;
  wire        _slots_11_io_out_uop_xcpt_pf_if;
  wire        _slots_11_io_out_uop_xcpt_ae_if;
  wire        _slots_11_io_out_uop_xcpt_ma_if;
  wire        _slots_11_io_out_uop_bp_debug_if;
  wire        _slots_11_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_11_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_11_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_11_io_uop_uopc;
  wire [31:0] _slots_11_io_uop_inst;
  wire [31:0] _slots_11_io_uop_debug_inst;
  wire        _slots_11_io_uop_is_rvc;
  wire [39:0] _slots_11_io_uop_debug_pc;
  wire [2:0]  _slots_11_io_uop_iq_type;
  wire [9:0]  _slots_11_io_uop_fu_code;
  wire [1:0]  _slots_11_io_uop_iw_state;
  wire        _slots_11_io_uop_iw_p1_poisoned;
  wire        _slots_11_io_uop_iw_p2_poisoned;
  wire        _slots_11_io_uop_is_br;
  wire        _slots_11_io_uop_is_jalr;
  wire        _slots_11_io_uop_is_jal;
  wire        _slots_11_io_uop_is_sfb;
  wire [19:0] _slots_11_io_uop_br_mask;
  wire [4:0]  _slots_11_io_uop_br_tag;
  wire [5:0]  _slots_11_io_uop_ftq_idx;
  wire        _slots_11_io_uop_edge_inst;
  wire [5:0]  _slots_11_io_uop_pc_lob;
  wire        _slots_11_io_uop_taken;
  wire [19:0] _slots_11_io_uop_imm_packed;
  wire [11:0] _slots_11_io_uop_csr_addr;
  wire [6:0]  _slots_11_io_uop_rob_idx;
  wire [4:0]  _slots_11_io_uop_ldq_idx;
  wire [4:0]  _slots_11_io_uop_stq_idx;
  wire [1:0]  _slots_11_io_uop_rxq_idx;
  wire [6:0]  _slots_11_io_uop_pdst;
  wire [6:0]  _slots_11_io_uop_prs1;
  wire [6:0]  _slots_11_io_uop_prs2;
  wire [6:0]  _slots_11_io_uop_prs3;
  wire [5:0]  _slots_11_io_uop_ppred;
  wire        _slots_11_io_uop_prs1_busy;
  wire        _slots_11_io_uop_prs2_busy;
  wire        _slots_11_io_uop_prs3_busy;
  wire        _slots_11_io_uop_ppred_busy;
  wire [6:0]  _slots_11_io_uop_stale_pdst;
  wire        _slots_11_io_uop_exception;
  wire [63:0] _slots_11_io_uop_exc_cause;
  wire        _slots_11_io_uop_bypassable;
  wire [4:0]  _slots_11_io_uop_mem_cmd;
  wire [1:0]  _slots_11_io_uop_mem_size;
  wire        _slots_11_io_uop_mem_signed;
  wire        _slots_11_io_uop_is_fence;
  wire        _slots_11_io_uop_is_fencei;
  wire        _slots_11_io_uop_is_amo;
  wire        _slots_11_io_uop_uses_ldq;
  wire        _slots_11_io_uop_uses_stq;
  wire        _slots_11_io_uop_is_sys_pc2epc;
  wire        _slots_11_io_uop_is_unique;
  wire        _slots_11_io_uop_flush_on_commit;
  wire        _slots_11_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_11_io_uop_ldst;
  wire [5:0]  _slots_11_io_uop_lrs1;
  wire [5:0]  _slots_11_io_uop_lrs2;
  wire [5:0]  _slots_11_io_uop_lrs3;
  wire        _slots_11_io_uop_ldst_val;
  wire [1:0]  _slots_11_io_uop_dst_rtype;
  wire [1:0]  _slots_11_io_uop_lrs1_rtype;
  wire [1:0]  _slots_11_io_uop_lrs2_rtype;
  wire        _slots_11_io_uop_frs3_en;
  wire        _slots_11_io_uop_fp_val;
  wire        _slots_11_io_uop_fp_single;
  wire        _slots_11_io_uop_xcpt_pf_if;
  wire        _slots_11_io_uop_xcpt_ae_if;
  wire        _slots_11_io_uop_xcpt_ma_if;
  wire        _slots_11_io_uop_bp_debug_if;
  wire        _slots_11_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_11_io_uop_debug_fsrc;
  wire [1:0]  _slots_11_io_uop_debug_tsrc;
  wire        _slots_10_io_valid;
  wire        _slots_10_io_will_be_valid;
  wire        _slots_10_io_request;
  wire [6:0]  _slots_10_io_out_uop_uopc;
  wire [31:0] _slots_10_io_out_uop_inst;
  wire [31:0] _slots_10_io_out_uop_debug_inst;
  wire        _slots_10_io_out_uop_is_rvc;
  wire [39:0] _slots_10_io_out_uop_debug_pc;
  wire [2:0]  _slots_10_io_out_uop_iq_type;
  wire [9:0]  _slots_10_io_out_uop_fu_code;
  wire [1:0]  _slots_10_io_out_uop_iw_state;
  wire        _slots_10_io_out_uop_iw_p1_poisoned;
  wire        _slots_10_io_out_uop_iw_p2_poisoned;
  wire        _slots_10_io_out_uop_is_br;
  wire        _slots_10_io_out_uop_is_jalr;
  wire        _slots_10_io_out_uop_is_jal;
  wire        _slots_10_io_out_uop_is_sfb;
  wire [19:0] _slots_10_io_out_uop_br_mask;
  wire [4:0]  _slots_10_io_out_uop_br_tag;
  wire [5:0]  _slots_10_io_out_uop_ftq_idx;
  wire        _slots_10_io_out_uop_edge_inst;
  wire [5:0]  _slots_10_io_out_uop_pc_lob;
  wire        _slots_10_io_out_uop_taken;
  wire [19:0] _slots_10_io_out_uop_imm_packed;
  wire [11:0] _slots_10_io_out_uop_csr_addr;
  wire [6:0]  _slots_10_io_out_uop_rob_idx;
  wire [4:0]  _slots_10_io_out_uop_ldq_idx;
  wire [4:0]  _slots_10_io_out_uop_stq_idx;
  wire [1:0]  _slots_10_io_out_uop_rxq_idx;
  wire [6:0]  _slots_10_io_out_uop_pdst;
  wire [6:0]  _slots_10_io_out_uop_prs1;
  wire [6:0]  _slots_10_io_out_uop_prs2;
  wire [6:0]  _slots_10_io_out_uop_prs3;
  wire [5:0]  _slots_10_io_out_uop_ppred;
  wire        _slots_10_io_out_uop_prs1_busy;
  wire        _slots_10_io_out_uop_prs2_busy;
  wire        _slots_10_io_out_uop_prs3_busy;
  wire        _slots_10_io_out_uop_ppred_busy;
  wire [6:0]  _slots_10_io_out_uop_stale_pdst;
  wire        _slots_10_io_out_uop_exception;
  wire [63:0] _slots_10_io_out_uop_exc_cause;
  wire        _slots_10_io_out_uop_bypassable;
  wire [4:0]  _slots_10_io_out_uop_mem_cmd;
  wire [1:0]  _slots_10_io_out_uop_mem_size;
  wire        _slots_10_io_out_uop_mem_signed;
  wire        _slots_10_io_out_uop_is_fence;
  wire        _slots_10_io_out_uop_is_fencei;
  wire        _slots_10_io_out_uop_is_amo;
  wire        _slots_10_io_out_uop_uses_ldq;
  wire        _slots_10_io_out_uop_uses_stq;
  wire        _slots_10_io_out_uop_is_sys_pc2epc;
  wire        _slots_10_io_out_uop_is_unique;
  wire        _slots_10_io_out_uop_flush_on_commit;
  wire        _slots_10_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_10_io_out_uop_ldst;
  wire [5:0]  _slots_10_io_out_uop_lrs1;
  wire [5:0]  _slots_10_io_out_uop_lrs2;
  wire [5:0]  _slots_10_io_out_uop_lrs3;
  wire        _slots_10_io_out_uop_ldst_val;
  wire [1:0]  _slots_10_io_out_uop_dst_rtype;
  wire [1:0]  _slots_10_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_10_io_out_uop_lrs2_rtype;
  wire        _slots_10_io_out_uop_frs3_en;
  wire        _slots_10_io_out_uop_fp_val;
  wire        _slots_10_io_out_uop_fp_single;
  wire        _slots_10_io_out_uop_xcpt_pf_if;
  wire        _slots_10_io_out_uop_xcpt_ae_if;
  wire        _slots_10_io_out_uop_xcpt_ma_if;
  wire        _slots_10_io_out_uop_bp_debug_if;
  wire        _slots_10_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_10_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_10_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_10_io_uop_uopc;
  wire [31:0] _slots_10_io_uop_inst;
  wire [31:0] _slots_10_io_uop_debug_inst;
  wire        _slots_10_io_uop_is_rvc;
  wire [39:0] _slots_10_io_uop_debug_pc;
  wire [2:0]  _slots_10_io_uop_iq_type;
  wire [9:0]  _slots_10_io_uop_fu_code;
  wire [1:0]  _slots_10_io_uop_iw_state;
  wire        _slots_10_io_uop_iw_p1_poisoned;
  wire        _slots_10_io_uop_iw_p2_poisoned;
  wire        _slots_10_io_uop_is_br;
  wire        _slots_10_io_uop_is_jalr;
  wire        _slots_10_io_uop_is_jal;
  wire        _slots_10_io_uop_is_sfb;
  wire [19:0] _slots_10_io_uop_br_mask;
  wire [4:0]  _slots_10_io_uop_br_tag;
  wire [5:0]  _slots_10_io_uop_ftq_idx;
  wire        _slots_10_io_uop_edge_inst;
  wire [5:0]  _slots_10_io_uop_pc_lob;
  wire        _slots_10_io_uop_taken;
  wire [19:0] _slots_10_io_uop_imm_packed;
  wire [11:0] _slots_10_io_uop_csr_addr;
  wire [6:0]  _slots_10_io_uop_rob_idx;
  wire [4:0]  _slots_10_io_uop_ldq_idx;
  wire [4:0]  _slots_10_io_uop_stq_idx;
  wire [1:0]  _slots_10_io_uop_rxq_idx;
  wire [6:0]  _slots_10_io_uop_pdst;
  wire [6:0]  _slots_10_io_uop_prs1;
  wire [6:0]  _slots_10_io_uop_prs2;
  wire [6:0]  _slots_10_io_uop_prs3;
  wire [5:0]  _slots_10_io_uop_ppred;
  wire        _slots_10_io_uop_prs1_busy;
  wire        _slots_10_io_uop_prs2_busy;
  wire        _slots_10_io_uop_prs3_busy;
  wire        _slots_10_io_uop_ppred_busy;
  wire [6:0]  _slots_10_io_uop_stale_pdst;
  wire        _slots_10_io_uop_exception;
  wire [63:0] _slots_10_io_uop_exc_cause;
  wire        _slots_10_io_uop_bypassable;
  wire [4:0]  _slots_10_io_uop_mem_cmd;
  wire [1:0]  _slots_10_io_uop_mem_size;
  wire        _slots_10_io_uop_mem_signed;
  wire        _slots_10_io_uop_is_fence;
  wire        _slots_10_io_uop_is_fencei;
  wire        _slots_10_io_uop_is_amo;
  wire        _slots_10_io_uop_uses_ldq;
  wire        _slots_10_io_uop_uses_stq;
  wire        _slots_10_io_uop_is_sys_pc2epc;
  wire        _slots_10_io_uop_is_unique;
  wire        _slots_10_io_uop_flush_on_commit;
  wire        _slots_10_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_10_io_uop_ldst;
  wire [5:0]  _slots_10_io_uop_lrs1;
  wire [5:0]  _slots_10_io_uop_lrs2;
  wire [5:0]  _slots_10_io_uop_lrs3;
  wire        _slots_10_io_uop_ldst_val;
  wire [1:0]  _slots_10_io_uop_dst_rtype;
  wire [1:0]  _slots_10_io_uop_lrs1_rtype;
  wire [1:0]  _slots_10_io_uop_lrs2_rtype;
  wire        _slots_10_io_uop_frs3_en;
  wire        _slots_10_io_uop_fp_val;
  wire        _slots_10_io_uop_fp_single;
  wire        _slots_10_io_uop_xcpt_pf_if;
  wire        _slots_10_io_uop_xcpt_ae_if;
  wire        _slots_10_io_uop_xcpt_ma_if;
  wire        _slots_10_io_uop_bp_debug_if;
  wire        _slots_10_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_10_io_uop_debug_fsrc;
  wire [1:0]  _slots_10_io_uop_debug_tsrc;
  wire        _slots_9_io_valid;
  wire        _slots_9_io_will_be_valid;
  wire        _slots_9_io_request;
  wire [6:0]  _slots_9_io_out_uop_uopc;
  wire [31:0] _slots_9_io_out_uop_inst;
  wire [31:0] _slots_9_io_out_uop_debug_inst;
  wire        _slots_9_io_out_uop_is_rvc;
  wire [39:0] _slots_9_io_out_uop_debug_pc;
  wire [2:0]  _slots_9_io_out_uop_iq_type;
  wire [9:0]  _slots_9_io_out_uop_fu_code;
  wire [1:0]  _slots_9_io_out_uop_iw_state;
  wire        _slots_9_io_out_uop_iw_p1_poisoned;
  wire        _slots_9_io_out_uop_iw_p2_poisoned;
  wire        _slots_9_io_out_uop_is_br;
  wire        _slots_9_io_out_uop_is_jalr;
  wire        _slots_9_io_out_uop_is_jal;
  wire        _slots_9_io_out_uop_is_sfb;
  wire [19:0] _slots_9_io_out_uop_br_mask;
  wire [4:0]  _slots_9_io_out_uop_br_tag;
  wire [5:0]  _slots_9_io_out_uop_ftq_idx;
  wire        _slots_9_io_out_uop_edge_inst;
  wire [5:0]  _slots_9_io_out_uop_pc_lob;
  wire        _slots_9_io_out_uop_taken;
  wire [19:0] _slots_9_io_out_uop_imm_packed;
  wire [11:0] _slots_9_io_out_uop_csr_addr;
  wire [6:0]  _slots_9_io_out_uop_rob_idx;
  wire [4:0]  _slots_9_io_out_uop_ldq_idx;
  wire [4:0]  _slots_9_io_out_uop_stq_idx;
  wire [1:0]  _slots_9_io_out_uop_rxq_idx;
  wire [6:0]  _slots_9_io_out_uop_pdst;
  wire [6:0]  _slots_9_io_out_uop_prs1;
  wire [6:0]  _slots_9_io_out_uop_prs2;
  wire [6:0]  _slots_9_io_out_uop_prs3;
  wire [5:0]  _slots_9_io_out_uop_ppred;
  wire        _slots_9_io_out_uop_prs1_busy;
  wire        _slots_9_io_out_uop_prs2_busy;
  wire        _slots_9_io_out_uop_prs3_busy;
  wire        _slots_9_io_out_uop_ppred_busy;
  wire [6:0]  _slots_9_io_out_uop_stale_pdst;
  wire        _slots_9_io_out_uop_exception;
  wire [63:0] _slots_9_io_out_uop_exc_cause;
  wire        _slots_9_io_out_uop_bypassable;
  wire [4:0]  _slots_9_io_out_uop_mem_cmd;
  wire [1:0]  _slots_9_io_out_uop_mem_size;
  wire        _slots_9_io_out_uop_mem_signed;
  wire        _slots_9_io_out_uop_is_fence;
  wire        _slots_9_io_out_uop_is_fencei;
  wire        _slots_9_io_out_uop_is_amo;
  wire        _slots_9_io_out_uop_uses_ldq;
  wire        _slots_9_io_out_uop_uses_stq;
  wire        _slots_9_io_out_uop_is_sys_pc2epc;
  wire        _slots_9_io_out_uop_is_unique;
  wire        _slots_9_io_out_uop_flush_on_commit;
  wire        _slots_9_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_9_io_out_uop_ldst;
  wire [5:0]  _slots_9_io_out_uop_lrs1;
  wire [5:0]  _slots_9_io_out_uop_lrs2;
  wire [5:0]  _slots_9_io_out_uop_lrs3;
  wire        _slots_9_io_out_uop_ldst_val;
  wire [1:0]  _slots_9_io_out_uop_dst_rtype;
  wire [1:0]  _slots_9_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_9_io_out_uop_lrs2_rtype;
  wire        _slots_9_io_out_uop_frs3_en;
  wire        _slots_9_io_out_uop_fp_val;
  wire        _slots_9_io_out_uop_fp_single;
  wire        _slots_9_io_out_uop_xcpt_pf_if;
  wire        _slots_9_io_out_uop_xcpt_ae_if;
  wire        _slots_9_io_out_uop_xcpt_ma_if;
  wire        _slots_9_io_out_uop_bp_debug_if;
  wire        _slots_9_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_9_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_9_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_9_io_uop_uopc;
  wire [31:0] _slots_9_io_uop_inst;
  wire [31:0] _slots_9_io_uop_debug_inst;
  wire        _slots_9_io_uop_is_rvc;
  wire [39:0] _slots_9_io_uop_debug_pc;
  wire [2:0]  _slots_9_io_uop_iq_type;
  wire [9:0]  _slots_9_io_uop_fu_code;
  wire [1:0]  _slots_9_io_uop_iw_state;
  wire        _slots_9_io_uop_iw_p1_poisoned;
  wire        _slots_9_io_uop_iw_p2_poisoned;
  wire        _slots_9_io_uop_is_br;
  wire        _slots_9_io_uop_is_jalr;
  wire        _slots_9_io_uop_is_jal;
  wire        _slots_9_io_uop_is_sfb;
  wire [19:0] _slots_9_io_uop_br_mask;
  wire [4:0]  _slots_9_io_uop_br_tag;
  wire [5:0]  _slots_9_io_uop_ftq_idx;
  wire        _slots_9_io_uop_edge_inst;
  wire [5:0]  _slots_9_io_uop_pc_lob;
  wire        _slots_9_io_uop_taken;
  wire [19:0] _slots_9_io_uop_imm_packed;
  wire [11:0] _slots_9_io_uop_csr_addr;
  wire [6:0]  _slots_9_io_uop_rob_idx;
  wire [4:0]  _slots_9_io_uop_ldq_idx;
  wire [4:0]  _slots_9_io_uop_stq_idx;
  wire [1:0]  _slots_9_io_uop_rxq_idx;
  wire [6:0]  _slots_9_io_uop_pdst;
  wire [6:0]  _slots_9_io_uop_prs1;
  wire [6:0]  _slots_9_io_uop_prs2;
  wire [6:0]  _slots_9_io_uop_prs3;
  wire [5:0]  _slots_9_io_uop_ppred;
  wire        _slots_9_io_uop_prs1_busy;
  wire        _slots_9_io_uop_prs2_busy;
  wire        _slots_9_io_uop_prs3_busy;
  wire        _slots_9_io_uop_ppred_busy;
  wire [6:0]  _slots_9_io_uop_stale_pdst;
  wire        _slots_9_io_uop_exception;
  wire [63:0] _slots_9_io_uop_exc_cause;
  wire        _slots_9_io_uop_bypassable;
  wire [4:0]  _slots_9_io_uop_mem_cmd;
  wire [1:0]  _slots_9_io_uop_mem_size;
  wire        _slots_9_io_uop_mem_signed;
  wire        _slots_9_io_uop_is_fence;
  wire        _slots_9_io_uop_is_fencei;
  wire        _slots_9_io_uop_is_amo;
  wire        _slots_9_io_uop_uses_ldq;
  wire        _slots_9_io_uop_uses_stq;
  wire        _slots_9_io_uop_is_sys_pc2epc;
  wire        _slots_9_io_uop_is_unique;
  wire        _slots_9_io_uop_flush_on_commit;
  wire        _slots_9_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_9_io_uop_ldst;
  wire [5:0]  _slots_9_io_uop_lrs1;
  wire [5:0]  _slots_9_io_uop_lrs2;
  wire [5:0]  _slots_9_io_uop_lrs3;
  wire        _slots_9_io_uop_ldst_val;
  wire [1:0]  _slots_9_io_uop_dst_rtype;
  wire [1:0]  _slots_9_io_uop_lrs1_rtype;
  wire [1:0]  _slots_9_io_uop_lrs2_rtype;
  wire        _slots_9_io_uop_frs3_en;
  wire        _slots_9_io_uop_fp_val;
  wire        _slots_9_io_uop_fp_single;
  wire        _slots_9_io_uop_xcpt_pf_if;
  wire        _slots_9_io_uop_xcpt_ae_if;
  wire        _slots_9_io_uop_xcpt_ma_if;
  wire        _slots_9_io_uop_bp_debug_if;
  wire        _slots_9_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_9_io_uop_debug_fsrc;
  wire [1:0]  _slots_9_io_uop_debug_tsrc;
  wire        _slots_8_io_valid;
  wire        _slots_8_io_will_be_valid;
  wire        _slots_8_io_request;
  wire [6:0]  _slots_8_io_out_uop_uopc;
  wire [31:0] _slots_8_io_out_uop_inst;
  wire [31:0] _slots_8_io_out_uop_debug_inst;
  wire        _slots_8_io_out_uop_is_rvc;
  wire [39:0] _slots_8_io_out_uop_debug_pc;
  wire [2:0]  _slots_8_io_out_uop_iq_type;
  wire [9:0]  _slots_8_io_out_uop_fu_code;
  wire [1:0]  _slots_8_io_out_uop_iw_state;
  wire        _slots_8_io_out_uop_iw_p1_poisoned;
  wire        _slots_8_io_out_uop_iw_p2_poisoned;
  wire        _slots_8_io_out_uop_is_br;
  wire        _slots_8_io_out_uop_is_jalr;
  wire        _slots_8_io_out_uop_is_jal;
  wire        _slots_8_io_out_uop_is_sfb;
  wire [19:0] _slots_8_io_out_uop_br_mask;
  wire [4:0]  _slots_8_io_out_uop_br_tag;
  wire [5:0]  _slots_8_io_out_uop_ftq_idx;
  wire        _slots_8_io_out_uop_edge_inst;
  wire [5:0]  _slots_8_io_out_uop_pc_lob;
  wire        _slots_8_io_out_uop_taken;
  wire [19:0] _slots_8_io_out_uop_imm_packed;
  wire [11:0] _slots_8_io_out_uop_csr_addr;
  wire [6:0]  _slots_8_io_out_uop_rob_idx;
  wire [4:0]  _slots_8_io_out_uop_ldq_idx;
  wire [4:0]  _slots_8_io_out_uop_stq_idx;
  wire [1:0]  _slots_8_io_out_uop_rxq_idx;
  wire [6:0]  _slots_8_io_out_uop_pdst;
  wire [6:0]  _slots_8_io_out_uop_prs1;
  wire [6:0]  _slots_8_io_out_uop_prs2;
  wire [6:0]  _slots_8_io_out_uop_prs3;
  wire [5:0]  _slots_8_io_out_uop_ppred;
  wire        _slots_8_io_out_uop_prs1_busy;
  wire        _slots_8_io_out_uop_prs2_busy;
  wire        _slots_8_io_out_uop_prs3_busy;
  wire        _slots_8_io_out_uop_ppred_busy;
  wire [6:0]  _slots_8_io_out_uop_stale_pdst;
  wire        _slots_8_io_out_uop_exception;
  wire [63:0] _slots_8_io_out_uop_exc_cause;
  wire        _slots_8_io_out_uop_bypassable;
  wire [4:0]  _slots_8_io_out_uop_mem_cmd;
  wire [1:0]  _slots_8_io_out_uop_mem_size;
  wire        _slots_8_io_out_uop_mem_signed;
  wire        _slots_8_io_out_uop_is_fence;
  wire        _slots_8_io_out_uop_is_fencei;
  wire        _slots_8_io_out_uop_is_amo;
  wire        _slots_8_io_out_uop_uses_ldq;
  wire        _slots_8_io_out_uop_uses_stq;
  wire        _slots_8_io_out_uop_is_sys_pc2epc;
  wire        _slots_8_io_out_uop_is_unique;
  wire        _slots_8_io_out_uop_flush_on_commit;
  wire        _slots_8_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_8_io_out_uop_ldst;
  wire [5:0]  _slots_8_io_out_uop_lrs1;
  wire [5:0]  _slots_8_io_out_uop_lrs2;
  wire [5:0]  _slots_8_io_out_uop_lrs3;
  wire        _slots_8_io_out_uop_ldst_val;
  wire [1:0]  _slots_8_io_out_uop_dst_rtype;
  wire [1:0]  _slots_8_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_8_io_out_uop_lrs2_rtype;
  wire        _slots_8_io_out_uop_frs3_en;
  wire        _slots_8_io_out_uop_fp_val;
  wire        _slots_8_io_out_uop_fp_single;
  wire        _slots_8_io_out_uop_xcpt_pf_if;
  wire        _slots_8_io_out_uop_xcpt_ae_if;
  wire        _slots_8_io_out_uop_xcpt_ma_if;
  wire        _slots_8_io_out_uop_bp_debug_if;
  wire        _slots_8_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_8_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_8_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_8_io_uop_uopc;
  wire [31:0] _slots_8_io_uop_inst;
  wire [31:0] _slots_8_io_uop_debug_inst;
  wire        _slots_8_io_uop_is_rvc;
  wire [39:0] _slots_8_io_uop_debug_pc;
  wire [2:0]  _slots_8_io_uop_iq_type;
  wire [9:0]  _slots_8_io_uop_fu_code;
  wire [1:0]  _slots_8_io_uop_iw_state;
  wire        _slots_8_io_uop_iw_p1_poisoned;
  wire        _slots_8_io_uop_iw_p2_poisoned;
  wire        _slots_8_io_uop_is_br;
  wire        _slots_8_io_uop_is_jalr;
  wire        _slots_8_io_uop_is_jal;
  wire        _slots_8_io_uop_is_sfb;
  wire [19:0] _slots_8_io_uop_br_mask;
  wire [4:0]  _slots_8_io_uop_br_tag;
  wire [5:0]  _slots_8_io_uop_ftq_idx;
  wire        _slots_8_io_uop_edge_inst;
  wire [5:0]  _slots_8_io_uop_pc_lob;
  wire        _slots_8_io_uop_taken;
  wire [19:0] _slots_8_io_uop_imm_packed;
  wire [11:0] _slots_8_io_uop_csr_addr;
  wire [6:0]  _slots_8_io_uop_rob_idx;
  wire [4:0]  _slots_8_io_uop_ldq_idx;
  wire [4:0]  _slots_8_io_uop_stq_idx;
  wire [1:0]  _slots_8_io_uop_rxq_idx;
  wire [6:0]  _slots_8_io_uop_pdst;
  wire [6:0]  _slots_8_io_uop_prs1;
  wire [6:0]  _slots_8_io_uop_prs2;
  wire [6:0]  _slots_8_io_uop_prs3;
  wire [5:0]  _slots_8_io_uop_ppred;
  wire        _slots_8_io_uop_prs1_busy;
  wire        _slots_8_io_uop_prs2_busy;
  wire        _slots_8_io_uop_prs3_busy;
  wire        _slots_8_io_uop_ppred_busy;
  wire [6:0]  _slots_8_io_uop_stale_pdst;
  wire        _slots_8_io_uop_exception;
  wire [63:0] _slots_8_io_uop_exc_cause;
  wire        _slots_8_io_uop_bypassable;
  wire [4:0]  _slots_8_io_uop_mem_cmd;
  wire [1:0]  _slots_8_io_uop_mem_size;
  wire        _slots_8_io_uop_mem_signed;
  wire        _slots_8_io_uop_is_fence;
  wire        _slots_8_io_uop_is_fencei;
  wire        _slots_8_io_uop_is_amo;
  wire        _slots_8_io_uop_uses_ldq;
  wire        _slots_8_io_uop_uses_stq;
  wire        _slots_8_io_uop_is_sys_pc2epc;
  wire        _slots_8_io_uop_is_unique;
  wire        _slots_8_io_uop_flush_on_commit;
  wire        _slots_8_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_8_io_uop_ldst;
  wire [5:0]  _slots_8_io_uop_lrs1;
  wire [5:0]  _slots_8_io_uop_lrs2;
  wire [5:0]  _slots_8_io_uop_lrs3;
  wire        _slots_8_io_uop_ldst_val;
  wire [1:0]  _slots_8_io_uop_dst_rtype;
  wire [1:0]  _slots_8_io_uop_lrs1_rtype;
  wire [1:0]  _slots_8_io_uop_lrs2_rtype;
  wire        _slots_8_io_uop_frs3_en;
  wire        _slots_8_io_uop_fp_val;
  wire        _slots_8_io_uop_fp_single;
  wire        _slots_8_io_uop_xcpt_pf_if;
  wire        _slots_8_io_uop_xcpt_ae_if;
  wire        _slots_8_io_uop_xcpt_ma_if;
  wire        _slots_8_io_uop_bp_debug_if;
  wire        _slots_8_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_8_io_uop_debug_fsrc;
  wire [1:0]  _slots_8_io_uop_debug_tsrc;
  wire        _slots_7_io_valid;
  wire        _slots_7_io_will_be_valid;
  wire        _slots_7_io_request;
  wire [6:0]  _slots_7_io_out_uop_uopc;
  wire [31:0] _slots_7_io_out_uop_inst;
  wire [31:0] _slots_7_io_out_uop_debug_inst;
  wire        _slots_7_io_out_uop_is_rvc;
  wire [39:0] _slots_7_io_out_uop_debug_pc;
  wire [2:0]  _slots_7_io_out_uop_iq_type;
  wire [9:0]  _slots_7_io_out_uop_fu_code;
  wire [1:0]  _slots_7_io_out_uop_iw_state;
  wire        _slots_7_io_out_uop_iw_p1_poisoned;
  wire        _slots_7_io_out_uop_iw_p2_poisoned;
  wire        _slots_7_io_out_uop_is_br;
  wire        _slots_7_io_out_uop_is_jalr;
  wire        _slots_7_io_out_uop_is_jal;
  wire        _slots_7_io_out_uop_is_sfb;
  wire [19:0] _slots_7_io_out_uop_br_mask;
  wire [4:0]  _slots_7_io_out_uop_br_tag;
  wire [5:0]  _slots_7_io_out_uop_ftq_idx;
  wire        _slots_7_io_out_uop_edge_inst;
  wire [5:0]  _slots_7_io_out_uop_pc_lob;
  wire        _slots_7_io_out_uop_taken;
  wire [19:0] _slots_7_io_out_uop_imm_packed;
  wire [11:0] _slots_7_io_out_uop_csr_addr;
  wire [6:0]  _slots_7_io_out_uop_rob_idx;
  wire [4:0]  _slots_7_io_out_uop_ldq_idx;
  wire [4:0]  _slots_7_io_out_uop_stq_idx;
  wire [1:0]  _slots_7_io_out_uop_rxq_idx;
  wire [6:0]  _slots_7_io_out_uop_pdst;
  wire [6:0]  _slots_7_io_out_uop_prs1;
  wire [6:0]  _slots_7_io_out_uop_prs2;
  wire [6:0]  _slots_7_io_out_uop_prs3;
  wire [5:0]  _slots_7_io_out_uop_ppred;
  wire        _slots_7_io_out_uop_prs1_busy;
  wire        _slots_7_io_out_uop_prs2_busy;
  wire        _slots_7_io_out_uop_prs3_busy;
  wire        _slots_7_io_out_uop_ppred_busy;
  wire [6:0]  _slots_7_io_out_uop_stale_pdst;
  wire        _slots_7_io_out_uop_exception;
  wire [63:0] _slots_7_io_out_uop_exc_cause;
  wire        _slots_7_io_out_uop_bypassable;
  wire [4:0]  _slots_7_io_out_uop_mem_cmd;
  wire [1:0]  _slots_7_io_out_uop_mem_size;
  wire        _slots_7_io_out_uop_mem_signed;
  wire        _slots_7_io_out_uop_is_fence;
  wire        _slots_7_io_out_uop_is_fencei;
  wire        _slots_7_io_out_uop_is_amo;
  wire        _slots_7_io_out_uop_uses_ldq;
  wire        _slots_7_io_out_uop_uses_stq;
  wire        _slots_7_io_out_uop_is_sys_pc2epc;
  wire        _slots_7_io_out_uop_is_unique;
  wire        _slots_7_io_out_uop_flush_on_commit;
  wire        _slots_7_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_7_io_out_uop_ldst;
  wire [5:0]  _slots_7_io_out_uop_lrs1;
  wire [5:0]  _slots_7_io_out_uop_lrs2;
  wire [5:0]  _slots_7_io_out_uop_lrs3;
  wire        _slots_7_io_out_uop_ldst_val;
  wire [1:0]  _slots_7_io_out_uop_dst_rtype;
  wire [1:0]  _slots_7_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_7_io_out_uop_lrs2_rtype;
  wire        _slots_7_io_out_uop_frs3_en;
  wire        _slots_7_io_out_uop_fp_val;
  wire        _slots_7_io_out_uop_fp_single;
  wire        _slots_7_io_out_uop_xcpt_pf_if;
  wire        _slots_7_io_out_uop_xcpt_ae_if;
  wire        _slots_7_io_out_uop_xcpt_ma_if;
  wire        _slots_7_io_out_uop_bp_debug_if;
  wire        _slots_7_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_7_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_7_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_7_io_uop_uopc;
  wire [31:0] _slots_7_io_uop_inst;
  wire [31:0] _slots_7_io_uop_debug_inst;
  wire        _slots_7_io_uop_is_rvc;
  wire [39:0] _slots_7_io_uop_debug_pc;
  wire [2:0]  _slots_7_io_uop_iq_type;
  wire [9:0]  _slots_7_io_uop_fu_code;
  wire [1:0]  _slots_7_io_uop_iw_state;
  wire        _slots_7_io_uop_iw_p1_poisoned;
  wire        _slots_7_io_uop_iw_p2_poisoned;
  wire        _slots_7_io_uop_is_br;
  wire        _slots_7_io_uop_is_jalr;
  wire        _slots_7_io_uop_is_jal;
  wire        _slots_7_io_uop_is_sfb;
  wire [19:0] _slots_7_io_uop_br_mask;
  wire [4:0]  _slots_7_io_uop_br_tag;
  wire [5:0]  _slots_7_io_uop_ftq_idx;
  wire        _slots_7_io_uop_edge_inst;
  wire [5:0]  _slots_7_io_uop_pc_lob;
  wire        _slots_7_io_uop_taken;
  wire [19:0] _slots_7_io_uop_imm_packed;
  wire [11:0] _slots_7_io_uop_csr_addr;
  wire [6:0]  _slots_7_io_uop_rob_idx;
  wire [4:0]  _slots_7_io_uop_ldq_idx;
  wire [4:0]  _slots_7_io_uop_stq_idx;
  wire [1:0]  _slots_7_io_uop_rxq_idx;
  wire [6:0]  _slots_7_io_uop_pdst;
  wire [6:0]  _slots_7_io_uop_prs1;
  wire [6:0]  _slots_7_io_uop_prs2;
  wire [6:0]  _slots_7_io_uop_prs3;
  wire [5:0]  _slots_7_io_uop_ppred;
  wire        _slots_7_io_uop_prs1_busy;
  wire        _slots_7_io_uop_prs2_busy;
  wire        _slots_7_io_uop_prs3_busy;
  wire        _slots_7_io_uop_ppred_busy;
  wire [6:0]  _slots_7_io_uop_stale_pdst;
  wire        _slots_7_io_uop_exception;
  wire [63:0] _slots_7_io_uop_exc_cause;
  wire        _slots_7_io_uop_bypassable;
  wire [4:0]  _slots_7_io_uop_mem_cmd;
  wire [1:0]  _slots_7_io_uop_mem_size;
  wire        _slots_7_io_uop_mem_signed;
  wire        _slots_7_io_uop_is_fence;
  wire        _slots_7_io_uop_is_fencei;
  wire        _slots_7_io_uop_is_amo;
  wire        _slots_7_io_uop_uses_ldq;
  wire        _slots_7_io_uop_uses_stq;
  wire        _slots_7_io_uop_is_sys_pc2epc;
  wire        _slots_7_io_uop_is_unique;
  wire        _slots_7_io_uop_flush_on_commit;
  wire        _slots_7_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_7_io_uop_ldst;
  wire [5:0]  _slots_7_io_uop_lrs1;
  wire [5:0]  _slots_7_io_uop_lrs2;
  wire [5:0]  _slots_7_io_uop_lrs3;
  wire        _slots_7_io_uop_ldst_val;
  wire [1:0]  _slots_7_io_uop_dst_rtype;
  wire [1:0]  _slots_7_io_uop_lrs1_rtype;
  wire [1:0]  _slots_7_io_uop_lrs2_rtype;
  wire        _slots_7_io_uop_frs3_en;
  wire        _slots_7_io_uop_fp_val;
  wire        _slots_7_io_uop_fp_single;
  wire        _slots_7_io_uop_xcpt_pf_if;
  wire        _slots_7_io_uop_xcpt_ae_if;
  wire        _slots_7_io_uop_xcpt_ma_if;
  wire        _slots_7_io_uop_bp_debug_if;
  wire        _slots_7_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_7_io_uop_debug_fsrc;
  wire [1:0]  _slots_7_io_uop_debug_tsrc;
  wire        _slots_6_io_valid;
  wire        _slots_6_io_will_be_valid;
  wire        _slots_6_io_request;
  wire [6:0]  _slots_6_io_out_uop_uopc;
  wire [31:0] _slots_6_io_out_uop_inst;
  wire [31:0] _slots_6_io_out_uop_debug_inst;
  wire        _slots_6_io_out_uop_is_rvc;
  wire [39:0] _slots_6_io_out_uop_debug_pc;
  wire [2:0]  _slots_6_io_out_uop_iq_type;
  wire [9:0]  _slots_6_io_out_uop_fu_code;
  wire [1:0]  _slots_6_io_out_uop_iw_state;
  wire        _slots_6_io_out_uop_iw_p1_poisoned;
  wire        _slots_6_io_out_uop_iw_p2_poisoned;
  wire        _slots_6_io_out_uop_is_br;
  wire        _slots_6_io_out_uop_is_jalr;
  wire        _slots_6_io_out_uop_is_jal;
  wire        _slots_6_io_out_uop_is_sfb;
  wire [19:0] _slots_6_io_out_uop_br_mask;
  wire [4:0]  _slots_6_io_out_uop_br_tag;
  wire [5:0]  _slots_6_io_out_uop_ftq_idx;
  wire        _slots_6_io_out_uop_edge_inst;
  wire [5:0]  _slots_6_io_out_uop_pc_lob;
  wire        _slots_6_io_out_uop_taken;
  wire [19:0] _slots_6_io_out_uop_imm_packed;
  wire [11:0] _slots_6_io_out_uop_csr_addr;
  wire [6:0]  _slots_6_io_out_uop_rob_idx;
  wire [4:0]  _slots_6_io_out_uop_ldq_idx;
  wire [4:0]  _slots_6_io_out_uop_stq_idx;
  wire [1:0]  _slots_6_io_out_uop_rxq_idx;
  wire [6:0]  _slots_6_io_out_uop_pdst;
  wire [6:0]  _slots_6_io_out_uop_prs1;
  wire [6:0]  _slots_6_io_out_uop_prs2;
  wire [6:0]  _slots_6_io_out_uop_prs3;
  wire [5:0]  _slots_6_io_out_uop_ppred;
  wire        _slots_6_io_out_uop_prs1_busy;
  wire        _slots_6_io_out_uop_prs2_busy;
  wire        _slots_6_io_out_uop_prs3_busy;
  wire        _slots_6_io_out_uop_ppred_busy;
  wire [6:0]  _slots_6_io_out_uop_stale_pdst;
  wire        _slots_6_io_out_uop_exception;
  wire [63:0] _slots_6_io_out_uop_exc_cause;
  wire        _slots_6_io_out_uop_bypassable;
  wire [4:0]  _slots_6_io_out_uop_mem_cmd;
  wire [1:0]  _slots_6_io_out_uop_mem_size;
  wire        _slots_6_io_out_uop_mem_signed;
  wire        _slots_6_io_out_uop_is_fence;
  wire        _slots_6_io_out_uop_is_fencei;
  wire        _slots_6_io_out_uop_is_amo;
  wire        _slots_6_io_out_uop_uses_ldq;
  wire        _slots_6_io_out_uop_uses_stq;
  wire        _slots_6_io_out_uop_is_sys_pc2epc;
  wire        _slots_6_io_out_uop_is_unique;
  wire        _slots_6_io_out_uop_flush_on_commit;
  wire        _slots_6_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_6_io_out_uop_ldst;
  wire [5:0]  _slots_6_io_out_uop_lrs1;
  wire [5:0]  _slots_6_io_out_uop_lrs2;
  wire [5:0]  _slots_6_io_out_uop_lrs3;
  wire        _slots_6_io_out_uop_ldst_val;
  wire [1:0]  _slots_6_io_out_uop_dst_rtype;
  wire [1:0]  _slots_6_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_6_io_out_uop_lrs2_rtype;
  wire        _slots_6_io_out_uop_frs3_en;
  wire        _slots_6_io_out_uop_fp_val;
  wire        _slots_6_io_out_uop_fp_single;
  wire        _slots_6_io_out_uop_xcpt_pf_if;
  wire        _slots_6_io_out_uop_xcpt_ae_if;
  wire        _slots_6_io_out_uop_xcpt_ma_if;
  wire        _slots_6_io_out_uop_bp_debug_if;
  wire        _slots_6_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_6_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_6_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_6_io_uop_uopc;
  wire [31:0] _slots_6_io_uop_inst;
  wire [31:0] _slots_6_io_uop_debug_inst;
  wire        _slots_6_io_uop_is_rvc;
  wire [39:0] _slots_6_io_uop_debug_pc;
  wire [2:0]  _slots_6_io_uop_iq_type;
  wire [9:0]  _slots_6_io_uop_fu_code;
  wire [1:0]  _slots_6_io_uop_iw_state;
  wire        _slots_6_io_uop_iw_p1_poisoned;
  wire        _slots_6_io_uop_iw_p2_poisoned;
  wire        _slots_6_io_uop_is_br;
  wire        _slots_6_io_uop_is_jalr;
  wire        _slots_6_io_uop_is_jal;
  wire        _slots_6_io_uop_is_sfb;
  wire [19:0] _slots_6_io_uop_br_mask;
  wire [4:0]  _slots_6_io_uop_br_tag;
  wire [5:0]  _slots_6_io_uop_ftq_idx;
  wire        _slots_6_io_uop_edge_inst;
  wire [5:0]  _slots_6_io_uop_pc_lob;
  wire        _slots_6_io_uop_taken;
  wire [19:0] _slots_6_io_uop_imm_packed;
  wire [11:0] _slots_6_io_uop_csr_addr;
  wire [6:0]  _slots_6_io_uop_rob_idx;
  wire [4:0]  _slots_6_io_uop_ldq_idx;
  wire [4:0]  _slots_6_io_uop_stq_idx;
  wire [1:0]  _slots_6_io_uop_rxq_idx;
  wire [6:0]  _slots_6_io_uop_pdst;
  wire [6:0]  _slots_6_io_uop_prs1;
  wire [6:0]  _slots_6_io_uop_prs2;
  wire [6:0]  _slots_6_io_uop_prs3;
  wire [5:0]  _slots_6_io_uop_ppred;
  wire        _slots_6_io_uop_prs1_busy;
  wire        _slots_6_io_uop_prs2_busy;
  wire        _slots_6_io_uop_prs3_busy;
  wire        _slots_6_io_uop_ppred_busy;
  wire [6:0]  _slots_6_io_uop_stale_pdst;
  wire        _slots_6_io_uop_exception;
  wire [63:0] _slots_6_io_uop_exc_cause;
  wire        _slots_6_io_uop_bypassable;
  wire [4:0]  _slots_6_io_uop_mem_cmd;
  wire [1:0]  _slots_6_io_uop_mem_size;
  wire        _slots_6_io_uop_mem_signed;
  wire        _slots_6_io_uop_is_fence;
  wire        _slots_6_io_uop_is_fencei;
  wire        _slots_6_io_uop_is_amo;
  wire        _slots_6_io_uop_uses_ldq;
  wire        _slots_6_io_uop_uses_stq;
  wire        _slots_6_io_uop_is_sys_pc2epc;
  wire        _slots_6_io_uop_is_unique;
  wire        _slots_6_io_uop_flush_on_commit;
  wire        _slots_6_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_6_io_uop_ldst;
  wire [5:0]  _slots_6_io_uop_lrs1;
  wire [5:0]  _slots_6_io_uop_lrs2;
  wire [5:0]  _slots_6_io_uop_lrs3;
  wire        _slots_6_io_uop_ldst_val;
  wire [1:0]  _slots_6_io_uop_dst_rtype;
  wire [1:0]  _slots_6_io_uop_lrs1_rtype;
  wire [1:0]  _slots_6_io_uop_lrs2_rtype;
  wire        _slots_6_io_uop_frs3_en;
  wire        _slots_6_io_uop_fp_val;
  wire        _slots_6_io_uop_fp_single;
  wire        _slots_6_io_uop_xcpt_pf_if;
  wire        _slots_6_io_uop_xcpt_ae_if;
  wire        _slots_6_io_uop_xcpt_ma_if;
  wire        _slots_6_io_uop_bp_debug_if;
  wire        _slots_6_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_6_io_uop_debug_fsrc;
  wire [1:0]  _slots_6_io_uop_debug_tsrc;
  wire        _slots_5_io_valid;
  wire        _slots_5_io_will_be_valid;
  wire        _slots_5_io_request;
  wire [6:0]  _slots_5_io_out_uop_uopc;
  wire [31:0] _slots_5_io_out_uop_inst;
  wire [31:0] _slots_5_io_out_uop_debug_inst;
  wire        _slots_5_io_out_uop_is_rvc;
  wire [39:0] _slots_5_io_out_uop_debug_pc;
  wire [2:0]  _slots_5_io_out_uop_iq_type;
  wire [9:0]  _slots_5_io_out_uop_fu_code;
  wire [1:0]  _slots_5_io_out_uop_iw_state;
  wire        _slots_5_io_out_uop_iw_p1_poisoned;
  wire        _slots_5_io_out_uop_iw_p2_poisoned;
  wire        _slots_5_io_out_uop_is_br;
  wire        _slots_5_io_out_uop_is_jalr;
  wire        _slots_5_io_out_uop_is_jal;
  wire        _slots_5_io_out_uop_is_sfb;
  wire [19:0] _slots_5_io_out_uop_br_mask;
  wire [4:0]  _slots_5_io_out_uop_br_tag;
  wire [5:0]  _slots_5_io_out_uop_ftq_idx;
  wire        _slots_5_io_out_uop_edge_inst;
  wire [5:0]  _slots_5_io_out_uop_pc_lob;
  wire        _slots_5_io_out_uop_taken;
  wire [19:0] _slots_5_io_out_uop_imm_packed;
  wire [11:0] _slots_5_io_out_uop_csr_addr;
  wire [6:0]  _slots_5_io_out_uop_rob_idx;
  wire [4:0]  _slots_5_io_out_uop_ldq_idx;
  wire [4:0]  _slots_5_io_out_uop_stq_idx;
  wire [1:0]  _slots_5_io_out_uop_rxq_idx;
  wire [6:0]  _slots_5_io_out_uop_pdst;
  wire [6:0]  _slots_5_io_out_uop_prs1;
  wire [6:0]  _slots_5_io_out_uop_prs2;
  wire [6:0]  _slots_5_io_out_uop_prs3;
  wire [5:0]  _slots_5_io_out_uop_ppred;
  wire        _slots_5_io_out_uop_prs1_busy;
  wire        _slots_5_io_out_uop_prs2_busy;
  wire        _slots_5_io_out_uop_prs3_busy;
  wire        _slots_5_io_out_uop_ppred_busy;
  wire [6:0]  _slots_5_io_out_uop_stale_pdst;
  wire        _slots_5_io_out_uop_exception;
  wire [63:0] _slots_5_io_out_uop_exc_cause;
  wire        _slots_5_io_out_uop_bypassable;
  wire [4:0]  _slots_5_io_out_uop_mem_cmd;
  wire [1:0]  _slots_5_io_out_uop_mem_size;
  wire        _slots_5_io_out_uop_mem_signed;
  wire        _slots_5_io_out_uop_is_fence;
  wire        _slots_5_io_out_uop_is_fencei;
  wire        _slots_5_io_out_uop_is_amo;
  wire        _slots_5_io_out_uop_uses_ldq;
  wire        _slots_5_io_out_uop_uses_stq;
  wire        _slots_5_io_out_uop_is_sys_pc2epc;
  wire        _slots_5_io_out_uop_is_unique;
  wire        _slots_5_io_out_uop_flush_on_commit;
  wire        _slots_5_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_5_io_out_uop_ldst;
  wire [5:0]  _slots_5_io_out_uop_lrs1;
  wire [5:0]  _slots_5_io_out_uop_lrs2;
  wire [5:0]  _slots_5_io_out_uop_lrs3;
  wire        _slots_5_io_out_uop_ldst_val;
  wire [1:0]  _slots_5_io_out_uop_dst_rtype;
  wire [1:0]  _slots_5_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_5_io_out_uop_lrs2_rtype;
  wire        _slots_5_io_out_uop_frs3_en;
  wire        _slots_5_io_out_uop_fp_val;
  wire        _slots_5_io_out_uop_fp_single;
  wire        _slots_5_io_out_uop_xcpt_pf_if;
  wire        _slots_5_io_out_uop_xcpt_ae_if;
  wire        _slots_5_io_out_uop_xcpt_ma_if;
  wire        _slots_5_io_out_uop_bp_debug_if;
  wire        _slots_5_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_5_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_5_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_5_io_uop_uopc;
  wire [31:0] _slots_5_io_uop_inst;
  wire [31:0] _slots_5_io_uop_debug_inst;
  wire        _slots_5_io_uop_is_rvc;
  wire [39:0] _slots_5_io_uop_debug_pc;
  wire [2:0]  _slots_5_io_uop_iq_type;
  wire [9:0]  _slots_5_io_uop_fu_code;
  wire [1:0]  _slots_5_io_uop_iw_state;
  wire        _slots_5_io_uop_iw_p1_poisoned;
  wire        _slots_5_io_uop_iw_p2_poisoned;
  wire        _slots_5_io_uop_is_br;
  wire        _slots_5_io_uop_is_jalr;
  wire        _slots_5_io_uop_is_jal;
  wire        _slots_5_io_uop_is_sfb;
  wire [19:0] _slots_5_io_uop_br_mask;
  wire [4:0]  _slots_5_io_uop_br_tag;
  wire [5:0]  _slots_5_io_uop_ftq_idx;
  wire        _slots_5_io_uop_edge_inst;
  wire [5:0]  _slots_5_io_uop_pc_lob;
  wire        _slots_5_io_uop_taken;
  wire [19:0] _slots_5_io_uop_imm_packed;
  wire [11:0] _slots_5_io_uop_csr_addr;
  wire [6:0]  _slots_5_io_uop_rob_idx;
  wire [4:0]  _slots_5_io_uop_ldq_idx;
  wire [4:0]  _slots_5_io_uop_stq_idx;
  wire [1:0]  _slots_5_io_uop_rxq_idx;
  wire [6:0]  _slots_5_io_uop_pdst;
  wire [6:0]  _slots_5_io_uop_prs1;
  wire [6:0]  _slots_5_io_uop_prs2;
  wire [6:0]  _slots_5_io_uop_prs3;
  wire [5:0]  _slots_5_io_uop_ppred;
  wire        _slots_5_io_uop_prs1_busy;
  wire        _slots_5_io_uop_prs2_busy;
  wire        _slots_5_io_uop_prs3_busy;
  wire        _slots_5_io_uop_ppred_busy;
  wire [6:0]  _slots_5_io_uop_stale_pdst;
  wire        _slots_5_io_uop_exception;
  wire [63:0] _slots_5_io_uop_exc_cause;
  wire        _slots_5_io_uop_bypassable;
  wire [4:0]  _slots_5_io_uop_mem_cmd;
  wire [1:0]  _slots_5_io_uop_mem_size;
  wire        _slots_5_io_uop_mem_signed;
  wire        _slots_5_io_uop_is_fence;
  wire        _slots_5_io_uop_is_fencei;
  wire        _slots_5_io_uop_is_amo;
  wire        _slots_5_io_uop_uses_ldq;
  wire        _slots_5_io_uop_uses_stq;
  wire        _slots_5_io_uop_is_sys_pc2epc;
  wire        _slots_5_io_uop_is_unique;
  wire        _slots_5_io_uop_flush_on_commit;
  wire        _slots_5_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_5_io_uop_ldst;
  wire [5:0]  _slots_5_io_uop_lrs1;
  wire [5:0]  _slots_5_io_uop_lrs2;
  wire [5:0]  _slots_5_io_uop_lrs3;
  wire        _slots_5_io_uop_ldst_val;
  wire [1:0]  _slots_5_io_uop_dst_rtype;
  wire [1:0]  _slots_5_io_uop_lrs1_rtype;
  wire [1:0]  _slots_5_io_uop_lrs2_rtype;
  wire        _slots_5_io_uop_frs3_en;
  wire        _slots_5_io_uop_fp_val;
  wire        _slots_5_io_uop_fp_single;
  wire        _slots_5_io_uop_xcpt_pf_if;
  wire        _slots_5_io_uop_xcpt_ae_if;
  wire        _slots_5_io_uop_xcpt_ma_if;
  wire        _slots_5_io_uop_bp_debug_if;
  wire        _slots_5_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_5_io_uop_debug_fsrc;
  wire [1:0]  _slots_5_io_uop_debug_tsrc;
  wire        _slots_4_io_valid;
  wire        _slots_4_io_will_be_valid;
  wire        _slots_4_io_request;
  wire [6:0]  _slots_4_io_out_uop_uopc;
  wire [31:0] _slots_4_io_out_uop_inst;
  wire [31:0] _slots_4_io_out_uop_debug_inst;
  wire        _slots_4_io_out_uop_is_rvc;
  wire [39:0] _slots_4_io_out_uop_debug_pc;
  wire [2:0]  _slots_4_io_out_uop_iq_type;
  wire [9:0]  _slots_4_io_out_uop_fu_code;
  wire [1:0]  _slots_4_io_out_uop_iw_state;
  wire        _slots_4_io_out_uop_iw_p1_poisoned;
  wire        _slots_4_io_out_uop_iw_p2_poisoned;
  wire        _slots_4_io_out_uop_is_br;
  wire        _slots_4_io_out_uop_is_jalr;
  wire        _slots_4_io_out_uop_is_jal;
  wire        _slots_4_io_out_uop_is_sfb;
  wire [19:0] _slots_4_io_out_uop_br_mask;
  wire [4:0]  _slots_4_io_out_uop_br_tag;
  wire [5:0]  _slots_4_io_out_uop_ftq_idx;
  wire        _slots_4_io_out_uop_edge_inst;
  wire [5:0]  _slots_4_io_out_uop_pc_lob;
  wire        _slots_4_io_out_uop_taken;
  wire [19:0] _slots_4_io_out_uop_imm_packed;
  wire [11:0] _slots_4_io_out_uop_csr_addr;
  wire [6:0]  _slots_4_io_out_uop_rob_idx;
  wire [4:0]  _slots_4_io_out_uop_ldq_idx;
  wire [4:0]  _slots_4_io_out_uop_stq_idx;
  wire [1:0]  _slots_4_io_out_uop_rxq_idx;
  wire [6:0]  _slots_4_io_out_uop_pdst;
  wire [6:0]  _slots_4_io_out_uop_prs1;
  wire [6:0]  _slots_4_io_out_uop_prs2;
  wire [6:0]  _slots_4_io_out_uop_prs3;
  wire [5:0]  _slots_4_io_out_uop_ppred;
  wire        _slots_4_io_out_uop_prs1_busy;
  wire        _slots_4_io_out_uop_prs2_busy;
  wire        _slots_4_io_out_uop_prs3_busy;
  wire        _slots_4_io_out_uop_ppred_busy;
  wire [6:0]  _slots_4_io_out_uop_stale_pdst;
  wire        _slots_4_io_out_uop_exception;
  wire [63:0] _slots_4_io_out_uop_exc_cause;
  wire        _slots_4_io_out_uop_bypassable;
  wire [4:0]  _slots_4_io_out_uop_mem_cmd;
  wire [1:0]  _slots_4_io_out_uop_mem_size;
  wire        _slots_4_io_out_uop_mem_signed;
  wire        _slots_4_io_out_uop_is_fence;
  wire        _slots_4_io_out_uop_is_fencei;
  wire        _slots_4_io_out_uop_is_amo;
  wire        _slots_4_io_out_uop_uses_ldq;
  wire        _slots_4_io_out_uop_uses_stq;
  wire        _slots_4_io_out_uop_is_sys_pc2epc;
  wire        _slots_4_io_out_uop_is_unique;
  wire        _slots_4_io_out_uop_flush_on_commit;
  wire        _slots_4_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_4_io_out_uop_ldst;
  wire [5:0]  _slots_4_io_out_uop_lrs1;
  wire [5:0]  _slots_4_io_out_uop_lrs2;
  wire [5:0]  _slots_4_io_out_uop_lrs3;
  wire        _slots_4_io_out_uop_ldst_val;
  wire [1:0]  _slots_4_io_out_uop_dst_rtype;
  wire [1:0]  _slots_4_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_4_io_out_uop_lrs2_rtype;
  wire        _slots_4_io_out_uop_frs3_en;
  wire        _slots_4_io_out_uop_fp_val;
  wire        _slots_4_io_out_uop_fp_single;
  wire        _slots_4_io_out_uop_xcpt_pf_if;
  wire        _slots_4_io_out_uop_xcpt_ae_if;
  wire        _slots_4_io_out_uop_xcpt_ma_if;
  wire        _slots_4_io_out_uop_bp_debug_if;
  wire        _slots_4_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_4_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_4_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_4_io_uop_uopc;
  wire [31:0] _slots_4_io_uop_inst;
  wire [31:0] _slots_4_io_uop_debug_inst;
  wire        _slots_4_io_uop_is_rvc;
  wire [39:0] _slots_4_io_uop_debug_pc;
  wire [2:0]  _slots_4_io_uop_iq_type;
  wire [9:0]  _slots_4_io_uop_fu_code;
  wire [1:0]  _slots_4_io_uop_iw_state;
  wire        _slots_4_io_uop_iw_p1_poisoned;
  wire        _slots_4_io_uop_iw_p2_poisoned;
  wire        _slots_4_io_uop_is_br;
  wire        _slots_4_io_uop_is_jalr;
  wire        _slots_4_io_uop_is_jal;
  wire        _slots_4_io_uop_is_sfb;
  wire [19:0] _slots_4_io_uop_br_mask;
  wire [4:0]  _slots_4_io_uop_br_tag;
  wire [5:0]  _slots_4_io_uop_ftq_idx;
  wire        _slots_4_io_uop_edge_inst;
  wire [5:0]  _slots_4_io_uop_pc_lob;
  wire        _slots_4_io_uop_taken;
  wire [19:0] _slots_4_io_uop_imm_packed;
  wire [11:0] _slots_4_io_uop_csr_addr;
  wire [6:0]  _slots_4_io_uop_rob_idx;
  wire [4:0]  _slots_4_io_uop_ldq_idx;
  wire [4:0]  _slots_4_io_uop_stq_idx;
  wire [1:0]  _slots_4_io_uop_rxq_idx;
  wire [6:0]  _slots_4_io_uop_pdst;
  wire [6:0]  _slots_4_io_uop_prs1;
  wire [6:0]  _slots_4_io_uop_prs2;
  wire [6:0]  _slots_4_io_uop_prs3;
  wire [5:0]  _slots_4_io_uop_ppred;
  wire        _slots_4_io_uop_prs1_busy;
  wire        _slots_4_io_uop_prs2_busy;
  wire        _slots_4_io_uop_prs3_busy;
  wire        _slots_4_io_uop_ppred_busy;
  wire [6:0]  _slots_4_io_uop_stale_pdst;
  wire        _slots_4_io_uop_exception;
  wire [63:0] _slots_4_io_uop_exc_cause;
  wire        _slots_4_io_uop_bypassable;
  wire [4:0]  _slots_4_io_uop_mem_cmd;
  wire [1:0]  _slots_4_io_uop_mem_size;
  wire        _slots_4_io_uop_mem_signed;
  wire        _slots_4_io_uop_is_fence;
  wire        _slots_4_io_uop_is_fencei;
  wire        _slots_4_io_uop_is_amo;
  wire        _slots_4_io_uop_uses_ldq;
  wire        _slots_4_io_uop_uses_stq;
  wire        _slots_4_io_uop_is_sys_pc2epc;
  wire        _slots_4_io_uop_is_unique;
  wire        _slots_4_io_uop_flush_on_commit;
  wire        _slots_4_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_4_io_uop_ldst;
  wire [5:0]  _slots_4_io_uop_lrs1;
  wire [5:0]  _slots_4_io_uop_lrs2;
  wire [5:0]  _slots_4_io_uop_lrs3;
  wire        _slots_4_io_uop_ldst_val;
  wire [1:0]  _slots_4_io_uop_dst_rtype;
  wire [1:0]  _slots_4_io_uop_lrs1_rtype;
  wire [1:0]  _slots_4_io_uop_lrs2_rtype;
  wire        _slots_4_io_uop_frs3_en;
  wire        _slots_4_io_uop_fp_val;
  wire        _slots_4_io_uop_fp_single;
  wire        _slots_4_io_uop_xcpt_pf_if;
  wire        _slots_4_io_uop_xcpt_ae_if;
  wire        _slots_4_io_uop_xcpt_ma_if;
  wire        _slots_4_io_uop_bp_debug_if;
  wire        _slots_4_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_4_io_uop_debug_fsrc;
  wire [1:0]  _slots_4_io_uop_debug_tsrc;
  wire        _slots_3_io_valid;
  wire        _slots_3_io_will_be_valid;
  wire        _slots_3_io_request;
  wire [6:0]  _slots_3_io_out_uop_uopc;
  wire [31:0] _slots_3_io_out_uop_inst;
  wire [31:0] _slots_3_io_out_uop_debug_inst;
  wire        _slots_3_io_out_uop_is_rvc;
  wire [39:0] _slots_3_io_out_uop_debug_pc;
  wire [2:0]  _slots_3_io_out_uop_iq_type;
  wire [9:0]  _slots_3_io_out_uop_fu_code;
  wire [1:0]  _slots_3_io_out_uop_iw_state;
  wire        _slots_3_io_out_uop_iw_p1_poisoned;
  wire        _slots_3_io_out_uop_iw_p2_poisoned;
  wire        _slots_3_io_out_uop_is_br;
  wire        _slots_3_io_out_uop_is_jalr;
  wire        _slots_3_io_out_uop_is_jal;
  wire        _slots_3_io_out_uop_is_sfb;
  wire [19:0] _slots_3_io_out_uop_br_mask;
  wire [4:0]  _slots_3_io_out_uop_br_tag;
  wire [5:0]  _slots_3_io_out_uop_ftq_idx;
  wire        _slots_3_io_out_uop_edge_inst;
  wire [5:0]  _slots_3_io_out_uop_pc_lob;
  wire        _slots_3_io_out_uop_taken;
  wire [19:0] _slots_3_io_out_uop_imm_packed;
  wire [11:0] _slots_3_io_out_uop_csr_addr;
  wire [6:0]  _slots_3_io_out_uop_rob_idx;
  wire [4:0]  _slots_3_io_out_uop_ldq_idx;
  wire [4:0]  _slots_3_io_out_uop_stq_idx;
  wire [1:0]  _slots_3_io_out_uop_rxq_idx;
  wire [6:0]  _slots_3_io_out_uop_pdst;
  wire [6:0]  _slots_3_io_out_uop_prs1;
  wire [6:0]  _slots_3_io_out_uop_prs2;
  wire [6:0]  _slots_3_io_out_uop_prs3;
  wire [5:0]  _slots_3_io_out_uop_ppred;
  wire        _slots_3_io_out_uop_prs1_busy;
  wire        _slots_3_io_out_uop_prs2_busy;
  wire        _slots_3_io_out_uop_prs3_busy;
  wire        _slots_3_io_out_uop_ppred_busy;
  wire [6:0]  _slots_3_io_out_uop_stale_pdst;
  wire        _slots_3_io_out_uop_exception;
  wire [63:0] _slots_3_io_out_uop_exc_cause;
  wire        _slots_3_io_out_uop_bypassable;
  wire [4:0]  _slots_3_io_out_uop_mem_cmd;
  wire [1:0]  _slots_3_io_out_uop_mem_size;
  wire        _slots_3_io_out_uop_mem_signed;
  wire        _slots_3_io_out_uop_is_fence;
  wire        _slots_3_io_out_uop_is_fencei;
  wire        _slots_3_io_out_uop_is_amo;
  wire        _slots_3_io_out_uop_uses_ldq;
  wire        _slots_3_io_out_uop_uses_stq;
  wire        _slots_3_io_out_uop_is_sys_pc2epc;
  wire        _slots_3_io_out_uop_is_unique;
  wire        _slots_3_io_out_uop_flush_on_commit;
  wire        _slots_3_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_3_io_out_uop_ldst;
  wire [5:0]  _slots_3_io_out_uop_lrs1;
  wire [5:0]  _slots_3_io_out_uop_lrs2;
  wire [5:0]  _slots_3_io_out_uop_lrs3;
  wire        _slots_3_io_out_uop_ldst_val;
  wire [1:0]  _slots_3_io_out_uop_dst_rtype;
  wire [1:0]  _slots_3_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_3_io_out_uop_lrs2_rtype;
  wire        _slots_3_io_out_uop_frs3_en;
  wire        _slots_3_io_out_uop_fp_val;
  wire        _slots_3_io_out_uop_fp_single;
  wire        _slots_3_io_out_uop_xcpt_pf_if;
  wire        _slots_3_io_out_uop_xcpt_ae_if;
  wire        _slots_3_io_out_uop_xcpt_ma_if;
  wire        _slots_3_io_out_uop_bp_debug_if;
  wire        _slots_3_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_3_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_3_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_3_io_uop_uopc;
  wire [31:0] _slots_3_io_uop_inst;
  wire [31:0] _slots_3_io_uop_debug_inst;
  wire        _slots_3_io_uop_is_rvc;
  wire [39:0] _slots_3_io_uop_debug_pc;
  wire [2:0]  _slots_3_io_uop_iq_type;
  wire [9:0]  _slots_3_io_uop_fu_code;
  wire [1:0]  _slots_3_io_uop_iw_state;
  wire        _slots_3_io_uop_iw_p1_poisoned;
  wire        _slots_3_io_uop_iw_p2_poisoned;
  wire        _slots_3_io_uop_is_br;
  wire        _slots_3_io_uop_is_jalr;
  wire        _slots_3_io_uop_is_jal;
  wire        _slots_3_io_uop_is_sfb;
  wire [19:0] _slots_3_io_uop_br_mask;
  wire [4:0]  _slots_3_io_uop_br_tag;
  wire [5:0]  _slots_3_io_uop_ftq_idx;
  wire        _slots_3_io_uop_edge_inst;
  wire [5:0]  _slots_3_io_uop_pc_lob;
  wire        _slots_3_io_uop_taken;
  wire [19:0] _slots_3_io_uop_imm_packed;
  wire [11:0] _slots_3_io_uop_csr_addr;
  wire [6:0]  _slots_3_io_uop_rob_idx;
  wire [4:0]  _slots_3_io_uop_ldq_idx;
  wire [4:0]  _slots_3_io_uop_stq_idx;
  wire [1:0]  _slots_3_io_uop_rxq_idx;
  wire [6:0]  _slots_3_io_uop_pdst;
  wire [6:0]  _slots_3_io_uop_prs1;
  wire [6:0]  _slots_3_io_uop_prs2;
  wire [6:0]  _slots_3_io_uop_prs3;
  wire [5:0]  _slots_3_io_uop_ppred;
  wire        _slots_3_io_uop_prs1_busy;
  wire        _slots_3_io_uop_prs2_busy;
  wire        _slots_3_io_uop_prs3_busy;
  wire        _slots_3_io_uop_ppred_busy;
  wire [6:0]  _slots_3_io_uop_stale_pdst;
  wire        _slots_3_io_uop_exception;
  wire [63:0] _slots_3_io_uop_exc_cause;
  wire        _slots_3_io_uop_bypassable;
  wire [4:0]  _slots_3_io_uop_mem_cmd;
  wire [1:0]  _slots_3_io_uop_mem_size;
  wire        _slots_3_io_uop_mem_signed;
  wire        _slots_3_io_uop_is_fence;
  wire        _slots_3_io_uop_is_fencei;
  wire        _slots_3_io_uop_is_amo;
  wire        _slots_3_io_uop_uses_ldq;
  wire        _slots_3_io_uop_uses_stq;
  wire        _slots_3_io_uop_is_sys_pc2epc;
  wire        _slots_3_io_uop_is_unique;
  wire        _slots_3_io_uop_flush_on_commit;
  wire        _slots_3_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_3_io_uop_ldst;
  wire [5:0]  _slots_3_io_uop_lrs1;
  wire [5:0]  _slots_3_io_uop_lrs2;
  wire [5:0]  _slots_3_io_uop_lrs3;
  wire        _slots_3_io_uop_ldst_val;
  wire [1:0]  _slots_3_io_uop_dst_rtype;
  wire [1:0]  _slots_3_io_uop_lrs1_rtype;
  wire [1:0]  _slots_3_io_uop_lrs2_rtype;
  wire        _slots_3_io_uop_frs3_en;
  wire        _slots_3_io_uop_fp_val;
  wire        _slots_3_io_uop_fp_single;
  wire        _slots_3_io_uop_xcpt_pf_if;
  wire        _slots_3_io_uop_xcpt_ae_if;
  wire        _slots_3_io_uop_xcpt_ma_if;
  wire        _slots_3_io_uop_bp_debug_if;
  wire        _slots_3_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_3_io_uop_debug_fsrc;
  wire [1:0]  _slots_3_io_uop_debug_tsrc;
  wire        _slots_2_io_valid;
  wire        _slots_2_io_will_be_valid;
  wire        _slots_2_io_request;
  wire [6:0]  _slots_2_io_out_uop_uopc;
  wire [31:0] _slots_2_io_out_uop_inst;
  wire [31:0] _slots_2_io_out_uop_debug_inst;
  wire        _slots_2_io_out_uop_is_rvc;
  wire [39:0] _slots_2_io_out_uop_debug_pc;
  wire [2:0]  _slots_2_io_out_uop_iq_type;
  wire [9:0]  _slots_2_io_out_uop_fu_code;
  wire [1:0]  _slots_2_io_out_uop_iw_state;
  wire        _slots_2_io_out_uop_iw_p1_poisoned;
  wire        _slots_2_io_out_uop_iw_p2_poisoned;
  wire        _slots_2_io_out_uop_is_br;
  wire        _slots_2_io_out_uop_is_jalr;
  wire        _slots_2_io_out_uop_is_jal;
  wire        _slots_2_io_out_uop_is_sfb;
  wire [19:0] _slots_2_io_out_uop_br_mask;
  wire [4:0]  _slots_2_io_out_uop_br_tag;
  wire [5:0]  _slots_2_io_out_uop_ftq_idx;
  wire        _slots_2_io_out_uop_edge_inst;
  wire [5:0]  _slots_2_io_out_uop_pc_lob;
  wire        _slots_2_io_out_uop_taken;
  wire [19:0] _slots_2_io_out_uop_imm_packed;
  wire [11:0] _slots_2_io_out_uop_csr_addr;
  wire [6:0]  _slots_2_io_out_uop_rob_idx;
  wire [4:0]  _slots_2_io_out_uop_ldq_idx;
  wire [4:0]  _slots_2_io_out_uop_stq_idx;
  wire [1:0]  _slots_2_io_out_uop_rxq_idx;
  wire [6:0]  _slots_2_io_out_uop_pdst;
  wire [6:0]  _slots_2_io_out_uop_prs1;
  wire [6:0]  _slots_2_io_out_uop_prs2;
  wire [6:0]  _slots_2_io_out_uop_prs3;
  wire [5:0]  _slots_2_io_out_uop_ppred;
  wire        _slots_2_io_out_uop_prs1_busy;
  wire        _slots_2_io_out_uop_prs2_busy;
  wire        _slots_2_io_out_uop_prs3_busy;
  wire        _slots_2_io_out_uop_ppred_busy;
  wire [6:0]  _slots_2_io_out_uop_stale_pdst;
  wire        _slots_2_io_out_uop_exception;
  wire [63:0] _slots_2_io_out_uop_exc_cause;
  wire        _slots_2_io_out_uop_bypassable;
  wire [4:0]  _slots_2_io_out_uop_mem_cmd;
  wire [1:0]  _slots_2_io_out_uop_mem_size;
  wire        _slots_2_io_out_uop_mem_signed;
  wire        _slots_2_io_out_uop_is_fence;
  wire        _slots_2_io_out_uop_is_fencei;
  wire        _slots_2_io_out_uop_is_amo;
  wire        _slots_2_io_out_uop_uses_ldq;
  wire        _slots_2_io_out_uop_uses_stq;
  wire        _slots_2_io_out_uop_is_sys_pc2epc;
  wire        _slots_2_io_out_uop_is_unique;
  wire        _slots_2_io_out_uop_flush_on_commit;
  wire        _slots_2_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_2_io_out_uop_ldst;
  wire [5:0]  _slots_2_io_out_uop_lrs1;
  wire [5:0]  _slots_2_io_out_uop_lrs2;
  wire [5:0]  _slots_2_io_out_uop_lrs3;
  wire        _slots_2_io_out_uop_ldst_val;
  wire [1:0]  _slots_2_io_out_uop_dst_rtype;
  wire [1:0]  _slots_2_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_2_io_out_uop_lrs2_rtype;
  wire        _slots_2_io_out_uop_frs3_en;
  wire        _slots_2_io_out_uop_fp_val;
  wire        _slots_2_io_out_uop_fp_single;
  wire        _slots_2_io_out_uop_xcpt_pf_if;
  wire        _slots_2_io_out_uop_xcpt_ae_if;
  wire        _slots_2_io_out_uop_xcpt_ma_if;
  wire        _slots_2_io_out_uop_bp_debug_if;
  wire        _slots_2_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_2_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_2_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_2_io_uop_uopc;
  wire [31:0] _slots_2_io_uop_inst;
  wire [31:0] _slots_2_io_uop_debug_inst;
  wire        _slots_2_io_uop_is_rvc;
  wire [39:0] _slots_2_io_uop_debug_pc;
  wire [2:0]  _slots_2_io_uop_iq_type;
  wire [9:0]  _slots_2_io_uop_fu_code;
  wire [1:0]  _slots_2_io_uop_iw_state;
  wire        _slots_2_io_uop_iw_p1_poisoned;
  wire        _slots_2_io_uop_iw_p2_poisoned;
  wire        _slots_2_io_uop_is_br;
  wire        _slots_2_io_uop_is_jalr;
  wire        _slots_2_io_uop_is_jal;
  wire        _slots_2_io_uop_is_sfb;
  wire [19:0] _slots_2_io_uop_br_mask;
  wire [4:0]  _slots_2_io_uop_br_tag;
  wire [5:0]  _slots_2_io_uop_ftq_idx;
  wire        _slots_2_io_uop_edge_inst;
  wire [5:0]  _slots_2_io_uop_pc_lob;
  wire        _slots_2_io_uop_taken;
  wire [19:0] _slots_2_io_uop_imm_packed;
  wire [11:0] _slots_2_io_uop_csr_addr;
  wire [6:0]  _slots_2_io_uop_rob_idx;
  wire [4:0]  _slots_2_io_uop_ldq_idx;
  wire [4:0]  _slots_2_io_uop_stq_idx;
  wire [1:0]  _slots_2_io_uop_rxq_idx;
  wire [6:0]  _slots_2_io_uop_pdst;
  wire [6:0]  _slots_2_io_uop_prs1;
  wire [6:0]  _slots_2_io_uop_prs2;
  wire [6:0]  _slots_2_io_uop_prs3;
  wire [5:0]  _slots_2_io_uop_ppred;
  wire        _slots_2_io_uop_prs1_busy;
  wire        _slots_2_io_uop_prs2_busy;
  wire        _slots_2_io_uop_prs3_busy;
  wire        _slots_2_io_uop_ppred_busy;
  wire [6:0]  _slots_2_io_uop_stale_pdst;
  wire        _slots_2_io_uop_exception;
  wire [63:0] _slots_2_io_uop_exc_cause;
  wire        _slots_2_io_uop_bypassable;
  wire [4:0]  _slots_2_io_uop_mem_cmd;
  wire [1:0]  _slots_2_io_uop_mem_size;
  wire        _slots_2_io_uop_mem_signed;
  wire        _slots_2_io_uop_is_fence;
  wire        _slots_2_io_uop_is_fencei;
  wire        _slots_2_io_uop_is_amo;
  wire        _slots_2_io_uop_uses_ldq;
  wire        _slots_2_io_uop_uses_stq;
  wire        _slots_2_io_uop_is_sys_pc2epc;
  wire        _slots_2_io_uop_is_unique;
  wire        _slots_2_io_uop_flush_on_commit;
  wire        _slots_2_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_2_io_uop_ldst;
  wire [5:0]  _slots_2_io_uop_lrs1;
  wire [5:0]  _slots_2_io_uop_lrs2;
  wire [5:0]  _slots_2_io_uop_lrs3;
  wire        _slots_2_io_uop_ldst_val;
  wire [1:0]  _slots_2_io_uop_dst_rtype;
  wire [1:0]  _slots_2_io_uop_lrs1_rtype;
  wire [1:0]  _slots_2_io_uop_lrs2_rtype;
  wire        _slots_2_io_uop_frs3_en;
  wire        _slots_2_io_uop_fp_val;
  wire        _slots_2_io_uop_fp_single;
  wire        _slots_2_io_uop_xcpt_pf_if;
  wire        _slots_2_io_uop_xcpt_ae_if;
  wire        _slots_2_io_uop_xcpt_ma_if;
  wire        _slots_2_io_uop_bp_debug_if;
  wire        _slots_2_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_2_io_uop_debug_fsrc;
  wire [1:0]  _slots_2_io_uop_debug_tsrc;
  wire        _slots_1_io_valid;
  wire        _slots_1_io_will_be_valid;
  wire        _slots_1_io_request;
  wire [6:0]  _slots_1_io_out_uop_uopc;
  wire [31:0] _slots_1_io_out_uop_inst;
  wire [31:0] _slots_1_io_out_uop_debug_inst;
  wire        _slots_1_io_out_uop_is_rvc;
  wire [39:0] _slots_1_io_out_uop_debug_pc;
  wire [2:0]  _slots_1_io_out_uop_iq_type;
  wire [9:0]  _slots_1_io_out_uop_fu_code;
  wire [1:0]  _slots_1_io_out_uop_iw_state;
  wire        _slots_1_io_out_uop_iw_p1_poisoned;
  wire        _slots_1_io_out_uop_iw_p2_poisoned;
  wire        _slots_1_io_out_uop_is_br;
  wire        _slots_1_io_out_uop_is_jalr;
  wire        _slots_1_io_out_uop_is_jal;
  wire        _slots_1_io_out_uop_is_sfb;
  wire [19:0] _slots_1_io_out_uop_br_mask;
  wire [4:0]  _slots_1_io_out_uop_br_tag;
  wire [5:0]  _slots_1_io_out_uop_ftq_idx;
  wire        _slots_1_io_out_uop_edge_inst;
  wire [5:0]  _slots_1_io_out_uop_pc_lob;
  wire        _slots_1_io_out_uop_taken;
  wire [19:0] _slots_1_io_out_uop_imm_packed;
  wire [11:0] _slots_1_io_out_uop_csr_addr;
  wire [6:0]  _slots_1_io_out_uop_rob_idx;
  wire [4:0]  _slots_1_io_out_uop_ldq_idx;
  wire [4:0]  _slots_1_io_out_uop_stq_idx;
  wire [1:0]  _slots_1_io_out_uop_rxq_idx;
  wire [6:0]  _slots_1_io_out_uop_pdst;
  wire [6:0]  _slots_1_io_out_uop_prs1;
  wire [6:0]  _slots_1_io_out_uop_prs2;
  wire [6:0]  _slots_1_io_out_uop_prs3;
  wire [5:0]  _slots_1_io_out_uop_ppred;
  wire        _slots_1_io_out_uop_prs1_busy;
  wire        _slots_1_io_out_uop_prs2_busy;
  wire        _slots_1_io_out_uop_prs3_busy;
  wire        _slots_1_io_out_uop_ppred_busy;
  wire [6:0]  _slots_1_io_out_uop_stale_pdst;
  wire        _slots_1_io_out_uop_exception;
  wire [63:0] _slots_1_io_out_uop_exc_cause;
  wire        _slots_1_io_out_uop_bypassable;
  wire [4:0]  _slots_1_io_out_uop_mem_cmd;
  wire [1:0]  _slots_1_io_out_uop_mem_size;
  wire        _slots_1_io_out_uop_mem_signed;
  wire        _slots_1_io_out_uop_is_fence;
  wire        _slots_1_io_out_uop_is_fencei;
  wire        _slots_1_io_out_uop_is_amo;
  wire        _slots_1_io_out_uop_uses_ldq;
  wire        _slots_1_io_out_uop_uses_stq;
  wire        _slots_1_io_out_uop_is_sys_pc2epc;
  wire        _slots_1_io_out_uop_is_unique;
  wire        _slots_1_io_out_uop_flush_on_commit;
  wire        _slots_1_io_out_uop_ldst_is_rs1;
  wire [5:0]  _slots_1_io_out_uop_ldst;
  wire [5:0]  _slots_1_io_out_uop_lrs1;
  wire [5:0]  _slots_1_io_out_uop_lrs2;
  wire [5:0]  _slots_1_io_out_uop_lrs3;
  wire        _slots_1_io_out_uop_ldst_val;
  wire [1:0]  _slots_1_io_out_uop_dst_rtype;
  wire [1:0]  _slots_1_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_1_io_out_uop_lrs2_rtype;
  wire        _slots_1_io_out_uop_frs3_en;
  wire        _slots_1_io_out_uop_fp_val;
  wire        _slots_1_io_out_uop_fp_single;
  wire        _slots_1_io_out_uop_xcpt_pf_if;
  wire        _slots_1_io_out_uop_xcpt_ae_if;
  wire        _slots_1_io_out_uop_xcpt_ma_if;
  wire        _slots_1_io_out_uop_bp_debug_if;
  wire        _slots_1_io_out_uop_bp_xcpt_if;
  wire [1:0]  _slots_1_io_out_uop_debug_fsrc;
  wire [1:0]  _slots_1_io_out_uop_debug_tsrc;
  wire [6:0]  _slots_1_io_uop_uopc;
  wire [31:0] _slots_1_io_uop_inst;
  wire [31:0] _slots_1_io_uop_debug_inst;
  wire        _slots_1_io_uop_is_rvc;
  wire [39:0] _slots_1_io_uop_debug_pc;
  wire [2:0]  _slots_1_io_uop_iq_type;
  wire [9:0]  _slots_1_io_uop_fu_code;
  wire [1:0]  _slots_1_io_uop_iw_state;
  wire        _slots_1_io_uop_iw_p1_poisoned;
  wire        _slots_1_io_uop_iw_p2_poisoned;
  wire        _slots_1_io_uop_is_br;
  wire        _slots_1_io_uop_is_jalr;
  wire        _slots_1_io_uop_is_jal;
  wire        _slots_1_io_uop_is_sfb;
  wire [19:0] _slots_1_io_uop_br_mask;
  wire [4:0]  _slots_1_io_uop_br_tag;
  wire [5:0]  _slots_1_io_uop_ftq_idx;
  wire        _slots_1_io_uop_edge_inst;
  wire [5:0]  _slots_1_io_uop_pc_lob;
  wire        _slots_1_io_uop_taken;
  wire [19:0] _slots_1_io_uop_imm_packed;
  wire [11:0] _slots_1_io_uop_csr_addr;
  wire [6:0]  _slots_1_io_uop_rob_idx;
  wire [4:0]  _slots_1_io_uop_ldq_idx;
  wire [4:0]  _slots_1_io_uop_stq_idx;
  wire [1:0]  _slots_1_io_uop_rxq_idx;
  wire [6:0]  _slots_1_io_uop_pdst;
  wire [6:0]  _slots_1_io_uop_prs1;
  wire [6:0]  _slots_1_io_uop_prs2;
  wire [6:0]  _slots_1_io_uop_prs3;
  wire [5:0]  _slots_1_io_uop_ppred;
  wire        _slots_1_io_uop_prs1_busy;
  wire        _slots_1_io_uop_prs2_busy;
  wire        _slots_1_io_uop_prs3_busy;
  wire        _slots_1_io_uop_ppred_busy;
  wire [6:0]  _slots_1_io_uop_stale_pdst;
  wire        _slots_1_io_uop_exception;
  wire [63:0] _slots_1_io_uop_exc_cause;
  wire        _slots_1_io_uop_bypassable;
  wire [4:0]  _slots_1_io_uop_mem_cmd;
  wire [1:0]  _slots_1_io_uop_mem_size;
  wire        _slots_1_io_uop_mem_signed;
  wire        _slots_1_io_uop_is_fence;
  wire        _slots_1_io_uop_is_fencei;
  wire        _slots_1_io_uop_is_amo;
  wire        _slots_1_io_uop_uses_ldq;
  wire        _slots_1_io_uop_uses_stq;
  wire        _slots_1_io_uop_is_sys_pc2epc;
  wire        _slots_1_io_uop_is_unique;
  wire        _slots_1_io_uop_flush_on_commit;
  wire        _slots_1_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_1_io_uop_ldst;
  wire [5:0]  _slots_1_io_uop_lrs1;
  wire [5:0]  _slots_1_io_uop_lrs2;
  wire [5:0]  _slots_1_io_uop_lrs3;
  wire        _slots_1_io_uop_ldst_val;
  wire [1:0]  _slots_1_io_uop_dst_rtype;
  wire [1:0]  _slots_1_io_uop_lrs1_rtype;
  wire [1:0]  _slots_1_io_uop_lrs2_rtype;
  wire        _slots_1_io_uop_frs3_en;
  wire        _slots_1_io_uop_fp_val;
  wire        _slots_1_io_uop_fp_single;
  wire        _slots_1_io_uop_xcpt_pf_if;
  wire        _slots_1_io_uop_xcpt_ae_if;
  wire        _slots_1_io_uop_xcpt_ma_if;
  wire        _slots_1_io_uop_bp_debug_if;
  wire        _slots_1_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_1_io_uop_debug_fsrc;
  wire [1:0]  _slots_1_io_uop_debug_tsrc;
  wire        _slots_0_io_valid;
  wire        _slots_0_io_will_be_valid;
  wire        _slots_0_io_request;
  wire [6:0]  _slots_0_io_uop_uopc;
  wire [31:0] _slots_0_io_uop_inst;
  wire [31:0] _slots_0_io_uop_debug_inst;
  wire        _slots_0_io_uop_is_rvc;
  wire [39:0] _slots_0_io_uop_debug_pc;
  wire [2:0]  _slots_0_io_uop_iq_type;
  wire [9:0]  _slots_0_io_uop_fu_code;
  wire [1:0]  _slots_0_io_uop_iw_state;
  wire        _slots_0_io_uop_iw_p1_poisoned;
  wire        _slots_0_io_uop_iw_p2_poisoned;
  wire        _slots_0_io_uop_is_br;
  wire        _slots_0_io_uop_is_jalr;
  wire        _slots_0_io_uop_is_jal;
  wire        _slots_0_io_uop_is_sfb;
  wire [19:0] _slots_0_io_uop_br_mask;
  wire [4:0]  _slots_0_io_uop_br_tag;
  wire [5:0]  _slots_0_io_uop_ftq_idx;
  wire        _slots_0_io_uop_edge_inst;
  wire [5:0]  _slots_0_io_uop_pc_lob;
  wire        _slots_0_io_uop_taken;
  wire [19:0] _slots_0_io_uop_imm_packed;
  wire [11:0] _slots_0_io_uop_csr_addr;
  wire [6:0]  _slots_0_io_uop_rob_idx;
  wire [4:0]  _slots_0_io_uop_ldq_idx;
  wire [4:0]  _slots_0_io_uop_stq_idx;
  wire [1:0]  _slots_0_io_uop_rxq_idx;
  wire [6:0]  _slots_0_io_uop_pdst;
  wire [6:0]  _slots_0_io_uop_prs1;
  wire [6:0]  _slots_0_io_uop_prs2;
  wire [6:0]  _slots_0_io_uop_prs3;
  wire [5:0]  _slots_0_io_uop_ppred;
  wire        _slots_0_io_uop_prs1_busy;
  wire        _slots_0_io_uop_prs2_busy;
  wire        _slots_0_io_uop_prs3_busy;
  wire        _slots_0_io_uop_ppred_busy;
  wire [6:0]  _slots_0_io_uop_stale_pdst;
  wire        _slots_0_io_uop_exception;
  wire [63:0] _slots_0_io_uop_exc_cause;
  wire        _slots_0_io_uop_bypassable;
  wire [4:0]  _slots_0_io_uop_mem_cmd;
  wire [1:0]  _slots_0_io_uop_mem_size;
  wire        _slots_0_io_uop_mem_signed;
  wire        _slots_0_io_uop_is_fence;
  wire        _slots_0_io_uop_is_fencei;
  wire        _slots_0_io_uop_is_amo;
  wire        _slots_0_io_uop_uses_ldq;
  wire        _slots_0_io_uop_uses_stq;
  wire        _slots_0_io_uop_is_sys_pc2epc;
  wire        _slots_0_io_uop_is_unique;
  wire        _slots_0_io_uop_flush_on_commit;
  wire        _slots_0_io_uop_ldst_is_rs1;
  wire [5:0]  _slots_0_io_uop_ldst;
  wire [5:0]  _slots_0_io_uop_lrs1;
  wire [5:0]  _slots_0_io_uop_lrs2;
  wire [5:0]  _slots_0_io_uop_lrs3;
  wire        _slots_0_io_uop_ldst_val;
  wire [1:0]  _slots_0_io_uop_dst_rtype;
  wire [1:0]  _slots_0_io_uop_lrs1_rtype;
  wire [1:0]  _slots_0_io_uop_lrs2_rtype;
  wire        _slots_0_io_uop_frs3_en;
  wire        _slots_0_io_uop_fp_val;
  wire        _slots_0_io_uop_fp_single;
  wire        _slots_0_io_uop_xcpt_pf_if;
  wire        _slots_0_io_uop_xcpt_ae_if;
  wire        _slots_0_io_uop_xcpt_ma_if;
  wire        _slots_0_io_uop_bp_debug_if;
  wire        _slots_0_io_uop_bp_xcpt_if;
  wire [1:0]  _slots_0_io_uop_debug_fsrc;
  wire [1:0]  _slots_0_io_uop_debug_tsrc;
  wire        _GEN = io_dis_uops_0_bits_uopc == 7'h2;
  wire        _GEN_0 = _GEN & ~(|io_dis_uops_0_bits_lrs2_rtype) | io_dis_uops_0_bits_uopc == 7'h43;
  wire [1:0]  _GEN_1 = _GEN_0 ? 2'h2 : 2'h1;
  wire        _GEN_2 = _GEN_0 | ~(_GEN & (|io_dis_uops_0_bits_lrs2_rtype));
  wire [1:0]  _GEN_3 = _GEN_2 ? io_dis_uops_0_bits_lrs2_rtype : 2'h2;
  wire        _GEN_4 = _GEN_2 & io_dis_uops_0_bits_prs2_busy;
  wire        _GEN_5 = io_dis_uops_1_bits_uopc == 7'h2;
  wire        _GEN_6 = _GEN_5 & ~(|io_dis_uops_1_bits_lrs2_rtype) | io_dis_uops_1_bits_uopc == 7'h43;
  wire [1:0]  _GEN_7 = _GEN_6 ? 2'h2 : 2'h1;
  wire        _GEN_8 = _GEN_6 | ~(_GEN_5 & (|io_dis_uops_1_bits_lrs2_rtype));
  wire [1:0]  _GEN_9 = _GEN_8 ? io_dis_uops_1_bits_lrs2_rtype : 2'h2;
  wire        _GEN_10 = _GEN_8 & io_dis_uops_1_bits_prs2_busy;
  wire        _GEN_11 = io_dis_uops_2_bits_uopc == 7'h2;
  wire        _GEN_12 = _GEN_11 & ~(|io_dis_uops_2_bits_lrs2_rtype) | io_dis_uops_2_bits_uopc == 7'h43;
  wire        _GEN_13 = _GEN_12 | ~(_GEN_11 & (|io_dis_uops_2_bits_lrs2_rtype));
  wire [1:0]  _GEN_14 = _GEN_13 ? io_dis_uops_2_bits_lrs2_rtype : 2'h2;
  wire        _GEN_15 = _GEN_13 & io_dis_uops_2_bits_prs2_busy;
  wire        _GEN_16 = io_dis_uops_3_bits_uopc == 7'h2;
  wire        _GEN_17 = _GEN_16 & ~(|io_dis_uops_3_bits_lrs2_rtype) | io_dis_uops_3_bits_uopc == 7'h43;
  wire        _GEN_18 = _GEN_17 | ~(_GEN_16 & (|io_dis_uops_3_bits_lrs2_rtype));
  wire [5:0]  count = {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, _slots_0_io_valid} + {1'h0, _slots_1_io_valid}} + {1'h0, {1'h0, _slots_2_io_valid} + {1'h0, _slots_3_io_valid} + {1'h0, _slots_4_io_valid}}} + {1'h0, {1'h0, {1'h0, _slots_5_io_valid} + {1'h0, _slots_6_io_valid}} + {1'h0, {1'h0, _slots_7_io_valid} + {1'h0, _slots_8_io_valid} + {1'h0, _slots_9_io_valid}}}} + {1'h0, {1'h0, {1'h0, {1'h0, _slots_10_io_valid} + {1'h0, _slots_11_io_valid}} + {1'h0, {1'h0, _slots_12_io_valid} + {1'h0, _slots_13_io_valid} + {1'h0, _slots_14_io_valid}}} + {1'h0, {1'h0, {1'h0, _slots_15_io_valid} + {1'h0, _slots_16_io_valid}} + {1'h0, {1'h0, _slots_17_io_valid} + {1'h0, _slots_18_io_valid} + {1'h0, _slots_19_io_valid}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, _slots_20_io_valid} + {1'h0, _slots_21_io_valid}} + {1'h0, {1'h0, _slots_22_io_valid} + {1'h0, _slots_23_io_valid} + {1'h0, _slots_24_io_valid}}} + {1'h0, {1'h0, {1'h0, _slots_25_io_valid} + {1'h0, _slots_26_io_valid}} + {1'h0, {1'h0, _slots_27_io_valid} + {1'h0, _slots_28_io_valid} + {1'h0, _slots_29_io_valid}}}} + {1'h0, {1'h0, {1'h0, {1'h0, _slots_30_io_valid} + {1'h0, _slots_31_io_valid}} + {1'h0, {1'h0, _slots_32_io_valid} + {1'h0, _slots_33_io_valid} + {1'h0, _slots_34_io_valid}}} + {1'h0, {1'h0, {1'h0, _slots_35_io_valid} + {1'h0, _slots_36_io_valid}} + {1'h0, {1'h0, _slots_37_io_valid} + {1'h0, _slots_38_io_valid} + {1'h0, _slots_39_io_valid}}}}};
  `ifndef SYNTHESIS
    always @(posedge clock) begin
      if (~reset & {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, issue_slots_0_grant} + {1'h0, issue_slots_1_grant}} + {1'h0, {1'h0, issue_slots_2_grant} + {1'h0, issue_slots_3_grant} + {1'h0, issue_slots_4_grant}}} + {1'h0, {1'h0, {1'h0, issue_slots_5_grant} + {1'h0, issue_slots_6_grant}} + {1'h0, {1'h0, issue_slots_7_grant} + {1'h0, issue_slots_8_grant} + {1'h0, issue_slots_9_grant}}}} + {1'h0, {1'h0, {1'h0, {1'h0, issue_slots_10_grant} + {1'h0, issue_slots_11_grant}} + {1'h0, {1'h0, issue_slots_12_grant} + {1'h0, issue_slots_13_grant} + {1'h0, issue_slots_14_grant}}} + {1'h0, {1'h0, {1'h0, issue_slots_15_grant} + {1'h0, issue_slots_16_grant}} + {1'h0, {1'h0, issue_slots_17_grant} + {1'h0, issue_slots_18_grant} + {1'h0, issue_slots_19_grant}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, issue_slots_20_grant} + {1'h0, issue_slots_21_grant}} + {1'h0, {1'h0, issue_slots_22_grant} + {1'h0, issue_slots_23_grant} + {1'h0, issue_slots_24_grant}}} + {1'h0, {1'h0, {1'h0, issue_slots_25_grant} + {1'h0, issue_slots_26_grant}} + {1'h0, {1'h0, issue_slots_27_grant} + {1'h0, issue_slots_28_grant} + {1'h0, issue_slots_29_grant}}}} + {1'h0, {1'h0, {1'h0, {1'h0, issue_slots_30_grant} + {1'h0, issue_slots_31_grant}} + {1'h0, {1'h0, issue_slots_32_grant} + {1'h0, issue_slots_33_grant} + {1'h0, issue_slots_34_grant}}} + {1'h0, {1'h0, {1'h0, issue_slots_35_grant} + {1'h0, issue_slots_36_grant}} + {1'h0, {1'h0, issue_slots_37_grant} + {1'h0, issue_slots_38_grant} + {1'h0, issue_slots_39_grant}}}}} > 6'h4) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [issue] window giving out too many grants.\n    at issue-unit.scala:172 assert (PopCount(issue_slots.map(s => s.grant)) <= issueWidth.U, \"[issue] window giving out too many grants.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire [3:0]  next_1 = _slots_0_io_valid & ~_slots_1_io_valid ? 4'h1 : _slots_1_io_valid ? {3'h0, ~_slots_0_io_valid} : {2'h0, ~_slots_0_io_valid, 1'h0};
  assign _next_1_1to0 = next_1[1:0];
  assign next_2 = _next_1_1to0 == 2'h0 & ~_slots_2_io_valid ? 4'h1 : next_1[3] | _slots_2_io_valid ? next_1 : {next_1[2:0], 1'h0};
  assign next_3 = next_2 == 4'h0 & ~_slots_3_io_valid ? 4'h1 : next_2[3] | _slots_3_io_valid ? next_2 : {next_2[2:0], 1'h0};
  assign next_4 = next_3 == 4'h0 & ~_slots_4_io_valid ? 4'h1 : next_3[3] | _slots_4_io_valid ? next_3 : {next_3[2:0], 1'h0};
  assign next_5 = next_4 == 4'h0 & ~_slots_5_io_valid ? 4'h1 : next_4[3] | _slots_5_io_valid ? next_4 : {next_4[2:0], 1'h0};
  assign next_6 = next_5 == 4'h0 & ~_slots_6_io_valid ? 4'h1 : next_5[3] | _slots_6_io_valid ? next_5 : {next_5[2:0], 1'h0};
  assign next_7 = next_6 == 4'h0 & ~_slots_7_io_valid ? 4'h1 : next_6[3] | _slots_7_io_valid ? next_6 : {next_6[2:0], 1'h0};
  assign next_8 = next_7 == 4'h0 & ~_slots_8_io_valid ? 4'h1 : next_7[3] | _slots_8_io_valid ? next_7 : {next_7[2:0], 1'h0};
  assign next_9 = next_8 == 4'h0 & ~_slots_9_io_valid ? 4'h1 : next_8[3] | _slots_9_io_valid ? next_8 : {next_8[2:0], 1'h0};
  assign next_10 = next_9 == 4'h0 & ~_slots_10_io_valid ? 4'h1 : next_9[3] | _slots_10_io_valid ? next_9 : {next_9[2:0], 1'h0};
  assign next_11 = next_10 == 4'h0 & ~_slots_11_io_valid ? 4'h1 : next_10[3] | _slots_11_io_valid ? next_10 : {next_10[2:0], 1'h0};
  assign next_12 = next_11 == 4'h0 & ~_slots_12_io_valid ? 4'h1 : next_11[3] | _slots_12_io_valid ? next_11 : {next_11[2:0], 1'h0};
  assign next_13 = next_12 == 4'h0 & ~_slots_13_io_valid ? 4'h1 : next_12[3] | _slots_13_io_valid ? next_12 : {next_12[2:0], 1'h0};
  assign next_14 = next_13 == 4'h0 & ~_slots_14_io_valid ? 4'h1 : next_13[3] | _slots_14_io_valid ? next_13 : {next_13[2:0], 1'h0};
  assign next_15 = next_14 == 4'h0 & ~_slots_15_io_valid ? 4'h1 : next_14[3] | _slots_15_io_valid ? next_14 : {next_14[2:0], 1'h0};
  assign next_16 = next_15 == 4'h0 & ~_slots_16_io_valid ? 4'h1 : next_15[3] | _slots_16_io_valid ? next_15 : {next_15[2:0], 1'h0};
  assign next_17 = next_16 == 4'h0 & ~_slots_17_io_valid ? 4'h1 : next_16[3] | _slots_17_io_valid ? next_16 : {next_16[2:0], 1'h0};
  assign next_18 = next_17 == 4'h0 & ~_slots_18_io_valid ? 4'h1 : next_17[3] | _slots_18_io_valid ? next_17 : {next_17[2:0], 1'h0};
  assign next_19 = next_18 == 4'h0 & ~_slots_19_io_valid ? 4'h1 : next_18[3] | _slots_19_io_valid ? next_18 : {next_18[2:0], 1'h0};
  assign next_20 = next_19 == 4'h0 & ~_slots_20_io_valid ? 4'h1 : next_19[3] | _slots_20_io_valid ? next_19 : {next_19[2:0], 1'h0};
  assign next_21 = next_20 == 4'h0 & ~_slots_21_io_valid ? 4'h1 : next_20[3] | _slots_21_io_valid ? next_20 : {next_20[2:0], 1'h0};
  assign next_22 = next_21 == 4'h0 & ~_slots_22_io_valid ? 4'h1 : next_21[3] | _slots_22_io_valid ? next_21 : {next_21[2:0], 1'h0};
  assign next_23 = next_22 == 4'h0 & ~_slots_23_io_valid ? 4'h1 : next_22[3] | _slots_23_io_valid ? next_22 : {next_22[2:0], 1'h0};
  assign next_24 = next_23 == 4'h0 & ~_slots_24_io_valid ? 4'h1 : next_23[3] | _slots_24_io_valid ? next_23 : {next_23[2:0], 1'h0};
  assign next_25 = next_24 == 4'h0 & ~_slots_25_io_valid ? 4'h1 : next_24[3] | _slots_25_io_valid ? next_24 : {next_24[2:0], 1'h0};
  assign next_26 = next_25 == 4'h0 & ~_slots_26_io_valid ? 4'h1 : next_25[3] | _slots_26_io_valid ? next_25 : {next_25[2:0], 1'h0};
  assign next_27 = next_26 == 4'h0 & ~_slots_27_io_valid ? 4'h1 : next_26[3] | _slots_27_io_valid ? next_26 : {next_26[2:0], 1'h0};
  assign next_28 = next_27 == 4'h0 & ~_slots_28_io_valid ? 4'h1 : next_27[3] | _slots_28_io_valid ? next_27 : {next_27[2:0], 1'h0};
  assign next_29 = next_28 == 4'h0 & ~_slots_29_io_valid ? 4'h1 : next_28[3] | _slots_29_io_valid ? next_28 : {next_28[2:0], 1'h0};
  assign next_30 = next_29 == 4'h0 & ~_slots_30_io_valid ? 4'h1 : next_29[3] | _slots_30_io_valid ? next_29 : {next_29[2:0], 1'h0};
  assign next_31 = next_30 == 4'h0 & ~_slots_31_io_valid ? 4'h1 : next_30[3] | _slots_31_io_valid ? next_30 : {next_30[2:0], 1'h0};
  assign next_32 = next_31 == 4'h0 & ~_slots_32_io_valid ? 4'h1 : next_31[3] | _slots_32_io_valid ? next_31 : {next_31[2:0], 1'h0};
  assign next_33 = next_32 == 4'h0 & ~_slots_33_io_valid ? 4'h1 : next_32[3] | _slots_33_io_valid ? next_32 : {next_32[2:0], 1'h0};
  assign next_34 = next_33 == 4'h0 & ~_slots_34_io_valid ? 4'h1 : next_33[3] | _slots_34_io_valid ? next_33 : {next_33[2:0], 1'h0};
  assign next_35 = next_34 == 4'h0 & ~_slots_35_io_valid ? 4'h1 : next_34[3] | _slots_35_io_valid ? next_34 : {next_34[2:0], 1'h0};
  assign next_36 = next_35 == 4'h0 & ~_slots_36_io_valid ? 4'h1 : next_35[3] | _slots_36_io_valid ? next_35 : {next_35[2:0], 1'h0};
  assign next_37 = next_36 == 4'h0 & ~_slots_37_io_valid ? 4'h1 : next_36[3] | _slots_37_io_valid ? next_36 : {next_36[2:0], 1'h0};
  assign next_38 = next_37 == 4'h0 & ~_slots_38_io_valid ? 4'h1 : next_37[3] | _slots_38_io_valid ? next_37 : {next_37[2:0], 1'h0};
  wire [3:0]  next_39 = next_38 == 4'h0 & ~_slots_39_io_valid ? 4'h1 : next_38[3] | _slots_39_io_valid ? next_38 : {next_38[2:0], 1'h0};
  wire [3:0]  next_40 = next_39 == 4'h0 & ~io_dis_uops_0_valid ? 4'h1 : next_39[3] | io_dis_uops_0_valid ? next_39 : {next_39[2:0], 1'h0};
  wire [3:0]  next_41 = next_40 == 4'h0 & ~io_dis_uops_1_valid ? 4'h1 : next_40[3] | io_dis_uops_1_valid ? next_40 : {next_40[2:0], 1'h0};
  wire        will_be_valid_40 = io_dis_uops_0_valid & ~io_dis_uops_0_bits_exception & ~io_dis_uops_0_bits_is_fence & ~io_dis_uops_0_bits_is_fencei;
  wire        will_be_valid_41 = io_dis_uops_1_valid & ~io_dis_uops_1_bits_exception & ~io_dis_uops_1_bits_is_fence & ~io_dis_uops_1_bits_is_fencei;
  wire        will_be_valid_42 = io_dis_uops_2_valid & ~io_dis_uops_2_bits_exception & ~io_dis_uops_2_bits_is_fence & ~io_dis_uops_2_bits_is_fencei;
  wire        _GEN_19 = _next_1_1to0 == 2'h2;
  wire        _GEN_20 = next_2 == 4'h4;
  wire        _GEN_21 = next_3 == 4'h8;
  wire        issue_slots_0_in_uop_valid = _GEN_21 ? _slots_4_io_will_be_valid : _GEN_20 ? _slots_3_io_will_be_valid : _GEN_19 ? _slots_2_io_will_be_valid : ~_slots_0_io_valid & _slots_1_io_will_be_valid;
  wire        _GEN_22 = next_2 == 4'h2;
  wire        _GEN_23 = next_3 == 4'h4;
  wire        _GEN_24 = next_4 == 4'h8;
  wire        issue_slots_1_in_uop_valid = _GEN_24 ? _slots_5_io_will_be_valid : _GEN_23 ? _slots_4_io_will_be_valid : _GEN_22 ? _slots_3_io_will_be_valid : _next_1_1to0 == 2'h1 & _slots_2_io_will_be_valid;
  wire        _GEN_25 = next_3 == 4'h2;
  wire        _GEN_26 = next_4 == 4'h4;
  wire        _GEN_27 = next_5 == 4'h8;
  wire        issue_slots_2_in_uop_valid = _GEN_27 ? _slots_6_io_will_be_valid : _GEN_26 ? _slots_5_io_will_be_valid : _GEN_25 ? _slots_4_io_will_be_valid : next_2 == 4'h1 & _slots_3_io_will_be_valid;
  wire        _GEN_28 = next_4 == 4'h2;
  wire        _GEN_29 = next_5 == 4'h4;
  wire        _GEN_30 = next_6 == 4'h8;
  wire        issue_slots_3_in_uop_valid = _GEN_30 ? _slots_7_io_will_be_valid : _GEN_29 ? _slots_6_io_will_be_valid : _GEN_28 ? _slots_5_io_will_be_valid : next_3 == 4'h1 & _slots_4_io_will_be_valid;
  wire        _GEN_31 = next_5 == 4'h2;
  wire        _GEN_32 = next_6 == 4'h4;
  wire        _GEN_33 = next_7 == 4'h8;
  wire        issue_slots_4_in_uop_valid = _GEN_33 ? _slots_8_io_will_be_valid : _GEN_32 ? _slots_7_io_will_be_valid : _GEN_31 ? _slots_6_io_will_be_valid : next_4 == 4'h1 & _slots_5_io_will_be_valid;
  wire        _GEN_34 = next_6 == 4'h2;
  wire        _GEN_35 = next_7 == 4'h4;
  wire        _GEN_36 = next_8 == 4'h8;
  wire        issue_slots_5_in_uop_valid = _GEN_36 ? _slots_9_io_will_be_valid : _GEN_35 ? _slots_8_io_will_be_valid : _GEN_34 ? _slots_7_io_will_be_valid : next_5 == 4'h1 & _slots_6_io_will_be_valid;
  wire        _GEN_37 = next_7 == 4'h2;
  wire        _GEN_38 = next_8 == 4'h4;
  wire        _GEN_39 = next_9 == 4'h8;
  wire        issue_slots_6_in_uop_valid = _GEN_39 ? _slots_10_io_will_be_valid : _GEN_38 ? _slots_9_io_will_be_valid : _GEN_37 ? _slots_8_io_will_be_valid : next_6 == 4'h1 & _slots_7_io_will_be_valid;
  wire        _GEN_40 = next_8 == 4'h2;
  wire        _GEN_41 = next_9 == 4'h4;
  wire        _GEN_42 = next_10 == 4'h8;
  wire        issue_slots_7_in_uop_valid = _GEN_42 ? _slots_11_io_will_be_valid : _GEN_41 ? _slots_10_io_will_be_valid : _GEN_40 ? _slots_9_io_will_be_valid : next_7 == 4'h1 & _slots_8_io_will_be_valid;
  wire        _GEN_43 = next_9 == 4'h2;
  wire        _GEN_44 = next_10 == 4'h4;
  wire        _GEN_45 = next_11 == 4'h8;
  wire        issue_slots_8_in_uop_valid = _GEN_45 ? _slots_12_io_will_be_valid : _GEN_44 ? _slots_11_io_will_be_valid : _GEN_43 ? _slots_10_io_will_be_valid : next_8 == 4'h1 & _slots_9_io_will_be_valid;
  wire        _GEN_46 = next_10 == 4'h2;
  wire        _GEN_47 = next_11 == 4'h4;
  wire        _GEN_48 = next_12 == 4'h8;
  wire        issue_slots_9_in_uop_valid = _GEN_48 ? _slots_13_io_will_be_valid : _GEN_47 ? _slots_12_io_will_be_valid : _GEN_46 ? _slots_11_io_will_be_valid : next_9 == 4'h1 & _slots_10_io_will_be_valid;
  wire        _GEN_49 = next_11 == 4'h2;
  wire        _GEN_50 = next_12 == 4'h4;
  wire        _GEN_51 = next_13 == 4'h8;
  wire        issue_slots_10_in_uop_valid = _GEN_51 ? _slots_14_io_will_be_valid : _GEN_50 ? _slots_13_io_will_be_valid : _GEN_49 ? _slots_12_io_will_be_valid : next_10 == 4'h1 & _slots_11_io_will_be_valid;
  wire        _GEN_52 = next_12 == 4'h2;
  wire        _GEN_53 = next_13 == 4'h4;
  wire        _GEN_54 = next_14 == 4'h8;
  wire        issue_slots_11_in_uop_valid = _GEN_54 ? _slots_15_io_will_be_valid : _GEN_53 ? _slots_14_io_will_be_valid : _GEN_52 ? _slots_13_io_will_be_valid : next_11 == 4'h1 & _slots_12_io_will_be_valid;
  wire        _GEN_55 = next_13 == 4'h2;
  wire        _GEN_56 = next_14 == 4'h4;
  wire        _GEN_57 = next_15 == 4'h8;
  wire        issue_slots_12_in_uop_valid = _GEN_57 ? _slots_16_io_will_be_valid : _GEN_56 ? _slots_15_io_will_be_valid : _GEN_55 ? _slots_14_io_will_be_valid : next_12 == 4'h1 & _slots_13_io_will_be_valid;
  wire        _GEN_58 = next_14 == 4'h2;
  wire        _GEN_59 = next_15 == 4'h4;
  wire        _GEN_60 = next_16 == 4'h8;
  wire        issue_slots_13_in_uop_valid = _GEN_60 ? _slots_17_io_will_be_valid : _GEN_59 ? _slots_16_io_will_be_valid : _GEN_58 ? _slots_15_io_will_be_valid : next_13 == 4'h1 & _slots_14_io_will_be_valid;
  wire        _GEN_61 = next_15 == 4'h2;
  wire        _GEN_62 = next_16 == 4'h4;
  wire        _GEN_63 = next_17 == 4'h8;
  wire        issue_slots_14_in_uop_valid = _GEN_63 ? _slots_18_io_will_be_valid : _GEN_62 ? _slots_17_io_will_be_valid : _GEN_61 ? _slots_16_io_will_be_valid : next_14 == 4'h1 & _slots_15_io_will_be_valid;
  wire        _GEN_64 = next_16 == 4'h2;
  wire        _GEN_65 = next_17 == 4'h4;
  wire        _GEN_66 = next_18 == 4'h8;
  wire        issue_slots_15_in_uop_valid = _GEN_66 ? _slots_19_io_will_be_valid : _GEN_65 ? _slots_18_io_will_be_valid : _GEN_64 ? _slots_17_io_will_be_valid : next_15 == 4'h1 & _slots_16_io_will_be_valid;
  wire        _GEN_67 = next_17 == 4'h2;
  wire        _GEN_68 = next_18 == 4'h4;
  wire        _GEN_69 = next_19 == 4'h8;
  wire        issue_slots_16_in_uop_valid = _GEN_69 ? _slots_20_io_will_be_valid : _GEN_68 ? _slots_19_io_will_be_valid : _GEN_67 ? _slots_18_io_will_be_valid : next_16 == 4'h1 & _slots_17_io_will_be_valid;
  wire        _GEN_70 = next_18 == 4'h2;
  wire        _GEN_71 = next_19 == 4'h4;
  wire        _GEN_72 = next_20 == 4'h8;
  wire        issue_slots_17_in_uop_valid = _GEN_72 ? _slots_21_io_will_be_valid : _GEN_71 ? _slots_20_io_will_be_valid : _GEN_70 ? _slots_19_io_will_be_valid : next_17 == 4'h1 & _slots_18_io_will_be_valid;
  wire        _GEN_73 = next_19 == 4'h2;
  wire        _GEN_74 = next_20 == 4'h4;
  wire        _GEN_75 = next_21 == 4'h8;
  wire        issue_slots_18_in_uop_valid = _GEN_75 ? _slots_22_io_will_be_valid : _GEN_74 ? _slots_21_io_will_be_valid : _GEN_73 ? _slots_20_io_will_be_valid : next_18 == 4'h1 & _slots_19_io_will_be_valid;
  wire        _GEN_76 = next_20 == 4'h2;
  wire        _GEN_77 = next_21 == 4'h4;
  wire        _GEN_78 = next_22 == 4'h8;
  wire        issue_slots_19_in_uop_valid = _GEN_78 ? _slots_23_io_will_be_valid : _GEN_77 ? _slots_22_io_will_be_valid : _GEN_76 ? _slots_21_io_will_be_valid : next_19 == 4'h1 & _slots_20_io_will_be_valid;
  wire        _GEN_79 = next_21 == 4'h2;
  wire        _GEN_80 = next_22 == 4'h4;
  wire        _GEN_81 = next_23 == 4'h8;
  wire        issue_slots_20_in_uop_valid = _GEN_81 ? _slots_24_io_will_be_valid : _GEN_80 ? _slots_23_io_will_be_valid : _GEN_79 ? _slots_22_io_will_be_valid : next_20 == 4'h1 & _slots_21_io_will_be_valid;
  wire        _GEN_82 = next_22 == 4'h2;
  wire        _GEN_83 = next_23 == 4'h4;
  wire        _GEN_84 = next_24 == 4'h8;
  wire        issue_slots_21_in_uop_valid = _GEN_84 ? _slots_25_io_will_be_valid : _GEN_83 ? _slots_24_io_will_be_valid : _GEN_82 ? _slots_23_io_will_be_valid : next_21 == 4'h1 & _slots_22_io_will_be_valid;
  wire        _GEN_85 = next_23 == 4'h2;
  wire        _GEN_86 = next_24 == 4'h4;
  wire        _GEN_87 = next_25 == 4'h8;
  wire        issue_slots_22_in_uop_valid = _GEN_87 ? _slots_26_io_will_be_valid : _GEN_86 ? _slots_25_io_will_be_valid : _GEN_85 ? _slots_24_io_will_be_valid : next_22 == 4'h1 & _slots_23_io_will_be_valid;
  wire        _GEN_88 = next_24 == 4'h2;
  wire        _GEN_89 = next_25 == 4'h4;
  wire        _GEN_90 = next_26 == 4'h8;
  wire        issue_slots_23_in_uop_valid = _GEN_90 ? _slots_27_io_will_be_valid : _GEN_89 ? _slots_26_io_will_be_valid : _GEN_88 ? _slots_25_io_will_be_valid : next_23 == 4'h1 & _slots_24_io_will_be_valid;
  wire        _GEN_91 = next_25 == 4'h2;
  wire        _GEN_92 = next_26 == 4'h4;
  wire        _GEN_93 = next_27 == 4'h8;
  wire        issue_slots_24_in_uop_valid = _GEN_93 ? _slots_28_io_will_be_valid : _GEN_92 ? _slots_27_io_will_be_valid : _GEN_91 ? _slots_26_io_will_be_valid : next_24 == 4'h1 & _slots_25_io_will_be_valid;
  wire        _GEN_94 = next_26 == 4'h2;
  wire        _GEN_95 = next_27 == 4'h4;
  wire        _GEN_96 = next_28 == 4'h8;
  wire        issue_slots_25_in_uop_valid = _GEN_96 ? _slots_29_io_will_be_valid : _GEN_95 ? _slots_28_io_will_be_valid : _GEN_94 ? _slots_27_io_will_be_valid : next_25 == 4'h1 & _slots_26_io_will_be_valid;
  wire        _GEN_97 = next_27 == 4'h2;
  wire        _GEN_98 = next_28 == 4'h4;
  wire        _GEN_99 = next_29 == 4'h8;
  wire        issue_slots_26_in_uop_valid = _GEN_99 ? _slots_30_io_will_be_valid : _GEN_98 ? _slots_29_io_will_be_valid : _GEN_97 ? _slots_28_io_will_be_valid : next_26 == 4'h1 & _slots_27_io_will_be_valid;
  wire        _GEN_100 = next_28 == 4'h2;
  wire        _GEN_101 = next_29 == 4'h4;
  wire        _GEN_102 = next_30 == 4'h8;
  wire        issue_slots_27_in_uop_valid = _GEN_102 ? _slots_31_io_will_be_valid : _GEN_101 ? _slots_30_io_will_be_valid : _GEN_100 ? _slots_29_io_will_be_valid : next_27 == 4'h1 & _slots_28_io_will_be_valid;
  wire        _GEN_103 = next_29 == 4'h2;
  wire        _GEN_104 = next_30 == 4'h4;
  wire        _GEN_105 = next_31 == 4'h8;
  wire        issue_slots_28_in_uop_valid = _GEN_105 ? _slots_32_io_will_be_valid : _GEN_104 ? _slots_31_io_will_be_valid : _GEN_103 ? _slots_30_io_will_be_valid : next_28 == 4'h1 & _slots_29_io_will_be_valid;
  wire        _GEN_106 = next_30 == 4'h2;
  wire        _GEN_107 = next_31 == 4'h4;
  wire        _GEN_108 = next_32 == 4'h8;
  wire        issue_slots_29_in_uop_valid = _GEN_108 ? _slots_33_io_will_be_valid : _GEN_107 ? _slots_32_io_will_be_valid : _GEN_106 ? _slots_31_io_will_be_valid : next_29 == 4'h1 & _slots_30_io_will_be_valid;
  wire        _GEN_109 = next_31 == 4'h2;
  wire        _GEN_110 = next_32 == 4'h4;
  wire        _GEN_111 = next_33 == 4'h8;
  wire        issue_slots_30_in_uop_valid = _GEN_111 ? _slots_34_io_will_be_valid : _GEN_110 ? _slots_33_io_will_be_valid : _GEN_109 ? _slots_32_io_will_be_valid : next_30 == 4'h1 & _slots_31_io_will_be_valid;
  wire        _GEN_112 = next_32 == 4'h2;
  wire        _GEN_113 = next_33 == 4'h4;
  wire        _GEN_114 = next_34 == 4'h8;
  wire        issue_slots_31_in_uop_valid = _GEN_114 ? _slots_35_io_will_be_valid : _GEN_113 ? _slots_34_io_will_be_valid : _GEN_112 ? _slots_33_io_will_be_valid : next_31 == 4'h1 & _slots_32_io_will_be_valid;
  wire        _GEN_115 = next_33 == 4'h2;
  wire        _GEN_116 = next_34 == 4'h4;
  wire        _GEN_117 = next_35 == 4'h8;
  wire        issue_slots_32_in_uop_valid = _GEN_117 ? _slots_36_io_will_be_valid : _GEN_116 ? _slots_35_io_will_be_valid : _GEN_115 ? _slots_34_io_will_be_valid : next_32 == 4'h1 & _slots_33_io_will_be_valid;
  wire        _GEN_118 = next_34 == 4'h2;
  wire        _GEN_119 = next_35 == 4'h4;
  wire        _GEN_120 = next_36 == 4'h8;
  wire        issue_slots_33_in_uop_valid = _GEN_120 ? _slots_37_io_will_be_valid : _GEN_119 ? _slots_36_io_will_be_valid : _GEN_118 ? _slots_35_io_will_be_valid : next_33 == 4'h1 & _slots_34_io_will_be_valid;
  wire        _GEN_121 = next_35 == 4'h2;
  wire        _GEN_122 = next_36 == 4'h4;
  wire        _GEN_123 = next_37 == 4'h8;
  wire        issue_slots_34_in_uop_valid = _GEN_123 ? _slots_38_io_will_be_valid : _GEN_122 ? _slots_37_io_will_be_valid : _GEN_121 ? _slots_36_io_will_be_valid : next_34 == 4'h1 & _slots_35_io_will_be_valid;
  wire        _GEN_124 = next_36 == 4'h2;
  wire        _GEN_125 = next_37 == 4'h4;
  wire        _GEN_126 = next_38 == 4'h8;
  wire        issue_slots_35_in_uop_valid = _GEN_126 ? _slots_39_io_will_be_valid : _GEN_125 ? _slots_38_io_will_be_valid : _GEN_124 ? _slots_37_io_will_be_valid : next_35 == 4'h1 & _slots_36_io_will_be_valid;
  wire        _GEN_127 = next_37 == 4'h2;
  wire        _GEN_128 = next_38 == 4'h4;
  wire        _GEN_129 = next_39 == 4'h8;
  wire        issue_slots_36_in_uop_valid = _GEN_129 ? will_be_valid_40 : _GEN_128 ? _slots_39_io_will_be_valid : _GEN_127 ? _slots_38_io_will_be_valid : next_36 == 4'h1 & _slots_37_io_will_be_valid;
  wire        _GEN_130 = next_38 == 4'h2;
  wire        _GEN_131 = next_39 == 4'h4;
  wire        _GEN_132 = next_40 == 4'h8;
  wire        issue_slots_37_in_uop_valid = _GEN_132 ? will_be_valid_41 : _GEN_131 ? will_be_valid_40 : _GEN_130 ? _slots_39_io_will_be_valid : next_37 == 4'h1 & _slots_38_io_will_be_valid;
  wire        _GEN_133 = _GEN_132 | _GEN_131;
  wire        _GEN_134 = next_39 == 4'h2;
  wire        _GEN_135 = next_40 == 4'h4;
  wire        _GEN_136 = next_41 == 4'h8;
  wire        issue_slots_38_in_uop_valid = _GEN_136 ? will_be_valid_42 : _GEN_135 ? will_be_valid_41 : _GEN_134 ? will_be_valid_40 : next_38 == 4'h1 & _slots_39_io_will_be_valid;
  wire        _GEN_137 = _GEN_136 | _GEN_135 | _GEN_134;
  wire        _GEN_138 = next_40 == 4'h2;
  wire        _GEN_139 = next_41 == 4'h4;
  wire        _GEN_140 = (next_41 == 4'h0 & ~io_dis_uops_2_valid ? 4'h1 : next_41[3] | io_dis_uops_2_valid ? next_41 : {next_41[2:0], 1'h0}) == 4'h8;
  wire        issue_slots_39_in_uop_valid = _GEN_140 ? io_dis_uops_3_valid & ~io_dis_uops_3_bits_exception & ~io_dis_uops_3_bits_is_fence & ~io_dis_uops_3_bits_is_fencei : _GEN_139 ? will_be_valid_42 : _GEN_138 ? will_be_valid_41 : next_39 == 4'h1 & will_be_valid_40;
  reg         io_dis_uops_0_ready_REG;
  reg         io_dis_uops_1_ready_REG;
  reg         io_dis_uops_2_ready_REG;
  reg         io_dis_uops_3_ready_REG;
  wire        _GEN_141 = _slots_0_io_request & (|(_slots_0_io_uop_fu_code & io_fu_types_0));
  wire [1:0]  _GEN_142 = {_slots_0_io_uop_fu_code[5], _slots_0_io_uop_fu_code[0]};
  wire        _GEN_143 = _slots_0_io_request & ~_GEN_141 & (|_GEN_142);
  wire        _GEN_144 = _slots_0_io_request & (|_GEN_142) | _GEN_141;
  wire [9:0]  _can_allocate_T_2 = _slots_0_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_145 = _slots_0_io_request & ~_GEN_144 & (|_can_allocate_T_2);
  wire        _GEN_146 = _slots_0_io_request & ~(_slots_0_io_request & (|_can_allocate_T_2) | _GEN_144) & (|(_slots_0_io_uop_fu_code & io_fu_types_3));
  assign issue_slots_0_grant = _GEN_146 | _GEN_145 | _GEN_143 | _GEN_141;
  wire        _GEN_147 = _slots_1_io_request & (|(_slots_1_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_148 = _GEN_147 & ~_GEN_141;
  wire        _GEN_149 = _GEN_147 | _GEN_141;
  wire [1:0]  _GEN_150 = {_slots_1_io_uop_fu_code[5], _slots_1_io_uop_fu_code[0]};
  wire        _GEN_151 = _slots_1_io_request & ~_GEN_148 & (|_GEN_150);
  wire        _GEN_152 = _GEN_151 & ~_GEN_143;
  wire        _GEN_153 = _GEN_151 | _GEN_143;
  wire        _GEN_154 = _slots_1_io_request & (|_GEN_150) & ~_GEN_143 | _GEN_148;
  wire [9:0]  _can_allocate_T_6 = _slots_1_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_155 = _slots_1_io_request & ~_GEN_154 & (|_can_allocate_T_6);
  wire        _GEN_156 = _GEN_155 & ~_GEN_145;
  wire        _GEN_157 = _GEN_155 | _GEN_145;
  wire        _GEN_158 = _slots_1_io_request & ~(_slots_1_io_request & (|_can_allocate_T_6) & ~_GEN_145 | _GEN_154) & (|(_slots_1_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_159 = _GEN_158 & ~_GEN_146;
  assign issue_slots_1_grant = _GEN_159 | _GEN_156 | _GEN_152 | _GEN_148;
  wire        _GEN_160 = _GEN_158 | _GEN_146;
  wire        _GEN_161 = _slots_2_io_request & (|(_slots_2_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_162 = _GEN_161 & ~_GEN_149;
  wire        _GEN_163 = _GEN_161 | _GEN_149;
  wire [1:0]  _GEN_164 = {_slots_2_io_uop_fu_code[5], _slots_2_io_uop_fu_code[0]};
  wire        _GEN_165 = _slots_2_io_request & ~_GEN_162 & (|_GEN_164);
  wire        _GEN_166 = _GEN_165 & ~_GEN_153;
  wire        _GEN_167 = _GEN_165 | _GEN_153;
  wire        _GEN_168 = _slots_2_io_request & (|_GEN_164) & ~_GEN_153 | _GEN_162;
  wire [9:0]  _can_allocate_T_10 = _slots_2_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_169 = _slots_2_io_request & ~_GEN_168 & (|_can_allocate_T_10);
  wire        _GEN_170 = _GEN_169 & ~_GEN_157;
  wire        _GEN_171 = _GEN_169 | _GEN_157;
  wire        _GEN_172 = _slots_2_io_request & ~(_slots_2_io_request & (|_can_allocate_T_10) & ~_GEN_157 | _GEN_168) & (|(_slots_2_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_173 = _GEN_172 & ~_GEN_160;
  assign issue_slots_2_grant = _GEN_173 | _GEN_170 | _GEN_166 | _GEN_162;
  wire        _GEN_174 = _GEN_172 | _GEN_160;
  wire        _GEN_175 = _slots_3_io_request & (|(_slots_3_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_176 = _GEN_175 & ~_GEN_163;
  wire        _GEN_177 = _GEN_175 | _GEN_163;
  wire [1:0]  _GEN_178 = {_slots_3_io_uop_fu_code[5], _slots_3_io_uop_fu_code[0]};
  wire        _GEN_179 = _slots_3_io_request & ~_GEN_176 & (|_GEN_178);
  wire        _GEN_180 = _GEN_179 & ~_GEN_167;
  wire        _GEN_181 = _GEN_179 | _GEN_167;
  wire        _GEN_182 = _slots_3_io_request & (|_GEN_178) & ~_GEN_167 | _GEN_176;
  wire [9:0]  _can_allocate_T_14 = _slots_3_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_183 = _slots_3_io_request & ~_GEN_182 & (|_can_allocate_T_14);
  wire        _GEN_184 = _GEN_183 & ~_GEN_171;
  wire        _GEN_185 = _GEN_183 | _GEN_171;
  wire        _GEN_186 = _slots_3_io_request & ~(_slots_3_io_request & (|_can_allocate_T_14) & ~_GEN_171 | _GEN_182) & (|(_slots_3_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_187 = _GEN_186 & ~_GEN_174;
  assign issue_slots_3_grant = _GEN_187 | _GEN_184 | _GEN_180 | _GEN_176;
  wire        _GEN_188 = _GEN_186 | _GEN_174;
  wire        _GEN_189 = _slots_4_io_request & (|(_slots_4_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_190 = _GEN_189 & ~_GEN_177;
  wire        _GEN_191 = _GEN_189 | _GEN_177;
  wire [1:0]  _GEN_192 = {_slots_4_io_uop_fu_code[5], _slots_4_io_uop_fu_code[0]};
  wire        _GEN_193 = _slots_4_io_request & ~_GEN_190 & (|_GEN_192);
  wire        _GEN_194 = _GEN_193 & ~_GEN_181;
  wire        _GEN_195 = _GEN_193 | _GEN_181;
  wire        _GEN_196 = _slots_4_io_request & (|_GEN_192) & ~_GEN_181 | _GEN_190;
  wire [9:0]  _can_allocate_T_18 = _slots_4_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_197 = _slots_4_io_request & ~_GEN_196 & (|_can_allocate_T_18);
  wire        _GEN_198 = _GEN_197 & ~_GEN_185;
  wire        _GEN_199 = _GEN_197 | _GEN_185;
  wire        _GEN_200 = _slots_4_io_request & ~(_slots_4_io_request & (|_can_allocate_T_18) & ~_GEN_185 | _GEN_196) & (|(_slots_4_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_201 = _GEN_200 & ~_GEN_188;
  assign issue_slots_4_grant = _GEN_201 | _GEN_198 | _GEN_194 | _GEN_190;
  wire        _GEN_202 = _GEN_200 | _GEN_188;
  wire        _GEN_203 = _slots_5_io_request & (|(_slots_5_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_204 = _GEN_203 & ~_GEN_191;
  wire        _GEN_205 = _GEN_203 | _GEN_191;
  wire [1:0]  _GEN_206 = {_slots_5_io_uop_fu_code[5], _slots_5_io_uop_fu_code[0]};
  wire        _GEN_207 = _slots_5_io_request & ~_GEN_204 & (|_GEN_206);
  wire        _GEN_208 = _GEN_207 & ~_GEN_195;
  wire        _GEN_209 = _GEN_207 | _GEN_195;
  wire        _GEN_210 = _slots_5_io_request & (|_GEN_206) & ~_GEN_195 | _GEN_204;
  wire [9:0]  _can_allocate_T_22 = _slots_5_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_211 = _slots_5_io_request & ~_GEN_210 & (|_can_allocate_T_22);
  wire        _GEN_212 = _GEN_211 & ~_GEN_199;
  wire        _GEN_213 = _GEN_211 | _GEN_199;
  wire        _GEN_214 = _slots_5_io_request & ~(_slots_5_io_request & (|_can_allocate_T_22) & ~_GEN_199 | _GEN_210) & (|(_slots_5_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_215 = _GEN_214 & ~_GEN_202;
  assign issue_slots_5_grant = _GEN_215 | _GEN_212 | _GEN_208 | _GEN_204;
  wire        _GEN_216 = _GEN_214 | _GEN_202;
  wire        _GEN_217 = _slots_6_io_request & (|(_slots_6_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_218 = _GEN_217 & ~_GEN_205;
  wire        _GEN_219 = _GEN_217 | _GEN_205;
  wire [1:0]  _GEN_220 = {_slots_6_io_uop_fu_code[5], _slots_6_io_uop_fu_code[0]};
  wire        _GEN_221 = _slots_6_io_request & ~_GEN_218 & (|_GEN_220);
  wire        _GEN_222 = _GEN_221 & ~_GEN_209;
  wire        _GEN_223 = _GEN_221 | _GEN_209;
  wire        _GEN_224 = _slots_6_io_request & (|_GEN_220) & ~_GEN_209 | _GEN_218;
  wire [9:0]  _can_allocate_T_26 = _slots_6_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_225 = _slots_6_io_request & ~_GEN_224 & (|_can_allocate_T_26);
  wire        _GEN_226 = _GEN_225 & ~_GEN_213;
  wire        _GEN_227 = _GEN_225 | _GEN_213;
  wire        _GEN_228 = _slots_6_io_request & ~(_slots_6_io_request & (|_can_allocate_T_26) & ~_GEN_213 | _GEN_224) & (|(_slots_6_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_229 = _GEN_228 & ~_GEN_216;
  assign issue_slots_6_grant = _GEN_229 | _GEN_226 | _GEN_222 | _GEN_218;
  wire        _GEN_230 = _GEN_228 | _GEN_216;
  wire        _GEN_231 = _slots_7_io_request & (|(_slots_7_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_232 = _GEN_231 & ~_GEN_219;
  wire        _GEN_233 = _GEN_231 | _GEN_219;
  wire [1:0]  _GEN_234 = {_slots_7_io_uop_fu_code[5], _slots_7_io_uop_fu_code[0]};
  wire        _GEN_235 = _slots_7_io_request & ~_GEN_232 & (|_GEN_234);
  wire        _GEN_236 = _GEN_235 & ~_GEN_223;
  wire        _GEN_237 = _GEN_235 | _GEN_223;
  wire        _GEN_238 = _slots_7_io_request & (|_GEN_234) & ~_GEN_223 | _GEN_232;
  wire [9:0]  _can_allocate_T_30 = _slots_7_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_239 = _slots_7_io_request & ~_GEN_238 & (|_can_allocate_T_30);
  wire        _GEN_240 = _GEN_239 & ~_GEN_227;
  wire        _GEN_241 = _GEN_239 | _GEN_227;
  wire        _GEN_242 = _slots_7_io_request & ~(_slots_7_io_request & (|_can_allocate_T_30) & ~_GEN_227 | _GEN_238) & (|(_slots_7_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_243 = _GEN_242 & ~_GEN_230;
  assign issue_slots_7_grant = _GEN_243 | _GEN_240 | _GEN_236 | _GEN_232;
  wire        _GEN_244 = _GEN_242 | _GEN_230;
  wire        _GEN_245 = _slots_8_io_request & (|(_slots_8_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_246 = _GEN_245 & ~_GEN_233;
  wire        _GEN_247 = _GEN_245 | _GEN_233;
  wire [1:0]  _GEN_248 = {_slots_8_io_uop_fu_code[5], _slots_8_io_uop_fu_code[0]};
  wire        _GEN_249 = _slots_8_io_request & ~_GEN_246 & (|_GEN_248);
  wire        _GEN_250 = _GEN_249 & ~_GEN_237;
  wire        _GEN_251 = _GEN_249 | _GEN_237;
  wire        _GEN_252 = _slots_8_io_request & (|_GEN_248) & ~_GEN_237 | _GEN_246;
  wire [9:0]  _can_allocate_T_34 = _slots_8_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_253 = _slots_8_io_request & ~_GEN_252 & (|_can_allocate_T_34);
  wire        _GEN_254 = _GEN_253 & ~_GEN_241;
  wire        _GEN_255 = _GEN_253 | _GEN_241;
  wire        _GEN_256 = _slots_8_io_request & ~(_slots_8_io_request & (|_can_allocate_T_34) & ~_GEN_241 | _GEN_252) & (|(_slots_8_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_257 = _GEN_256 & ~_GEN_244;
  assign issue_slots_8_grant = _GEN_257 | _GEN_254 | _GEN_250 | _GEN_246;
  wire        _GEN_258 = _GEN_256 | _GEN_244;
  wire        _GEN_259 = _slots_9_io_request & (|(_slots_9_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_260 = _GEN_259 & ~_GEN_247;
  wire        _GEN_261 = _GEN_259 | _GEN_247;
  wire [1:0]  _GEN_262 = {_slots_9_io_uop_fu_code[5], _slots_9_io_uop_fu_code[0]};
  wire        _GEN_263 = _slots_9_io_request & ~_GEN_260 & (|_GEN_262);
  wire        _GEN_264 = _GEN_263 & ~_GEN_251;
  wire        _GEN_265 = _GEN_263 | _GEN_251;
  wire        _GEN_266 = _slots_9_io_request & (|_GEN_262) & ~_GEN_251 | _GEN_260;
  wire [9:0]  _can_allocate_T_38 = _slots_9_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_267 = _slots_9_io_request & ~_GEN_266 & (|_can_allocate_T_38);
  wire        _GEN_268 = _GEN_267 & ~_GEN_255;
  wire        _GEN_269 = _GEN_267 | _GEN_255;
  wire        _GEN_270 = _slots_9_io_request & ~(_slots_9_io_request & (|_can_allocate_T_38) & ~_GEN_255 | _GEN_266) & (|(_slots_9_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_271 = _GEN_270 & ~_GEN_258;
  assign issue_slots_9_grant = _GEN_271 | _GEN_268 | _GEN_264 | _GEN_260;
  wire        _GEN_272 = _GEN_270 | _GEN_258;
  wire        _GEN_273 = _slots_10_io_request & (|(_slots_10_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_274 = _GEN_273 & ~_GEN_261;
  wire        _GEN_275 = _GEN_273 | _GEN_261;
  wire [1:0]  _GEN_276 = {_slots_10_io_uop_fu_code[5], _slots_10_io_uop_fu_code[0]};
  wire        _GEN_277 = _slots_10_io_request & ~_GEN_274 & (|_GEN_276);
  wire        _GEN_278 = _GEN_277 & ~_GEN_265;
  wire        _GEN_279 = _GEN_277 | _GEN_265;
  wire        _GEN_280 = _slots_10_io_request & (|_GEN_276) & ~_GEN_265 | _GEN_274;
  wire [9:0]  _can_allocate_T_42 = _slots_10_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_281 = _slots_10_io_request & ~_GEN_280 & (|_can_allocate_T_42);
  wire        _GEN_282 = _GEN_281 & ~_GEN_269;
  wire        _GEN_283 = _GEN_281 | _GEN_269;
  wire        _GEN_284 = _slots_10_io_request & ~(_slots_10_io_request & (|_can_allocate_T_42) & ~_GEN_269 | _GEN_280) & (|(_slots_10_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_285 = _GEN_284 & ~_GEN_272;
  assign issue_slots_10_grant = _GEN_285 | _GEN_282 | _GEN_278 | _GEN_274;
  wire        _GEN_286 = _GEN_284 | _GEN_272;
  wire        _GEN_287 = _slots_11_io_request & (|(_slots_11_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_288 = _GEN_287 & ~_GEN_275;
  wire        _GEN_289 = _GEN_287 | _GEN_275;
  wire [1:0]  _GEN_290 = {_slots_11_io_uop_fu_code[5], _slots_11_io_uop_fu_code[0]};
  wire        _GEN_291 = _slots_11_io_request & ~_GEN_288 & (|_GEN_290);
  wire        _GEN_292 = _GEN_291 & ~_GEN_279;
  wire        _GEN_293 = _GEN_291 | _GEN_279;
  wire        _GEN_294 = _slots_11_io_request & (|_GEN_290) & ~_GEN_279 | _GEN_288;
  wire [9:0]  _can_allocate_T_46 = _slots_11_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_295 = _slots_11_io_request & ~_GEN_294 & (|_can_allocate_T_46);
  wire        _GEN_296 = _GEN_295 & ~_GEN_283;
  wire        _GEN_297 = _GEN_295 | _GEN_283;
  wire        _GEN_298 = _slots_11_io_request & ~(_slots_11_io_request & (|_can_allocate_T_46) & ~_GEN_283 | _GEN_294) & (|(_slots_11_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_299 = _GEN_298 & ~_GEN_286;
  assign issue_slots_11_grant = _GEN_299 | _GEN_296 | _GEN_292 | _GEN_288;
  wire        _GEN_300 = _GEN_298 | _GEN_286;
  wire        _GEN_301 = _slots_12_io_request & (|(_slots_12_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_302 = _GEN_301 & ~_GEN_289;
  wire        _GEN_303 = _GEN_301 | _GEN_289;
  wire [1:0]  _GEN_304 = {_slots_12_io_uop_fu_code[5], _slots_12_io_uop_fu_code[0]};
  wire        _GEN_305 = _slots_12_io_request & ~_GEN_302 & (|_GEN_304);
  wire        _GEN_306 = _GEN_305 & ~_GEN_293;
  wire        _GEN_307 = _GEN_305 | _GEN_293;
  wire        _GEN_308 = _slots_12_io_request & (|_GEN_304) & ~_GEN_293 | _GEN_302;
  wire [9:0]  _can_allocate_T_50 = _slots_12_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_309 = _slots_12_io_request & ~_GEN_308 & (|_can_allocate_T_50);
  wire        _GEN_310 = _GEN_309 & ~_GEN_297;
  wire        _GEN_311 = _GEN_309 | _GEN_297;
  wire        _GEN_312 = _slots_12_io_request & ~(_slots_12_io_request & (|_can_allocate_T_50) & ~_GEN_297 | _GEN_308) & (|(_slots_12_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_313 = _GEN_312 & ~_GEN_300;
  assign issue_slots_12_grant = _GEN_313 | _GEN_310 | _GEN_306 | _GEN_302;
  wire        _GEN_314 = _GEN_312 | _GEN_300;
  wire        _GEN_315 = _slots_13_io_request & (|(_slots_13_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_316 = _GEN_315 & ~_GEN_303;
  wire        _GEN_317 = _GEN_315 | _GEN_303;
  wire [1:0]  _GEN_318 = {_slots_13_io_uop_fu_code[5], _slots_13_io_uop_fu_code[0]};
  wire        _GEN_319 = _slots_13_io_request & ~_GEN_316 & (|_GEN_318);
  wire        _GEN_320 = _GEN_319 & ~_GEN_307;
  wire        _GEN_321 = _GEN_319 | _GEN_307;
  wire        _GEN_322 = _slots_13_io_request & (|_GEN_318) & ~_GEN_307 | _GEN_316;
  wire [9:0]  _can_allocate_T_54 = _slots_13_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_323 = _slots_13_io_request & ~_GEN_322 & (|_can_allocate_T_54);
  wire        _GEN_324 = _GEN_323 & ~_GEN_311;
  wire        _GEN_325 = _GEN_323 | _GEN_311;
  wire        _GEN_326 = _slots_13_io_request & ~(_slots_13_io_request & (|_can_allocate_T_54) & ~_GEN_311 | _GEN_322) & (|(_slots_13_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_327 = _GEN_326 & ~_GEN_314;
  assign issue_slots_13_grant = _GEN_327 | _GEN_324 | _GEN_320 | _GEN_316;
  wire        _GEN_328 = _GEN_326 | _GEN_314;
  wire        _GEN_329 = _slots_14_io_request & (|(_slots_14_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_330 = _GEN_329 & ~_GEN_317;
  wire        _GEN_331 = _GEN_329 | _GEN_317;
  wire [1:0]  _GEN_332 = {_slots_14_io_uop_fu_code[5], _slots_14_io_uop_fu_code[0]};
  wire        _GEN_333 = _slots_14_io_request & ~_GEN_330 & (|_GEN_332);
  wire        _GEN_334 = _GEN_333 & ~_GEN_321;
  wire        _GEN_335 = _GEN_333 | _GEN_321;
  wire        _GEN_336 = _slots_14_io_request & (|_GEN_332) & ~_GEN_321 | _GEN_330;
  wire [9:0]  _can_allocate_T_58 = _slots_14_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_337 = _slots_14_io_request & ~_GEN_336 & (|_can_allocate_T_58);
  wire        _GEN_338 = _GEN_337 & ~_GEN_325;
  wire        _GEN_339 = _GEN_337 | _GEN_325;
  wire        _GEN_340 = _slots_14_io_request & ~(_slots_14_io_request & (|_can_allocate_T_58) & ~_GEN_325 | _GEN_336) & (|(_slots_14_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_341 = _GEN_340 & ~_GEN_328;
  assign issue_slots_14_grant = _GEN_341 | _GEN_338 | _GEN_334 | _GEN_330;
  wire        _GEN_342 = _GEN_340 | _GEN_328;
  wire        _GEN_343 = _slots_15_io_request & (|(_slots_15_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_344 = _GEN_343 & ~_GEN_331;
  wire        _GEN_345 = _GEN_343 | _GEN_331;
  wire [1:0]  _GEN_346 = {_slots_15_io_uop_fu_code[5], _slots_15_io_uop_fu_code[0]};
  wire        _GEN_347 = _slots_15_io_request & ~_GEN_344 & (|_GEN_346);
  wire        _GEN_348 = _GEN_347 & ~_GEN_335;
  wire        _GEN_349 = _GEN_347 | _GEN_335;
  wire        _GEN_350 = _slots_15_io_request & (|_GEN_346) & ~_GEN_335 | _GEN_344;
  wire [9:0]  _can_allocate_T_62 = _slots_15_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_351 = _slots_15_io_request & ~_GEN_350 & (|_can_allocate_T_62);
  wire        _GEN_352 = _GEN_351 & ~_GEN_339;
  wire        _GEN_353 = _GEN_351 | _GEN_339;
  wire        _GEN_354 = _slots_15_io_request & ~(_slots_15_io_request & (|_can_allocate_T_62) & ~_GEN_339 | _GEN_350) & (|(_slots_15_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_355 = _GEN_354 & ~_GEN_342;
  assign issue_slots_15_grant = _GEN_355 | _GEN_352 | _GEN_348 | _GEN_344;
  wire        _GEN_356 = _GEN_354 | _GEN_342;
  wire        _GEN_357 = _slots_16_io_request & (|(_slots_16_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_358 = _GEN_357 & ~_GEN_345;
  wire        _GEN_359 = _GEN_357 | _GEN_345;
  wire [1:0]  _GEN_360 = {_slots_16_io_uop_fu_code[5], _slots_16_io_uop_fu_code[0]};
  wire        _GEN_361 = _slots_16_io_request & ~_GEN_358 & (|_GEN_360);
  wire        _GEN_362 = _GEN_361 & ~_GEN_349;
  wire        _GEN_363 = _GEN_361 | _GEN_349;
  wire        _GEN_364 = _slots_16_io_request & (|_GEN_360) & ~_GEN_349 | _GEN_358;
  wire [9:0]  _can_allocate_T_66 = _slots_16_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_365 = _slots_16_io_request & ~_GEN_364 & (|_can_allocate_T_66);
  wire        _GEN_366 = _GEN_365 & ~_GEN_353;
  wire        _GEN_367 = _GEN_365 | _GEN_353;
  wire        _GEN_368 = _slots_16_io_request & ~(_slots_16_io_request & (|_can_allocate_T_66) & ~_GEN_353 | _GEN_364) & (|(_slots_16_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_369 = _GEN_368 & ~_GEN_356;
  assign issue_slots_16_grant = _GEN_369 | _GEN_366 | _GEN_362 | _GEN_358;
  wire        _GEN_370 = _GEN_368 | _GEN_356;
  wire        _GEN_371 = _slots_17_io_request & (|(_slots_17_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_372 = _GEN_371 & ~_GEN_359;
  wire        _GEN_373 = _GEN_371 | _GEN_359;
  wire [1:0]  _GEN_374 = {_slots_17_io_uop_fu_code[5], _slots_17_io_uop_fu_code[0]};
  wire        _GEN_375 = _slots_17_io_request & ~_GEN_372 & (|_GEN_374);
  wire        _GEN_376 = _GEN_375 & ~_GEN_363;
  wire        _GEN_377 = _GEN_375 | _GEN_363;
  wire        _GEN_378 = _slots_17_io_request & (|_GEN_374) & ~_GEN_363 | _GEN_372;
  wire [9:0]  _can_allocate_T_70 = _slots_17_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_379 = _slots_17_io_request & ~_GEN_378 & (|_can_allocate_T_70);
  wire        _GEN_380 = _GEN_379 & ~_GEN_367;
  wire        _GEN_381 = _GEN_379 | _GEN_367;
  wire        _GEN_382 = _slots_17_io_request & ~(_slots_17_io_request & (|_can_allocate_T_70) & ~_GEN_367 | _GEN_378) & (|(_slots_17_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_383 = _GEN_382 & ~_GEN_370;
  assign issue_slots_17_grant = _GEN_383 | _GEN_380 | _GEN_376 | _GEN_372;
  wire        _GEN_384 = _GEN_382 | _GEN_370;
  wire        _GEN_385 = _slots_18_io_request & (|(_slots_18_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_386 = _GEN_385 & ~_GEN_373;
  wire        _GEN_387 = _GEN_385 | _GEN_373;
  wire [1:0]  _GEN_388 = {_slots_18_io_uop_fu_code[5], _slots_18_io_uop_fu_code[0]};
  wire        _GEN_389 = _slots_18_io_request & ~_GEN_386 & (|_GEN_388);
  wire        _GEN_390 = _GEN_389 & ~_GEN_377;
  wire        _GEN_391 = _GEN_389 | _GEN_377;
  wire        _GEN_392 = _slots_18_io_request & (|_GEN_388) & ~_GEN_377 | _GEN_386;
  wire [9:0]  _can_allocate_T_74 = _slots_18_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_393 = _slots_18_io_request & ~_GEN_392 & (|_can_allocate_T_74);
  wire        _GEN_394 = _GEN_393 & ~_GEN_381;
  wire        _GEN_395 = _GEN_393 | _GEN_381;
  wire        _GEN_396 = _slots_18_io_request & ~(_slots_18_io_request & (|_can_allocate_T_74) & ~_GEN_381 | _GEN_392) & (|(_slots_18_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_397 = _GEN_396 & ~_GEN_384;
  assign issue_slots_18_grant = _GEN_397 | _GEN_394 | _GEN_390 | _GEN_386;
  wire        _GEN_398 = _GEN_396 | _GEN_384;
  wire        _GEN_399 = _slots_19_io_request & (|(_slots_19_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_400 = _GEN_399 & ~_GEN_387;
  wire        _GEN_401 = _GEN_399 | _GEN_387;
  wire [1:0]  _GEN_402 = {_slots_19_io_uop_fu_code[5], _slots_19_io_uop_fu_code[0]};
  wire        _GEN_403 = _slots_19_io_request & ~_GEN_400 & (|_GEN_402);
  wire        _GEN_404 = _GEN_403 & ~_GEN_391;
  wire        _GEN_405 = _GEN_403 | _GEN_391;
  wire        _GEN_406 = _slots_19_io_request & (|_GEN_402) & ~_GEN_391 | _GEN_400;
  wire [9:0]  _can_allocate_T_78 = _slots_19_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_407 = _slots_19_io_request & ~_GEN_406 & (|_can_allocate_T_78);
  wire        _GEN_408 = _GEN_407 & ~_GEN_395;
  wire        _GEN_409 = _GEN_407 | _GEN_395;
  wire        _GEN_410 = _slots_19_io_request & ~(_slots_19_io_request & (|_can_allocate_T_78) & ~_GEN_395 | _GEN_406) & (|(_slots_19_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_411 = _GEN_410 & ~_GEN_398;
  assign issue_slots_19_grant = _GEN_411 | _GEN_408 | _GEN_404 | _GEN_400;
  wire        _GEN_412 = _GEN_410 | _GEN_398;
  wire        _GEN_413 = _slots_20_io_request & (|(_slots_20_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_414 = _GEN_413 & ~_GEN_401;
  wire        _GEN_415 = _GEN_413 | _GEN_401;
  wire [1:0]  _GEN_416 = {_slots_20_io_uop_fu_code[5], _slots_20_io_uop_fu_code[0]};
  wire        _GEN_417 = _slots_20_io_request & ~_GEN_414 & (|_GEN_416);
  wire        _GEN_418 = _GEN_417 & ~_GEN_405;
  wire        _GEN_419 = _GEN_417 | _GEN_405;
  wire        _GEN_420 = _slots_20_io_request & (|_GEN_416) & ~_GEN_405 | _GEN_414;
  wire [9:0]  _can_allocate_T_82 = _slots_20_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_421 = _slots_20_io_request & ~_GEN_420 & (|_can_allocate_T_82);
  wire        _GEN_422 = _GEN_421 & ~_GEN_409;
  wire        _GEN_423 = _GEN_421 | _GEN_409;
  wire        _GEN_424 = _slots_20_io_request & ~(_slots_20_io_request & (|_can_allocate_T_82) & ~_GEN_409 | _GEN_420) & (|(_slots_20_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_425 = _GEN_424 & ~_GEN_412;
  assign issue_slots_20_grant = _GEN_425 | _GEN_422 | _GEN_418 | _GEN_414;
  wire        _GEN_426 = _GEN_424 | _GEN_412;
  wire        _GEN_427 = _slots_21_io_request & (|(_slots_21_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_428 = _GEN_427 & ~_GEN_415;
  wire        _GEN_429 = _GEN_427 | _GEN_415;
  wire [1:0]  _GEN_430 = {_slots_21_io_uop_fu_code[5], _slots_21_io_uop_fu_code[0]};
  wire        _GEN_431 = _slots_21_io_request & ~_GEN_428 & (|_GEN_430);
  wire        _GEN_432 = _GEN_431 & ~_GEN_419;
  wire        _GEN_433 = _GEN_431 | _GEN_419;
  wire        _GEN_434 = _slots_21_io_request & (|_GEN_430) & ~_GEN_419 | _GEN_428;
  wire [9:0]  _can_allocate_T_86 = _slots_21_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_435 = _slots_21_io_request & ~_GEN_434 & (|_can_allocate_T_86);
  wire        _GEN_436 = _GEN_435 & ~_GEN_423;
  wire        _GEN_437 = _GEN_435 | _GEN_423;
  wire        _GEN_438 = _slots_21_io_request & ~(_slots_21_io_request & (|_can_allocate_T_86) & ~_GEN_423 | _GEN_434) & (|(_slots_21_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_439 = _GEN_438 & ~_GEN_426;
  assign issue_slots_21_grant = _GEN_439 | _GEN_436 | _GEN_432 | _GEN_428;
  wire        _GEN_440 = _GEN_438 | _GEN_426;
  wire        _GEN_441 = _slots_22_io_request & (|(_slots_22_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_442 = _GEN_441 & ~_GEN_429;
  wire        _GEN_443 = _GEN_441 | _GEN_429;
  wire [1:0]  _GEN_444 = {_slots_22_io_uop_fu_code[5], _slots_22_io_uop_fu_code[0]};
  wire        _GEN_445 = _slots_22_io_request & ~_GEN_442 & (|_GEN_444);
  wire        _GEN_446 = _GEN_445 & ~_GEN_433;
  wire        _GEN_447 = _GEN_445 | _GEN_433;
  wire        _GEN_448 = _slots_22_io_request & (|_GEN_444) & ~_GEN_433 | _GEN_442;
  wire [9:0]  _can_allocate_T_90 = _slots_22_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_449 = _slots_22_io_request & ~_GEN_448 & (|_can_allocate_T_90);
  wire        _GEN_450 = _GEN_449 & ~_GEN_437;
  wire        _GEN_451 = _GEN_449 | _GEN_437;
  wire        _GEN_452 = _slots_22_io_request & ~(_slots_22_io_request & (|_can_allocate_T_90) & ~_GEN_437 | _GEN_448) & (|(_slots_22_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_453 = _GEN_452 & ~_GEN_440;
  assign issue_slots_22_grant = _GEN_453 | _GEN_450 | _GEN_446 | _GEN_442;
  wire        _GEN_454 = _GEN_452 | _GEN_440;
  wire        _GEN_455 = _slots_23_io_request & (|(_slots_23_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_456 = _GEN_455 & ~_GEN_443;
  wire        _GEN_457 = _GEN_455 | _GEN_443;
  wire [1:0]  _GEN_458 = {_slots_23_io_uop_fu_code[5], _slots_23_io_uop_fu_code[0]};
  wire        _GEN_459 = _slots_23_io_request & ~_GEN_456 & (|_GEN_458);
  wire        _GEN_460 = _GEN_459 & ~_GEN_447;
  wire        _GEN_461 = _GEN_459 | _GEN_447;
  wire        _GEN_462 = _slots_23_io_request & (|_GEN_458) & ~_GEN_447 | _GEN_456;
  wire [9:0]  _can_allocate_T_94 = _slots_23_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_463 = _slots_23_io_request & ~_GEN_462 & (|_can_allocate_T_94);
  wire        _GEN_464 = _GEN_463 & ~_GEN_451;
  wire        _GEN_465 = _GEN_463 | _GEN_451;
  wire        _GEN_466 = _slots_23_io_request & ~(_slots_23_io_request & (|_can_allocate_T_94) & ~_GEN_451 | _GEN_462) & (|(_slots_23_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_467 = _GEN_466 & ~_GEN_454;
  assign issue_slots_23_grant = _GEN_467 | _GEN_464 | _GEN_460 | _GEN_456;
  wire        _GEN_468 = _GEN_466 | _GEN_454;
  wire        _GEN_469 = _slots_24_io_request & (|(_slots_24_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_470 = _GEN_469 & ~_GEN_457;
  wire        _GEN_471 = _GEN_469 | _GEN_457;
  wire [1:0]  _GEN_472 = {_slots_24_io_uop_fu_code[5], _slots_24_io_uop_fu_code[0]};
  wire        _GEN_473 = _slots_24_io_request & ~_GEN_470 & (|_GEN_472);
  wire        _GEN_474 = _GEN_473 & ~_GEN_461;
  wire        _GEN_475 = _GEN_473 | _GEN_461;
  wire        _GEN_476 = _slots_24_io_request & (|_GEN_472) & ~_GEN_461 | _GEN_470;
  wire [9:0]  _can_allocate_T_98 = _slots_24_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_477 = _slots_24_io_request & ~_GEN_476 & (|_can_allocate_T_98);
  wire        _GEN_478 = _GEN_477 & ~_GEN_465;
  wire        _GEN_479 = _GEN_477 | _GEN_465;
  wire        _GEN_480 = _slots_24_io_request & ~(_slots_24_io_request & (|_can_allocate_T_98) & ~_GEN_465 | _GEN_476) & (|(_slots_24_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_481 = _GEN_480 & ~_GEN_468;
  assign issue_slots_24_grant = _GEN_481 | _GEN_478 | _GEN_474 | _GEN_470;
  wire        _GEN_482 = _GEN_480 | _GEN_468;
  wire        _GEN_483 = _slots_25_io_request & (|(_slots_25_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_484 = _GEN_483 & ~_GEN_471;
  wire        _GEN_485 = _GEN_483 | _GEN_471;
  wire [1:0]  _GEN_486 = {_slots_25_io_uop_fu_code[5], _slots_25_io_uop_fu_code[0]};
  wire        _GEN_487 = _slots_25_io_request & ~_GEN_484 & (|_GEN_486);
  wire        _GEN_488 = _GEN_487 & ~_GEN_475;
  wire        _GEN_489 = _GEN_487 | _GEN_475;
  wire        _GEN_490 = _slots_25_io_request & (|_GEN_486) & ~_GEN_475 | _GEN_484;
  wire [9:0]  _can_allocate_T_102 = _slots_25_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_491 = _slots_25_io_request & ~_GEN_490 & (|_can_allocate_T_102);
  wire        _GEN_492 = _GEN_491 & ~_GEN_479;
  wire        _GEN_493 = _GEN_491 | _GEN_479;
  wire        _GEN_494 = _slots_25_io_request & ~(_slots_25_io_request & (|_can_allocate_T_102) & ~_GEN_479 | _GEN_490) & (|(_slots_25_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_495 = _GEN_494 & ~_GEN_482;
  assign issue_slots_25_grant = _GEN_495 | _GEN_492 | _GEN_488 | _GEN_484;
  wire        _GEN_496 = _GEN_494 | _GEN_482;
  wire        _GEN_497 = _slots_26_io_request & (|(_slots_26_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_498 = _GEN_497 & ~_GEN_485;
  wire        _GEN_499 = _GEN_497 | _GEN_485;
  wire [1:0]  _GEN_500 = {_slots_26_io_uop_fu_code[5], _slots_26_io_uop_fu_code[0]};
  wire        _GEN_501 = _slots_26_io_request & ~_GEN_498 & (|_GEN_500);
  wire        _GEN_502 = _GEN_501 & ~_GEN_489;
  wire        _GEN_503 = _GEN_501 | _GEN_489;
  wire        _GEN_504 = _slots_26_io_request & (|_GEN_500) & ~_GEN_489 | _GEN_498;
  wire [9:0]  _can_allocate_T_106 = _slots_26_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_505 = _slots_26_io_request & ~_GEN_504 & (|_can_allocate_T_106);
  wire        _GEN_506 = _GEN_505 & ~_GEN_493;
  wire        _GEN_507 = _GEN_505 | _GEN_493;
  wire        _GEN_508 = _slots_26_io_request & ~(_slots_26_io_request & (|_can_allocate_T_106) & ~_GEN_493 | _GEN_504) & (|(_slots_26_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_509 = _GEN_508 & ~_GEN_496;
  assign issue_slots_26_grant = _GEN_509 | _GEN_506 | _GEN_502 | _GEN_498;
  wire        _GEN_510 = _GEN_508 | _GEN_496;
  wire        _GEN_511 = _slots_27_io_request & (|(_slots_27_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_512 = _GEN_511 & ~_GEN_499;
  wire        _GEN_513 = _GEN_511 | _GEN_499;
  wire [1:0]  _GEN_514 = {_slots_27_io_uop_fu_code[5], _slots_27_io_uop_fu_code[0]};
  wire        _GEN_515 = _slots_27_io_request & ~_GEN_512 & (|_GEN_514);
  wire        _GEN_516 = _GEN_515 & ~_GEN_503;
  wire        _GEN_517 = _GEN_515 | _GEN_503;
  wire        _GEN_518 = _slots_27_io_request & (|_GEN_514) & ~_GEN_503 | _GEN_512;
  wire [9:0]  _can_allocate_T_110 = _slots_27_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_519 = _slots_27_io_request & ~_GEN_518 & (|_can_allocate_T_110);
  wire        _GEN_520 = _GEN_519 & ~_GEN_507;
  wire        _GEN_521 = _GEN_519 | _GEN_507;
  wire        _GEN_522 = _slots_27_io_request & ~(_slots_27_io_request & (|_can_allocate_T_110) & ~_GEN_507 | _GEN_518) & (|(_slots_27_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_523 = _GEN_522 & ~_GEN_510;
  assign issue_slots_27_grant = _GEN_523 | _GEN_520 | _GEN_516 | _GEN_512;
  wire        _GEN_524 = _GEN_522 | _GEN_510;
  wire        _GEN_525 = _slots_28_io_request & (|(_slots_28_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_526 = _GEN_525 & ~_GEN_513;
  wire        _GEN_527 = _GEN_525 | _GEN_513;
  wire [1:0]  _GEN_528 = {_slots_28_io_uop_fu_code[5], _slots_28_io_uop_fu_code[0]};
  wire        _GEN_529 = _slots_28_io_request & ~_GEN_526 & (|_GEN_528);
  wire        _GEN_530 = _GEN_529 & ~_GEN_517;
  wire        _GEN_531 = _GEN_529 | _GEN_517;
  wire        _GEN_532 = _slots_28_io_request & (|_GEN_528) & ~_GEN_517 | _GEN_526;
  wire [9:0]  _can_allocate_T_114 = _slots_28_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_533 = _slots_28_io_request & ~_GEN_532 & (|_can_allocate_T_114);
  wire        _GEN_534 = _GEN_533 & ~_GEN_521;
  wire        _GEN_535 = _GEN_533 | _GEN_521;
  wire        _GEN_536 = _slots_28_io_request & ~(_slots_28_io_request & (|_can_allocate_T_114) & ~_GEN_521 | _GEN_532) & (|(_slots_28_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_537 = _GEN_536 & ~_GEN_524;
  assign issue_slots_28_grant = _GEN_537 | _GEN_534 | _GEN_530 | _GEN_526;
  wire        _GEN_538 = _GEN_536 | _GEN_524;
  wire        _GEN_539 = _slots_29_io_request & (|(_slots_29_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_540 = _GEN_539 & ~_GEN_527;
  wire        _GEN_541 = _GEN_539 | _GEN_527;
  wire [1:0]  _GEN_542 = {_slots_29_io_uop_fu_code[5], _slots_29_io_uop_fu_code[0]};
  wire        _GEN_543 = _slots_29_io_request & ~_GEN_540 & (|_GEN_542);
  wire        _GEN_544 = _GEN_543 & ~_GEN_531;
  wire        _GEN_545 = _GEN_543 | _GEN_531;
  wire        _GEN_546 = _slots_29_io_request & (|_GEN_542) & ~_GEN_531 | _GEN_540;
  wire [9:0]  _can_allocate_T_118 = _slots_29_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_547 = _slots_29_io_request & ~_GEN_546 & (|_can_allocate_T_118);
  wire        _GEN_548 = _GEN_547 & ~_GEN_535;
  wire        _GEN_549 = _GEN_547 | _GEN_535;
  wire        _GEN_550 = _slots_29_io_request & ~(_slots_29_io_request & (|_can_allocate_T_118) & ~_GEN_535 | _GEN_546) & (|(_slots_29_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_551 = _GEN_550 & ~_GEN_538;
  assign issue_slots_29_grant = _GEN_551 | _GEN_548 | _GEN_544 | _GEN_540;
  wire        _GEN_552 = _GEN_550 | _GEN_538;
  wire        _GEN_553 = _slots_30_io_request & (|(_slots_30_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_554 = _GEN_553 & ~_GEN_541;
  wire        _GEN_555 = _GEN_553 | _GEN_541;
  wire [1:0]  _GEN_556 = {_slots_30_io_uop_fu_code[5], _slots_30_io_uop_fu_code[0]};
  wire        _GEN_557 = _slots_30_io_request & ~_GEN_554 & (|_GEN_556);
  wire        _GEN_558 = _GEN_557 & ~_GEN_545;
  wire        _GEN_559 = _GEN_557 | _GEN_545;
  wire        _GEN_560 = _slots_30_io_request & (|_GEN_556) & ~_GEN_545 | _GEN_554;
  wire [9:0]  _can_allocate_T_122 = _slots_30_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_561 = _slots_30_io_request & ~_GEN_560 & (|_can_allocate_T_122);
  wire        _GEN_562 = _GEN_561 & ~_GEN_549;
  wire        _GEN_563 = _GEN_561 | _GEN_549;
  wire        _GEN_564 = _slots_30_io_request & ~(_slots_30_io_request & (|_can_allocate_T_122) & ~_GEN_549 | _GEN_560) & (|(_slots_30_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_565 = _GEN_564 & ~_GEN_552;
  assign issue_slots_30_grant = _GEN_565 | _GEN_562 | _GEN_558 | _GEN_554;
  wire        _GEN_566 = _GEN_564 | _GEN_552;
  wire        _GEN_567 = _slots_31_io_request & (|(_slots_31_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_568 = _GEN_567 & ~_GEN_555;
  wire        _GEN_569 = _GEN_567 | _GEN_555;
  wire [1:0]  _GEN_570 = {_slots_31_io_uop_fu_code[5], _slots_31_io_uop_fu_code[0]};
  wire        _GEN_571 = _slots_31_io_request & ~_GEN_568 & (|_GEN_570);
  wire        _GEN_572 = _GEN_571 & ~_GEN_559;
  wire        _GEN_573 = _GEN_571 | _GEN_559;
  wire        _GEN_574 = _slots_31_io_request & (|_GEN_570) & ~_GEN_559 | _GEN_568;
  wire [9:0]  _can_allocate_T_126 = _slots_31_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_575 = _slots_31_io_request & ~_GEN_574 & (|_can_allocate_T_126);
  wire        _GEN_576 = _GEN_575 & ~_GEN_563;
  wire        _GEN_577 = _GEN_575 | _GEN_563;
  wire        _GEN_578 = _slots_31_io_request & ~(_slots_31_io_request & (|_can_allocate_T_126) & ~_GEN_563 | _GEN_574) & (|(_slots_31_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_579 = _GEN_578 & ~_GEN_566;
  assign issue_slots_31_grant = _GEN_579 | _GEN_576 | _GEN_572 | _GEN_568;
  wire        _GEN_580 = _GEN_578 | _GEN_566;
  wire        _GEN_581 = _slots_32_io_request & (|(_slots_32_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_582 = _GEN_581 & ~_GEN_569;
  wire        _GEN_583 = _GEN_581 | _GEN_569;
  wire [1:0]  _GEN_584 = {_slots_32_io_uop_fu_code[5], _slots_32_io_uop_fu_code[0]};
  wire        _GEN_585 = _slots_32_io_request & ~_GEN_582 & (|_GEN_584);
  wire        _GEN_586 = _GEN_585 & ~_GEN_573;
  wire        _GEN_587 = _GEN_585 | _GEN_573;
  wire        _GEN_588 = _slots_32_io_request & (|_GEN_584) & ~_GEN_573 | _GEN_582;
  wire [9:0]  _can_allocate_T_130 = _slots_32_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_589 = _slots_32_io_request & ~_GEN_588 & (|_can_allocate_T_130);
  wire        _GEN_590 = _GEN_589 & ~_GEN_577;
  wire        _GEN_591 = _GEN_589 | _GEN_577;
  wire        _GEN_592 = _slots_32_io_request & ~(_slots_32_io_request & (|_can_allocate_T_130) & ~_GEN_577 | _GEN_588) & (|(_slots_32_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_593 = _GEN_592 & ~_GEN_580;
  assign issue_slots_32_grant = _GEN_593 | _GEN_590 | _GEN_586 | _GEN_582;
  wire        _GEN_594 = _GEN_592 | _GEN_580;
  wire        _GEN_595 = _slots_33_io_request & (|(_slots_33_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_596 = _GEN_595 & ~_GEN_583;
  wire        _GEN_597 = _GEN_595 | _GEN_583;
  wire [1:0]  _GEN_598 = {_slots_33_io_uop_fu_code[5], _slots_33_io_uop_fu_code[0]};
  wire        _GEN_599 = _slots_33_io_request & ~_GEN_596 & (|_GEN_598);
  wire        _GEN_600 = _GEN_599 & ~_GEN_587;
  wire        _GEN_601 = _GEN_599 | _GEN_587;
  wire        _GEN_602 = _slots_33_io_request & (|_GEN_598) & ~_GEN_587 | _GEN_596;
  wire [9:0]  _can_allocate_T_134 = _slots_33_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_603 = _slots_33_io_request & ~_GEN_602 & (|_can_allocate_T_134);
  wire        _GEN_604 = _GEN_603 & ~_GEN_591;
  wire        _GEN_605 = _GEN_603 | _GEN_591;
  wire        _GEN_606 = _slots_33_io_request & ~(_slots_33_io_request & (|_can_allocate_T_134) & ~_GEN_591 | _GEN_602) & (|(_slots_33_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_607 = _GEN_606 & ~_GEN_594;
  assign issue_slots_33_grant = _GEN_607 | _GEN_604 | _GEN_600 | _GEN_596;
  wire        _GEN_608 = _GEN_606 | _GEN_594;
  wire        _GEN_609 = _slots_34_io_request & (|(_slots_34_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_610 = _GEN_609 & ~_GEN_597;
  wire        _GEN_611 = _GEN_609 | _GEN_597;
  wire [1:0]  _GEN_612 = {_slots_34_io_uop_fu_code[5], _slots_34_io_uop_fu_code[0]};
  wire        _GEN_613 = _slots_34_io_request & ~_GEN_610 & (|_GEN_612);
  wire        _GEN_614 = _GEN_613 & ~_GEN_601;
  wire        _GEN_615 = _GEN_613 | _GEN_601;
  wire        _GEN_616 = _slots_34_io_request & (|_GEN_612) & ~_GEN_601 | _GEN_610;
  wire [9:0]  _can_allocate_T_138 = _slots_34_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_617 = _slots_34_io_request & ~_GEN_616 & (|_can_allocate_T_138);
  wire        _GEN_618 = _GEN_617 & ~_GEN_605;
  wire        _GEN_619 = _GEN_617 | _GEN_605;
  wire        _GEN_620 = _slots_34_io_request & ~(_slots_34_io_request & (|_can_allocate_T_138) & ~_GEN_605 | _GEN_616) & (|(_slots_34_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_621 = _GEN_620 & ~_GEN_608;
  assign issue_slots_34_grant = _GEN_621 | _GEN_618 | _GEN_614 | _GEN_610;
  wire        _GEN_622 = _GEN_620 | _GEN_608;
  wire        _GEN_623 = _slots_35_io_request & (|(_slots_35_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_624 = _GEN_623 & ~_GEN_611;
  wire        _GEN_625 = _GEN_623 | _GEN_611;
  wire [1:0]  _GEN_626 = {_slots_35_io_uop_fu_code[5], _slots_35_io_uop_fu_code[0]};
  wire        _GEN_627 = _slots_35_io_request & ~_GEN_624 & (|_GEN_626);
  wire        _GEN_628 = _GEN_627 & ~_GEN_615;
  wire        _GEN_629 = _GEN_627 | _GEN_615;
  wire        _GEN_630 = _slots_35_io_request & (|_GEN_626) & ~_GEN_615 | _GEN_624;
  wire [9:0]  _can_allocate_T_142 = _slots_35_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_631 = _slots_35_io_request & ~_GEN_630 & (|_can_allocate_T_142);
  wire        _GEN_632 = _GEN_631 & ~_GEN_619;
  wire        _GEN_633 = _GEN_631 | _GEN_619;
  wire        _GEN_634 = _slots_35_io_request & ~(_slots_35_io_request & (|_can_allocate_T_142) & ~_GEN_619 | _GEN_630) & (|(_slots_35_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_635 = _GEN_634 & ~_GEN_622;
  assign issue_slots_35_grant = _GEN_635 | _GEN_632 | _GEN_628 | _GEN_624;
  wire        _GEN_636 = _GEN_634 | _GEN_622;
  wire        _GEN_637 = _slots_36_io_request & (|(_slots_36_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_638 = _GEN_637 & ~_GEN_625;
  wire        _GEN_639 = _GEN_637 | _GEN_625;
  wire [1:0]  _GEN_640 = {_slots_36_io_uop_fu_code[5], _slots_36_io_uop_fu_code[0]};
  wire        _GEN_641 = _slots_36_io_request & ~_GEN_638 & (|_GEN_640);
  wire        _GEN_642 = _GEN_641 & ~_GEN_629;
  wire        _GEN_643 = _GEN_641 | _GEN_629;
  wire        _GEN_644 = _slots_36_io_request & (|_GEN_640) & ~_GEN_629 | _GEN_638;
  wire [9:0]  _can_allocate_T_146 = _slots_36_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_645 = _slots_36_io_request & ~_GEN_644 & (|_can_allocate_T_146);
  wire        _GEN_646 = _GEN_645 & ~_GEN_633;
  wire        _GEN_647 = _GEN_645 | _GEN_633;
  wire        _GEN_648 = _slots_36_io_request & ~(_slots_36_io_request & (|_can_allocate_T_146) & ~_GEN_633 | _GEN_644) & (|(_slots_36_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_649 = _GEN_648 & ~_GEN_636;
  assign issue_slots_36_grant = _GEN_649 | _GEN_646 | _GEN_642 | _GEN_638;
  wire        _GEN_650 = _GEN_648 | _GEN_636;
  wire        _GEN_651 = _slots_37_io_request & (|(_slots_37_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_652 = _GEN_651 & ~_GEN_639;
  wire        _GEN_653 = _GEN_651 | _GEN_639;
  wire [1:0]  _GEN_654 = {_slots_37_io_uop_fu_code[5], _slots_37_io_uop_fu_code[0]};
  wire        _GEN_655 = _slots_37_io_request & ~_GEN_652 & (|_GEN_654);
  wire        _GEN_656 = _GEN_655 & ~_GEN_643;
  wire        _GEN_657 = _GEN_655 | _GEN_643;
  wire        _GEN_658 = _slots_37_io_request & (|_GEN_654) & ~_GEN_643 | _GEN_652;
  wire [9:0]  _can_allocate_T_150 = _slots_37_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_659 = _slots_37_io_request & ~_GEN_658 & (|_can_allocate_T_150);
  wire        _GEN_660 = _GEN_659 & ~_GEN_647;
  wire        _GEN_661 = _GEN_659 | _GEN_647;
  wire        _GEN_662 = _slots_37_io_request & ~(_slots_37_io_request & (|_can_allocate_T_150) & ~_GEN_647 | _GEN_658) & (|(_slots_37_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_663 = _GEN_662 & ~_GEN_650;
  assign issue_slots_37_grant = _GEN_663 | _GEN_660 | _GEN_656 | _GEN_652;
  wire        _GEN_664 = _GEN_662 | _GEN_650;
  wire        _GEN_665 = _slots_38_io_request & (|(_slots_38_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_666 = _GEN_665 & ~_GEN_653;
  wire [1:0]  _GEN_667 = {_slots_38_io_uop_fu_code[5], _slots_38_io_uop_fu_code[0]};
  wire        _GEN_668 = _slots_38_io_request & ~_GEN_666 & (|_GEN_667);
  wire        _GEN_669 = _GEN_668 & ~_GEN_657;
  wire        _GEN_670 = _GEN_668 | _GEN_657;
  wire        _GEN_671 = _slots_38_io_request & (|_GEN_667) & ~_GEN_657 | _GEN_666;
  wire [9:0]  _can_allocate_T_154 = _slots_38_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_672 = _slots_38_io_request & ~_GEN_671 & (|_can_allocate_T_154);
  wire        _GEN_673 = _GEN_672 & ~_GEN_661;
  wire        _GEN_674 = _GEN_672 | _GEN_661;
  wire        _GEN_675 = _slots_38_io_request & ~(_slots_38_io_request & (|_can_allocate_T_154) & ~_GEN_661 | _GEN_671) & (|(_slots_38_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_676 = _GEN_675 & ~_GEN_664;
  assign issue_slots_38_grant = _GEN_676 | _GEN_673 | _GEN_669 | _GEN_666;
  wire        _GEN_677 = _slots_39_io_request & (|(_slots_39_io_uop_fu_code & io_fu_types_0)) & ~(_GEN_665 | _GEN_653);
  wire [1:0]  _GEN_678 = {_slots_39_io_uop_fu_code[5], _slots_39_io_uop_fu_code[0]};
  wire        _GEN_679 = _slots_39_io_request & ~_GEN_677 & (|_GEN_678) & ~_GEN_670;
  wire        _GEN_680 = _slots_39_io_request & (|_GEN_678) & ~_GEN_670 | _GEN_677;
  wire [9:0]  _can_allocate_T_158 = _slots_39_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_681 = _slots_39_io_request & ~_GEN_680 & (|_can_allocate_T_158) & ~_GEN_674;
  wire        _GEN_682 = _slots_39_io_request & ~(_slots_39_io_request & (|_can_allocate_T_158) & ~_GEN_674 | _GEN_680) & (|(_slots_39_io_uop_fu_code & io_fu_types_3)) & ~(_GEN_675 | _GEN_664);
  assign issue_slots_39_grant = _GEN_682 | _GEN_681 | _GEN_679 | _GEN_677;
  wire [5:0]  num_available =
    {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, ~_slots_0_io_will_be_valid & ~issue_slots_0_in_uop_valid} + {1'h0, (~_slots_1_io_will_be_valid | ~_slots_0_io_valid) & ~issue_slots_1_in_uop_valid}} + {1'h0, {1'h0, (~_slots_2_io_will_be_valid | (|_next_1_1to0)) & ~issue_slots_2_in_uop_valid} + {1'h0, (~_slots_3_io_will_be_valid | (|next_2)) & ~issue_slots_3_in_uop_valid} + {1'h0, (~_slots_4_io_will_be_valid | (|next_3)) & ~issue_slots_4_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_5_io_will_be_valid | (|next_4)) & ~issue_slots_5_in_uop_valid} + {1'h0, (~_slots_6_io_will_be_valid | (|next_5)) & ~issue_slots_6_in_uop_valid}} + {1'h0, {1'h0, (~_slots_7_io_will_be_valid | (|next_6)) & ~issue_slots_7_in_uop_valid} + {1'h0, (~_slots_8_io_will_be_valid | (|next_7)) & ~issue_slots_8_in_uop_valid} + {1'h0, (~_slots_9_io_will_be_valid | (|next_8)) & ~issue_slots_9_in_uop_valid}}}} + {1'h0, {1'h0, {1'h0, {1'h0, (~_slots_10_io_will_be_valid | (|next_9)) & ~issue_slots_10_in_uop_valid} + {1'h0, (~_slots_11_io_will_be_valid | (|next_10)) & ~issue_slots_11_in_uop_valid}} + {1'h0, {1'h0, (~_slots_12_io_will_be_valid | (|next_11)) & ~issue_slots_12_in_uop_valid} + {1'h0, (~_slots_13_io_will_be_valid | (|next_12)) & ~issue_slots_13_in_uop_valid} + {1'h0, (~_slots_14_io_will_be_valid | (|next_13)) & ~issue_slots_14_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_15_io_will_be_valid | (|next_14)) & ~issue_slots_15_in_uop_valid} + {1'h0, (~_slots_16_io_will_be_valid | (|next_15)) & ~issue_slots_16_in_uop_valid}} + {1'h0, {1'h0, (~_slots_17_io_will_be_valid | (|next_16)) & ~issue_slots_17_in_uop_valid} + {1'h0, (~_slots_18_io_will_be_valid | (|next_17)) & ~issue_slots_18_in_uop_valid} + {1'h0, (~_slots_19_io_will_be_valid | (|next_18)) & ~issue_slots_19_in_uop_valid}}}}}
    + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, (~_slots_20_io_will_be_valid | (|next_19)) & ~issue_slots_20_in_uop_valid} + {1'h0, (~_slots_21_io_will_be_valid | (|next_20)) & ~issue_slots_21_in_uop_valid}} + {1'h0, {1'h0, (~_slots_22_io_will_be_valid | (|next_21)) & ~issue_slots_22_in_uop_valid} + {1'h0, (~_slots_23_io_will_be_valid | (|next_22)) & ~issue_slots_23_in_uop_valid} + {1'h0, (~_slots_24_io_will_be_valid | (|next_23)) & ~issue_slots_24_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_25_io_will_be_valid | (|next_24)) & ~issue_slots_25_in_uop_valid} + {1'h0, (~_slots_26_io_will_be_valid | (|next_25)) & ~issue_slots_26_in_uop_valid}} + {1'h0, {1'h0, (~_slots_27_io_will_be_valid | (|next_26)) & ~issue_slots_27_in_uop_valid} + {1'h0, (~_slots_28_io_will_be_valid | (|next_27)) & ~issue_slots_28_in_uop_valid} + {1'h0, (~_slots_29_io_will_be_valid | (|next_28)) & ~issue_slots_29_in_uop_valid}}}} + {1'h0, {1'h0, {1'h0, {1'h0, (~_slots_30_io_will_be_valid | (|next_29)) & ~issue_slots_30_in_uop_valid} + {1'h0, (~_slots_31_io_will_be_valid | (|next_30)) & ~issue_slots_31_in_uop_valid}} + {1'h0, {1'h0, (~_slots_32_io_will_be_valid | (|next_31)) & ~issue_slots_32_in_uop_valid} + {1'h0, (~_slots_33_io_will_be_valid | (|next_32)) & ~issue_slots_33_in_uop_valid} + {1'h0, (~_slots_34_io_will_be_valid | (|next_33)) & ~issue_slots_34_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_35_io_will_be_valid | (|next_34)) & ~issue_slots_35_in_uop_valid} + {1'h0, (~_slots_36_io_will_be_valid | (|next_35)) & ~issue_slots_36_in_uop_valid}} + {1'h0, {1'h0, (~_slots_37_io_will_be_valid | (|next_36)) & ~issue_slots_37_in_uop_valid} + {1'h0, (~_slots_38_io_will_be_valid | (|next_37)) & ~issue_slots_38_in_uop_valid} + {1'h0, (~_slots_39_io_will_be_valid | (|next_38)) & ~issue_slots_39_in_uop_valid}}}}};
  always @(posedge clock) begin
    io_dis_uops_0_ready_REG <= |num_available;
    io_dis_uops_1_ready_REG <= |(num_available[5:1]);
    io_dis_uops_2_ready_REG <= num_available > 6'h2;
    io_dis_uops_3_ready_REG <= |(num_available[5:2]);
  end // always @(posedge)
  IssueSlot_32 slots_0 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_0_io_valid),
    .io_will_be_valid               (_slots_0_io_will_be_valid),
    .io_request                     (_slots_0_io_request),
    .io_grant                       (issue_slots_0_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (1'h0),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_0_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_21 ? _slots_4_io_out_uop_uopc : _GEN_20 ? _slots_3_io_out_uop_uopc : _GEN_19 ? _slots_2_io_out_uop_uopc : _slots_1_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_21 ? _slots_4_io_out_uop_inst : _GEN_20 ? _slots_3_io_out_uop_inst : _GEN_19 ? _slots_2_io_out_uop_inst : _slots_1_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_21 ? _slots_4_io_out_uop_debug_inst : _GEN_20 ? _slots_3_io_out_uop_debug_inst : _GEN_19 ? _slots_2_io_out_uop_debug_inst : _slots_1_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_21 ? _slots_4_io_out_uop_is_rvc : _GEN_20 ? _slots_3_io_out_uop_is_rvc : _GEN_19 ? _slots_2_io_out_uop_is_rvc : _slots_1_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_21 ? _slots_4_io_out_uop_debug_pc : _GEN_20 ? _slots_3_io_out_uop_debug_pc : _GEN_19 ? _slots_2_io_out_uop_debug_pc : _slots_1_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_21 ? _slots_4_io_out_uop_iq_type : _GEN_20 ? _slots_3_io_out_uop_iq_type : _GEN_19 ? _slots_2_io_out_uop_iq_type : _slots_1_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_21 ? _slots_4_io_out_uop_fu_code : _GEN_20 ? _slots_3_io_out_uop_fu_code : _GEN_19 ? _slots_2_io_out_uop_fu_code : _slots_1_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_21 ? _slots_4_io_out_uop_iw_state : _GEN_20 ? _slots_3_io_out_uop_iw_state : _GEN_19 ? _slots_2_io_out_uop_iw_state : _slots_1_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_21 ? _slots_4_io_out_uop_iw_p1_poisoned : _GEN_20 ? _slots_3_io_out_uop_iw_p1_poisoned : _GEN_19 ? _slots_2_io_out_uop_iw_p1_poisoned : _slots_1_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_21 ? _slots_4_io_out_uop_iw_p2_poisoned : _GEN_20 ? _slots_3_io_out_uop_iw_p2_poisoned : _GEN_19 ? _slots_2_io_out_uop_iw_p2_poisoned : _slots_1_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_21 ? _slots_4_io_out_uop_is_br : _GEN_20 ? _slots_3_io_out_uop_is_br : _GEN_19 ? _slots_2_io_out_uop_is_br : _slots_1_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_21 ? _slots_4_io_out_uop_is_jalr : _GEN_20 ? _slots_3_io_out_uop_is_jalr : _GEN_19 ? _slots_2_io_out_uop_is_jalr : _slots_1_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_21 ? _slots_4_io_out_uop_is_jal : _GEN_20 ? _slots_3_io_out_uop_is_jal : _GEN_19 ? _slots_2_io_out_uop_is_jal : _slots_1_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_21 ? _slots_4_io_out_uop_is_sfb : _GEN_20 ? _slots_3_io_out_uop_is_sfb : _GEN_19 ? _slots_2_io_out_uop_is_sfb : _slots_1_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_21 ? _slots_4_io_out_uop_br_mask : _GEN_20 ? _slots_3_io_out_uop_br_mask : _GEN_19 ? _slots_2_io_out_uop_br_mask : _slots_1_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_21 ? _slots_4_io_out_uop_br_tag : _GEN_20 ? _slots_3_io_out_uop_br_tag : _GEN_19 ? _slots_2_io_out_uop_br_tag : _slots_1_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_21 ? _slots_4_io_out_uop_ftq_idx : _GEN_20 ? _slots_3_io_out_uop_ftq_idx : _GEN_19 ? _slots_2_io_out_uop_ftq_idx : _slots_1_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_21 ? _slots_4_io_out_uop_edge_inst : _GEN_20 ? _slots_3_io_out_uop_edge_inst : _GEN_19 ? _slots_2_io_out_uop_edge_inst : _slots_1_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_21 ? _slots_4_io_out_uop_pc_lob : _GEN_20 ? _slots_3_io_out_uop_pc_lob : _GEN_19 ? _slots_2_io_out_uop_pc_lob : _slots_1_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_21 ? _slots_4_io_out_uop_taken : _GEN_20 ? _slots_3_io_out_uop_taken : _GEN_19 ? _slots_2_io_out_uop_taken : _slots_1_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_21 ? _slots_4_io_out_uop_imm_packed : _GEN_20 ? _slots_3_io_out_uop_imm_packed : _GEN_19 ? _slots_2_io_out_uop_imm_packed : _slots_1_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_21 ? _slots_4_io_out_uop_csr_addr : _GEN_20 ? _slots_3_io_out_uop_csr_addr : _GEN_19 ? _slots_2_io_out_uop_csr_addr : _slots_1_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_21 ? _slots_4_io_out_uop_rob_idx : _GEN_20 ? _slots_3_io_out_uop_rob_idx : _GEN_19 ? _slots_2_io_out_uop_rob_idx : _slots_1_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_21 ? _slots_4_io_out_uop_ldq_idx : _GEN_20 ? _slots_3_io_out_uop_ldq_idx : _GEN_19 ? _slots_2_io_out_uop_ldq_idx : _slots_1_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_21 ? _slots_4_io_out_uop_stq_idx : _GEN_20 ? _slots_3_io_out_uop_stq_idx : _GEN_19 ? _slots_2_io_out_uop_stq_idx : _slots_1_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_21 ? _slots_4_io_out_uop_rxq_idx : _GEN_20 ? _slots_3_io_out_uop_rxq_idx : _GEN_19 ? _slots_2_io_out_uop_rxq_idx : _slots_1_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_21 ? _slots_4_io_out_uop_pdst : _GEN_20 ? _slots_3_io_out_uop_pdst : _GEN_19 ? _slots_2_io_out_uop_pdst : _slots_1_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_21 ? _slots_4_io_out_uop_prs1 : _GEN_20 ? _slots_3_io_out_uop_prs1 : _GEN_19 ? _slots_2_io_out_uop_prs1 : _slots_1_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_21 ? _slots_4_io_out_uop_prs2 : _GEN_20 ? _slots_3_io_out_uop_prs2 : _GEN_19 ? _slots_2_io_out_uop_prs2 : _slots_1_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_21 ? _slots_4_io_out_uop_prs3 : _GEN_20 ? _slots_3_io_out_uop_prs3 : _GEN_19 ? _slots_2_io_out_uop_prs3 : _slots_1_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_21 ? _slots_4_io_out_uop_ppred : _GEN_20 ? _slots_3_io_out_uop_ppred : _GEN_19 ? _slots_2_io_out_uop_ppred : _slots_1_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_21 ? _slots_4_io_out_uop_prs1_busy : _GEN_20 ? _slots_3_io_out_uop_prs1_busy : _GEN_19 ? _slots_2_io_out_uop_prs1_busy : _slots_1_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_21 ? _slots_4_io_out_uop_prs2_busy : _GEN_20 ? _slots_3_io_out_uop_prs2_busy : _GEN_19 ? _slots_2_io_out_uop_prs2_busy : _slots_1_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_21 ? _slots_4_io_out_uop_prs3_busy : _GEN_20 ? _slots_3_io_out_uop_prs3_busy : _GEN_19 ? _slots_2_io_out_uop_prs3_busy : _slots_1_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_21 ? _slots_4_io_out_uop_ppred_busy : _GEN_20 ? _slots_3_io_out_uop_ppred_busy : _GEN_19 ? _slots_2_io_out_uop_ppred_busy : _slots_1_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_21 ? _slots_4_io_out_uop_stale_pdst : _GEN_20 ? _slots_3_io_out_uop_stale_pdst : _GEN_19 ? _slots_2_io_out_uop_stale_pdst : _slots_1_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_21 ? _slots_4_io_out_uop_exception : _GEN_20 ? _slots_3_io_out_uop_exception : _GEN_19 ? _slots_2_io_out_uop_exception : _slots_1_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_21 ? _slots_4_io_out_uop_exc_cause : _GEN_20 ? _slots_3_io_out_uop_exc_cause : _GEN_19 ? _slots_2_io_out_uop_exc_cause : _slots_1_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_21 ? _slots_4_io_out_uop_bypassable : _GEN_20 ? _slots_3_io_out_uop_bypassable : _GEN_19 ? _slots_2_io_out_uop_bypassable : _slots_1_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_21 ? _slots_4_io_out_uop_mem_cmd : _GEN_20 ? _slots_3_io_out_uop_mem_cmd : _GEN_19 ? _slots_2_io_out_uop_mem_cmd : _slots_1_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_21 ? _slots_4_io_out_uop_mem_size : _GEN_20 ? _slots_3_io_out_uop_mem_size : _GEN_19 ? _slots_2_io_out_uop_mem_size : _slots_1_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_21 ? _slots_4_io_out_uop_mem_signed : _GEN_20 ? _slots_3_io_out_uop_mem_signed : _GEN_19 ? _slots_2_io_out_uop_mem_signed : _slots_1_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_21 ? _slots_4_io_out_uop_is_fence : _GEN_20 ? _slots_3_io_out_uop_is_fence : _GEN_19 ? _slots_2_io_out_uop_is_fence : _slots_1_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_21 ? _slots_4_io_out_uop_is_fencei : _GEN_20 ? _slots_3_io_out_uop_is_fencei : _GEN_19 ? _slots_2_io_out_uop_is_fencei : _slots_1_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_21 ? _slots_4_io_out_uop_is_amo : _GEN_20 ? _slots_3_io_out_uop_is_amo : _GEN_19 ? _slots_2_io_out_uop_is_amo : _slots_1_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_21 ? _slots_4_io_out_uop_uses_ldq : _GEN_20 ? _slots_3_io_out_uop_uses_ldq : _GEN_19 ? _slots_2_io_out_uop_uses_ldq : _slots_1_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_21 ? _slots_4_io_out_uop_uses_stq : _GEN_20 ? _slots_3_io_out_uop_uses_stq : _GEN_19 ? _slots_2_io_out_uop_uses_stq : _slots_1_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_21 ? _slots_4_io_out_uop_is_sys_pc2epc : _GEN_20 ? _slots_3_io_out_uop_is_sys_pc2epc : _GEN_19 ? _slots_2_io_out_uop_is_sys_pc2epc : _slots_1_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_21 ? _slots_4_io_out_uop_is_unique : _GEN_20 ? _slots_3_io_out_uop_is_unique : _GEN_19 ? _slots_2_io_out_uop_is_unique : _slots_1_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_21 ? _slots_4_io_out_uop_flush_on_commit : _GEN_20 ? _slots_3_io_out_uop_flush_on_commit : _GEN_19 ? _slots_2_io_out_uop_flush_on_commit : _slots_1_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_21 ? _slots_4_io_out_uop_ldst_is_rs1 : _GEN_20 ? _slots_3_io_out_uop_ldst_is_rs1 : _GEN_19 ? _slots_2_io_out_uop_ldst_is_rs1 : _slots_1_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_21 ? _slots_4_io_out_uop_ldst : _GEN_20 ? _slots_3_io_out_uop_ldst : _GEN_19 ? _slots_2_io_out_uop_ldst : _slots_1_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_21 ? _slots_4_io_out_uop_lrs1 : _GEN_20 ? _slots_3_io_out_uop_lrs1 : _GEN_19 ? _slots_2_io_out_uop_lrs1 : _slots_1_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_21 ? _slots_4_io_out_uop_lrs2 : _GEN_20 ? _slots_3_io_out_uop_lrs2 : _GEN_19 ? _slots_2_io_out_uop_lrs2 : _slots_1_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_21 ? _slots_4_io_out_uop_lrs3 : _GEN_20 ? _slots_3_io_out_uop_lrs3 : _GEN_19 ? _slots_2_io_out_uop_lrs3 : _slots_1_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_21 ? _slots_4_io_out_uop_ldst_val : _GEN_20 ? _slots_3_io_out_uop_ldst_val : _GEN_19 ? _slots_2_io_out_uop_ldst_val : _slots_1_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_21 ? _slots_4_io_out_uop_dst_rtype : _GEN_20 ? _slots_3_io_out_uop_dst_rtype : _GEN_19 ? _slots_2_io_out_uop_dst_rtype : _slots_1_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_21 ? _slots_4_io_out_uop_lrs1_rtype : _GEN_20 ? _slots_3_io_out_uop_lrs1_rtype : _GEN_19 ? _slots_2_io_out_uop_lrs1_rtype : _slots_1_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_21 ? _slots_4_io_out_uop_lrs2_rtype : _GEN_20 ? _slots_3_io_out_uop_lrs2_rtype : _GEN_19 ? _slots_2_io_out_uop_lrs2_rtype : _slots_1_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_21 ? _slots_4_io_out_uop_frs3_en : _GEN_20 ? _slots_3_io_out_uop_frs3_en : _GEN_19 ? _slots_2_io_out_uop_frs3_en : _slots_1_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_21 ? _slots_4_io_out_uop_fp_val : _GEN_20 ? _slots_3_io_out_uop_fp_val : _GEN_19 ? _slots_2_io_out_uop_fp_val : _slots_1_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_21 ? _slots_4_io_out_uop_fp_single : _GEN_20 ? _slots_3_io_out_uop_fp_single : _GEN_19 ? _slots_2_io_out_uop_fp_single : _slots_1_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_21 ? _slots_4_io_out_uop_xcpt_pf_if : _GEN_20 ? _slots_3_io_out_uop_xcpt_pf_if : _GEN_19 ? _slots_2_io_out_uop_xcpt_pf_if : _slots_1_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_21 ? _slots_4_io_out_uop_xcpt_ae_if : _GEN_20 ? _slots_3_io_out_uop_xcpt_ae_if : _GEN_19 ? _slots_2_io_out_uop_xcpt_ae_if : _slots_1_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_21 ? _slots_4_io_out_uop_xcpt_ma_if : _GEN_20 ? _slots_3_io_out_uop_xcpt_ma_if : _GEN_19 ? _slots_2_io_out_uop_xcpt_ma_if : _slots_1_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_21 ? _slots_4_io_out_uop_bp_debug_if : _GEN_20 ? _slots_3_io_out_uop_bp_debug_if : _GEN_19 ? _slots_2_io_out_uop_bp_debug_if : _slots_1_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_21 ? _slots_4_io_out_uop_bp_xcpt_if : _GEN_20 ? _slots_3_io_out_uop_bp_xcpt_if : _GEN_19 ? _slots_2_io_out_uop_bp_xcpt_if : _slots_1_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_21 ? _slots_4_io_out_uop_debug_fsrc : _GEN_20 ? _slots_3_io_out_uop_debug_fsrc : _GEN_19 ? _slots_2_io_out_uop_debug_fsrc : _slots_1_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_21 ? _slots_4_io_out_uop_debug_tsrc : _GEN_20 ? _slots_3_io_out_uop_debug_tsrc : _GEN_19 ? _slots_2_io_out_uop_debug_tsrc : _slots_1_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (/* unused */),
    .io_out_uop_inst                (/* unused */),
    .io_out_uop_debug_inst          (/* unused */),
    .io_out_uop_is_rvc              (/* unused */),
    .io_out_uop_debug_pc            (/* unused */),
    .io_out_uop_iq_type             (/* unused */),
    .io_out_uop_fu_code             (/* unused */),
    .io_out_uop_iw_state            (/* unused */),
    .io_out_uop_iw_p1_poisoned      (/* unused */),
    .io_out_uop_iw_p2_poisoned      (/* unused */),
    .io_out_uop_is_br               (/* unused */),
    .io_out_uop_is_jalr             (/* unused */),
    .io_out_uop_is_jal              (/* unused */),
    .io_out_uop_is_sfb              (/* unused */),
    .io_out_uop_br_mask             (/* unused */),
    .io_out_uop_br_tag              (/* unused */),
    .io_out_uop_ftq_idx             (/* unused */),
    .io_out_uop_edge_inst           (/* unused */),
    .io_out_uop_pc_lob              (/* unused */),
    .io_out_uop_taken               (/* unused */),
    .io_out_uop_imm_packed          (/* unused */),
    .io_out_uop_csr_addr            (/* unused */),
    .io_out_uop_rob_idx             (/* unused */),
    .io_out_uop_ldq_idx             (/* unused */),
    .io_out_uop_stq_idx             (/* unused */),
    .io_out_uop_rxq_idx             (/* unused */),
    .io_out_uop_pdst                (/* unused */),
    .io_out_uop_prs1                (/* unused */),
    .io_out_uop_prs2                (/* unused */),
    .io_out_uop_prs3                (/* unused */),
    .io_out_uop_ppred               (/* unused */),
    .io_out_uop_prs1_busy           (/* unused */),
    .io_out_uop_prs2_busy           (/* unused */),
    .io_out_uop_prs3_busy           (/* unused */),
    .io_out_uop_ppred_busy          (/* unused */),
    .io_out_uop_stale_pdst          (/* unused */),
    .io_out_uop_exception           (/* unused */),
    .io_out_uop_exc_cause           (/* unused */),
    .io_out_uop_bypassable          (/* unused */),
    .io_out_uop_mem_cmd             (/* unused */),
    .io_out_uop_mem_size            (/* unused */),
    .io_out_uop_mem_signed          (/* unused */),
    .io_out_uop_is_fence            (/* unused */),
    .io_out_uop_is_fencei           (/* unused */),
    .io_out_uop_is_amo              (/* unused */),
    .io_out_uop_uses_ldq            (/* unused */),
    .io_out_uop_uses_stq            (/* unused */),
    .io_out_uop_is_sys_pc2epc       (/* unused */),
    .io_out_uop_is_unique           (/* unused */),
    .io_out_uop_flush_on_commit     (/* unused */),
    .io_out_uop_ldst_is_rs1         (/* unused */),
    .io_out_uop_ldst                (/* unused */),
    .io_out_uop_lrs1                (/* unused */),
    .io_out_uop_lrs2                (/* unused */),
    .io_out_uop_lrs3                (/* unused */),
    .io_out_uop_ldst_val            (/* unused */),
    .io_out_uop_dst_rtype           (/* unused */),
    .io_out_uop_lrs1_rtype          (/* unused */),
    .io_out_uop_lrs2_rtype          (/* unused */),
    .io_out_uop_frs3_en             (/* unused */),
    .io_out_uop_fp_val              (/* unused */),
    .io_out_uop_fp_single           (/* unused */),
    .io_out_uop_xcpt_pf_if          (/* unused */),
    .io_out_uop_xcpt_ae_if          (/* unused */),
    .io_out_uop_xcpt_ma_if          (/* unused */),
    .io_out_uop_bp_debug_if         (/* unused */),
    .io_out_uop_bp_xcpt_if          (/* unused */),
    .io_out_uop_debug_fsrc          (/* unused */),
    .io_out_uop_debug_tsrc          (/* unused */),
    .io_uop_uopc                    (_slots_0_io_uop_uopc),
    .io_uop_inst                    (_slots_0_io_uop_inst),
    .io_uop_debug_inst              (_slots_0_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_0_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_0_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_0_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_0_io_uop_fu_code),
    .io_uop_iw_state                (_slots_0_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_0_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_0_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_0_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_0_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_0_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_0_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_0_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_0_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_0_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_0_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_0_io_uop_pc_lob),
    .io_uop_taken                   (_slots_0_io_uop_taken),
    .io_uop_imm_packed              (_slots_0_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_0_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_0_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_0_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_0_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_0_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_0_io_uop_pdst),
    .io_uop_prs1                    (_slots_0_io_uop_prs1),
    .io_uop_prs2                    (_slots_0_io_uop_prs2),
    .io_uop_prs3                    (_slots_0_io_uop_prs3),
    .io_uop_ppred                   (_slots_0_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_0_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_0_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_0_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_0_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_0_io_uop_stale_pdst),
    .io_uop_exception               (_slots_0_io_uop_exception),
    .io_uop_exc_cause               (_slots_0_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_0_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_0_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_0_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_0_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_0_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_0_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_0_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_0_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_0_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_0_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_0_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_0_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_0_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_0_io_uop_ldst),
    .io_uop_lrs1                    (_slots_0_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_0_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_0_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_0_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_0_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_0_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_0_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_0_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_0_io_uop_fp_val),
    .io_uop_fp_single               (_slots_0_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_0_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_0_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_0_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_0_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_0_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_0_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_0_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_1 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_1_io_valid),
    .io_will_be_valid               (_slots_1_io_will_be_valid),
    .io_request                     (_slots_1_io_request),
    .io_grant                       (issue_slots_1_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (~_slots_0_io_valid),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_1_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_24 ? _slots_5_io_out_uop_uopc : _GEN_23 ? _slots_4_io_out_uop_uopc : _GEN_22 ? _slots_3_io_out_uop_uopc : _slots_2_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_24 ? _slots_5_io_out_uop_inst : _GEN_23 ? _slots_4_io_out_uop_inst : _GEN_22 ? _slots_3_io_out_uop_inst : _slots_2_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_24 ? _slots_5_io_out_uop_debug_inst : _GEN_23 ? _slots_4_io_out_uop_debug_inst : _GEN_22 ? _slots_3_io_out_uop_debug_inst : _slots_2_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_24 ? _slots_5_io_out_uop_is_rvc : _GEN_23 ? _slots_4_io_out_uop_is_rvc : _GEN_22 ? _slots_3_io_out_uop_is_rvc : _slots_2_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_24 ? _slots_5_io_out_uop_debug_pc : _GEN_23 ? _slots_4_io_out_uop_debug_pc : _GEN_22 ? _slots_3_io_out_uop_debug_pc : _slots_2_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_24 ? _slots_5_io_out_uop_iq_type : _GEN_23 ? _slots_4_io_out_uop_iq_type : _GEN_22 ? _slots_3_io_out_uop_iq_type : _slots_2_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_24 ? _slots_5_io_out_uop_fu_code : _GEN_23 ? _slots_4_io_out_uop_fu_code : _GEN_22 ? _slots_3_io_out_uop_fu_code : _slots_2_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_24 ? _slots_5_io_out_uop_iw_state : _GEN_23 ? _slots_4_io_out_uop_iw_state : _GEN_22 ? _slots_3_io_out_uop_iw_state : _slots_2_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_24 ? _slots_5_io_out_uop_iw_p1_poisoned : _GEN_23 ? _slots_4_io_out_uop_iw_p1_poisoned : _GEN_22 ? _slots_3_io_out_uop_iw_p1_poisoned : _slots_2_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_24 ? _slots_5_io_out_uop_iw_p2_poisoned : _GEN_23 ? _slots_4_io_out_uop_iw_p2_poisoned : _GEN_22 ? _slots_3_io_out_uop_iw_p2_poisoned : _slots_2_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_24 ? _slots_5_io_out_uop_is_br : _GEN_23 ? _slots_4_io_out_uop_is_br : _GEN_22 ? _slots_3_io_out_uop_is_br : _slots_2_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_24 ? _slots_5_io_out_uop_is_jalr : _GEN_23 ? _slots_4_io_out_uop_is_jalr : _GEN_22 ? _slots_3_io_out_uop_is_jalr : _slots_2_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_24 ? _slots_5_io_out_uop_is_jal : _GEN_23 ? _slots_4_io_out_uop_is_jal : _GEN_22 ? _slots_3_io_out_uop_is_jal : _slots_2_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_24 ? _slots_5_io_out_uop_is_sfb : _GEN_23 ? _slots_4_io_out_uop_is_sfb : _GEN_22 ? _slots_3_io_out_uop_is_sfb : _slots_2_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_24 ? _slots_5_io_out_uop_br_mask : _GEN_23 ? _slots_4_io_out_uop_br_mask : _GEN_22 ? _slots_3_io_out_uop_br_mask : _slots_2_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_24 ? _slots_5_io_out_uop_br_tag : _GEN_23 ? _slots_4_io_out_uop_br_tag : _GEN_22 ? _slots_3_io_out_uop_br_tag : _slots_2_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_24 ? _slots_5_io_out_uop_ftq_idx : _GEN_23 ? _slots_4_io_out_uop_ftq_idx : _GEN_22 ? _slots_3_io_out_uop_ftq_idx : _slots_2_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_24 ? _slots_5_io_out_uop_edge_inst : _GEN_23 ? _slots_4_io_out_uop_edge_inst : _GEN_22 ? _slots_3_io_out_uop_edge_inst : _slots_2_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_24 ? _slots_5_io_out_uop_pc_lob : _GEN_23 ? _slots_4_io_out_uop_pc_lob : _GEN_22 ? _slots_3_io_out_uop_pc_lob : _slots_2_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_24 ? _slots_5_io_out_uop_taken : _GEN_23 ? _slots_4_io_out_uop_taken : _GEN_22 ? _slots_3_io_out_uop_taken : _slots_2_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_24 ? _slots_5_io_out_uop_imm_packed : _GEN_23 ? _slots_4_io_out_uop_imm_packed : _GEN_22 ? _slots_3_io_out_uop_imm_packed : _slots_2_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_24 ? _slots_5_io_out_uop_csr_addr : _GEN_23 ? _slots_4_io_out_uop_csr_addr : _GEN_22 ? _slots_3_io_out_uop_csr_addr : _slots_2_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_24 ? _slots_5_io_out_uop_rob_idx : _GEN_23 ? _slots_4_io_out_uop_rob_idx : _GEN_22 ? _slots_3_io_out_uop_rob_idx : _slots_2_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_24 ? _slots_5_io_out_uop_ldq_idx : _GEN_23 ? _slots_4_io_out_uop_ldq_idx : _GEN_22 ? _slots_3_io_out_uop_ldq_idx : _slots_2_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_24 ? _slots_5_io_out_uop_stq_idx : _GEN_23 ? _slots_4_io_out_uop_stq_idx : _GEN_22 ? _slots_3_io_out_uop_stq_idx : _slots_2_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_24 ? _slots_5_io_out_uop_rxq_idx : _GEN_23 ? _slots_4_io_out_uop_rxq_idx : _GEN_22 ? _slots_3_io_out_uop_rxq_idx : _slots_2_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_24 ? _slots_5_io_out_uop_pdst : _GEN_23 ? _slots_4_io_out_uop_pdst : _GEN_22 ? _slots_3_io_out_uop_pdst : _slots_2_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_24 ? _slots_5_io_out_uop_prs1 : _GEN_23 ? _slots_4_io_out_uop_prs1 : _GEN_22 ? _slots_3_io_out_uop_prs1 : _slots_2_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_24 ? _slots_5_io_out_uop_prs2 : _GEN_23 ? _slots_4_io_out_uop_prs2 : _GEN_22 ? _slots_3_io_out_uop_prs2 : _slots_2_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_24 ? _slots_5_io_out_uop_prs3 : _GEN_23 ? _slots_4_io_out_uop_prs3 : _GEN_22 ? _slots_3_io_out_uop_prs3 : _slots_2_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_24 ? _slots_5_io_out_uop_ppred : _GEN_23 ? _slots_4_io_out_uop_ppred : _GEN_22 ? _slots_3_io_out_uop_ppred : _slots_2_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_24 ? _slots_5_io_out_uop_prs1_busy : _GEN_23 ? _slots_4_io_out_uop_prs1_busy : _GEN_22 ? _slots_3_io_out_uop_prs1_busy : _slots_2_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_24 ? _slots_5_io_out_uop_prs2_busy : _GEN_23 ? _slots_4_io_out_uop_prs2_busy : _GEN_22 ? _slots_3_io_out_uop_prs2_busy : _slots_2_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_24 ? _slots_5_io_out_uop_prs3_busy : _GEN_23 ? _slots_4_io_out_uop_prs3_busy : _GEN_22 ? _slots_3_io_out_uop_prs3_busy : _slots_2_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_24 ? _slots_5_io_out_uop_ppred_busy : _GEN_23 ? _slots_4_io_out_uop_ppred_busy : _GEN_22 ? _slots_3_io_out_uop_ppred_busy : _slots_2_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_24 ? _slots_5_io_out_uop_stale_pdst : _GEN_23 ? _slots_4_io_out_uop_stale_pdst : _GEN_22 ? _slots_3_io_out_uop_stale_pdst : _slots_2_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_24 ? _slots_5_io_out_uop_exception : _GEN_23 ? _slots_4_io_out_uop_exception : _GEN_22 ? _slots_3_io_out_uop_exception : _slots_2_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_24 ? _slots_5_io_out_uop_exc_cause : _GEN_23 ? _slots_4_io_out_uop_exc_cause : _GEN_22 ? _slots_3_io_out_uop_exc_cause : _slots_2_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_24 ? _slots_5_io_out_uop_bypassable : _GEN_23 ? _slots_4_io_out_uop_bypassable : _GEN_22 ? _slots_3_io_out_uop_bypassable : _slots_2_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_24 ? _slots_5_io_out_uop_mem_cmd : _GEN_23 ? _slots_4_io_out_uop_mem_cmd : _GEN_22 ? _slots_3_io_out_uop_mem_cmd : _slots_2_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_24 ? _slots_5_io_out_uop_mem_size : _GEN_23 ? _slots_4_io_out_uop_mem_size : _GEN_22 ? _slots_3_io_out_uop_mem_size : _slots_2_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_24 ? _slots_5_io_out_uop_mem_signed : _GEN_23 ? _slots_4_io_out_uop_mem_signed : _GEN_22 ? _slots_3_io_out_uop_mem_signed : _slots_2_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_24 ? _slots_5_io_out_uop_is_fence : _GEN_23 ? _slots_4_io_out_uop_is_fence : _GEN_22 ? _slots_3_io_out_uop_is_fence : _slots_2_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_24 ? _slots_5_io_out_uop_is_fencei : _GEN_23 ? _slots_4_io_out_uop_is_fencei : _GEN_22 ? _slots_3_io_out_uop_is_fencei : _slots_2_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_24 ? _slots_5_io_out_uop_is_amo : _GEN_23 ? _slots_4_io_out_uop_is_amo : _GEN_22 ? _slots_3_io_out_uop_is_amo : _slots_2_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_24 ? _slots_5_io_out_uop_uses_ldq : _GEN_23 ? _slots_4_io_out_uop_uses_ldq : _GEN_22 ? _slots_3_io_out_uop_uses_ldq : _slots_2_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_24 ? _slots_5_io_out_uop_uses_stq : _GEN_23 ? _slots_4_io_out_uop_uses_stq : _GEN_22 ? _slots_3_io_out_uop_uses_stq : _slots_2_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_24 ? _slots_5_io_out_uop_is_sys_pc2epc : _GEN_23 ? _slots_4_io_out_uop_is_sys_pc2epc : _GEN_22 ? _slots_3_io_out_uop_is_sys_pc2epc : _slots_2_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_24 ? _slots_5_io_out_uop_is_unique : _GEN_23 ? _slots_4_io_out_uop_is_unique : _GEN_22 ? _slots_3_io_out_uop_is_unique : _slots_2_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_24 ? _slots_5_io_out_uop_flush_on_commit : _GEN_23 ? _slots_4_io_out_uop_flush_on_commit : _GEN_22 ? _slots_3_io_out_uop_flush_on_commit : _slots_2_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_24 ? _slots_5_io_out_uop_ldst_is_rs1 : _GEN_23 ? _slots_4_io_out_uop_ldst_is_rs1 : _GEN_22 ? _slots_3_io_out_uop_ldst_is_rs1 : _slots_2_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_24 ? _slots_5_io_out_uop_ldst : _GEN_23 ? _slots_4_io_out_uop_ldst : _GEN_22 ? _slots_3_io_out_uop_ldst : _slots_2_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_24 ? _slots_5_io_out_uop_lrs1 : _GEN_23 ? _slots_4_io_out_uop_lrs1 : _GEN_22 ? _slots_3_io_out_uop_lrs1 : _slots_2_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_24 ? _slots_5_io_out_uop_lrs2 : _GEN_23 ? _slots_4_io_out_uop_lrs2 : _GEN_22 ? _slots_3_io_out_uop_lrs2 : _slots_2_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_24 ? _slots_5_io_out_uop_lrs3 : _GEN_23 ? _slots_4_io_out_uop_lrs3 : _GEN_22 ? _slots_3_io_out_uop_lrs3 : _slots_2_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_24 ? _slots_5_io_out_uop_ldst_val : _GEN_23 ? _slots_4_io_out_uop_ldst_val : _GEN_22 ? _slots_3_io_out_uop_ldst_val : _slots_2_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_24 ? _slots_5_io_out_uop_dst_rtype : _GEN_23 ? _slots_4_io_out_uop_dst_rtype : _GEN_22 ? _slots_3_io_out_uop_dst_rtype : _slots_2_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_24 ? _slots_5_io_out_uop_lrs1_rtype : _GEN_23 ? _slots_4_io_out_uop_lrs1_rtype : _GEN_22 ? _slots_3_io_out_uop_lrs1_rtype : _slots_2_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_24 ? _slots_5_io_out_uop_lrs2_rtype : _GEN_23 ? _slots_4_io_out_uop_lrs2_rtype : _GEN_22 ? _slots_3_io_out_uop_lrs2_rtype : _slots_2_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_24 ? _slots_5_io_out_uop_frs3_en : _GEN_23 ? _slots_4_io_out_uop_frs3_en : _GEN_22 ? _slots_3_io_out_uop_frs3_en : _slots_2_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_24 ? _slots_5_io_out_uop_fp_val : _GEN_23 ? _slots_4_io_out_uop_fp_val : _GEN_22 ? _slots_3_io_out_uop_fp_val : _slots_2_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_24 ? _slots_5_io_out_uop_fp_single : _GEN_23 ? _slots_4_io_out_uop_fp_single : _GEN_22 ? _slots_3_io_out_uop_fp_single : _slots_2_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_24 ? _slots_5_io_out_uop_xcpt_pf_if : _GEN_23 ? _slots_4_io_out_uop_xcpt_pf_if : _GEN_22 ? _slots_3_io_out_uop_xcpt_pf_if : _slots_2_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_24 ? _slots_5_io_out_uop_xcpt_ae_if : _GEN_23 ? _slots_4_io_out_uop_xcpt_ae_if : _GEN_22 ? _slots_3_io_out_uop_xcpt_ae_if : _slots_2_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_24 ? _slots_5_io_out_uop_xcpt_ma_if : _GEN_23 ? _slots_4_io_out_uop_xcpt_ma_if : _GEN_22 ? _slots_3_io_out_uop_xcpt_ma_if : _slots_2_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_24 ? _slots_5_io_out_uop_bp_debug_if : _GEN_23 ? _slots_4_io_out_uop_bp_debug_if : _GEN_22 ? _slots_3_io_out_uop_bp_debug_if : _slots_2_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_24 ? _slots_5_io_out_uop_bp_xcpt_if : _GEN_23 ? _slots_4_io_out_uop_bp_xcpt_if : _GEN_22 ? _slots_3_io_out_uop_bp_xcpt_if : _slots_2_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_24 ? _slots_5_io_out_uop_debug_fsrc : _GEN_23 ? _slots_4_io_out_uop_debug_fsrc : _GEN_22 ? _slots_3_io_out_uop_debug_fsrc : _slots_2_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_24 ? _slots_5_io_out_uop_debug_tsrc : _GEN_23 ? _slots_4_io_out_uop_debug_tsrc : _GEN_22 ? _slots_3_io_out_uop_debug_tsrc : _slots_2_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_1_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_1_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_1_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_1_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_1_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_1_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_1_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_1_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_1_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_1_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_1_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_1_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_1_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_1_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_1_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_1_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_1_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_1_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_1_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_1_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_1_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_1_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_1_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_1_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_1_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_1_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_1_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_1_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_1_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_1_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_1_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_1_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_1_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_1_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_1_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_1_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_1_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_1_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_1_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_1_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_1_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_1_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_1_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_1_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_1_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_1_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_1_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_1_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_1_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_1_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_1_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_1_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_1_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_1_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_1_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_1_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_1_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_1_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_1_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_1_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_1_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_1_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_1_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_1_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_1_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_1_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_1_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_1_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_1_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_1_io_uop_uopc),
    .io_uop_inst                    (_slots_1_io_uop_inst),
    .io_uop_debug_inst              (_slots_1_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_1_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_1_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_1_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_1_io_uop_fu_code),
    .io_uop_iw_state                (_slots_1_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_1_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_1_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_1_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_1_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_1_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_1_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_1_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_1_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_1_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_1_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_1_io_uop_pc_lob),
    .io_uop_taken                   (_slots_1_io_uop_taken),
    .io_uop_imm_packed              (_slots_1_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_1_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_1_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_1_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_1_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_1_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_1_io_uop_pdst),
    .io_uop_prs1                    (_slots_1_io_uop_prs1),
    .io_uop_prs2                    (_slots_1_io_uop_prs2),
    .io_uop_prs3                    (_slots_1_io_uop_prs3),
    .io_uop_ppred                   (_slots_1_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_1_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_1_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_1_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_1_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_1_io_uop_stale_pdst),
    .io_uop_exception               (_slots_1_io_uop_exception),
    .io_uop_exc_cause               (_slots_1_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_1_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_1_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_1_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_1_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_1_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_1_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_1_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_1_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_1_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_1_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_1_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_1_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_1_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_1_io_uop_ldst),
    .io_uop_lrs1                    (_slots_1_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_1_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_1_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_1_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_1_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_1_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_1_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_1_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_1_io_uop_fp_val),
    .io_uop_fp_single               (_slots_1_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_1_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_1_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_1_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_1_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_1_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_1_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_1_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_2 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_2_io_valid),
    .io_will_be_valid               (_slots_2_io_will_be_valid),
    .io_request                     (_slots_2_io_request),
    .io_grant                       (issue_slots_2_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_next_1_1to0),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_2_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_27 ? _slots_6_io_out_uop_uopc : _GEN_26 ? _slots_5_io_out_uop_uopc : _GEN_25 ? _slots_4_io_out_uop_uopc : _slots_3_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_27 ? _slots_6_io_out_uop_inst : _GEN_26 ? _slots_5_io_out_uop_inst : _GEN_25 ? _slots_4_io_out_uop_inst : _slots_3_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_27 ? _slots_6_io_out_uop_debug_inst : _GEN_26 ? _slots_5_io_out_uop_debug_inst : _GEN_25 ? _slots_4_io_out_uop_debug_inst : _slots_3_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_27 ? _slots_6_io_out_uop_is_rvc : _GEN_26 ? _slots_5_io_out_uop_is_rvc : _GEN_25 ? _slots_4_io_out_uop_is_rvc : _slots_3_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_27 ? _slots_6_io_out_uop_debug_pc : _GEN_26 ? _slots_5_io_out_uop_debug_pc : _GEN_25 ? _slots_4_io_out_uop_debug_pc : _slots_3_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_27 ? _slots_6_io_out_uop_iq_type : _GEN_26 ? _slots_5_io_out_uop_iq_type : _GEN_25 ? _slots_4_io_out_uop_iq_type : _slots_3_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_27 ? _slots_6_io_out_uop_fu_code : _GEN_26 ? _slots_5_io_out_uop_fu_code : _GEN_25 ? _slots_4_io_out_uop_fu_code : _slots_3_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_27 ? _slots_6_io_out_uop_iw_state : _GEN_26 ? _slots_5_io_out_uop_iw_state : _GEN_25 ? _slots_4_io_out_uop_iw_state : _slots_3_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_27 ? _slots_6_io_out_uop_iw_p1_poisoned : _GEN_26 ? _slots_5_io_out_uop_iw_p1_poisoned : _GEN_25 ? _slots_4_io_out_uop_iw_p1_poisoned : _slots_3_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_27 ? _slots_6_io_out_uop_iw_p2_poisoned : _GEN_26 ? _slots_5_io_out_uop_iw_p2_poisoned : _GEN_25 ? _slots_4_io_out_uop_iw_p2_poisoned : _slots_3_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_27 ? _slots_6_io_out_uop_is_br : _GEN_26 ? _slots_5_io_out_uop_is_br : _GEN_25 ? _slots_4_io_out_uop_is_br : _slots_3_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_27 ? _slots_6_io_out_uop_is_jalr : _GEN_26 ? _slots_5_io_out_uop_is_jalr : _GEN_25 ? _slots_4_io_out_uop_is_jalr : _slots_3_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_27 ? _slots_6_io_out_uop_is_jal : _GEN_26 ? _slots_5_io_out_uop_is_jal : _GEN_25 ? _slots_4_io_out_uop_is_jal : _slots_3_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_27 ? _slots_6_io_out_uop_is_sfb : _GEN_26 ? _slots_5_io_out_uop_is_sfb : _GEN_25 ? _slots_4_io_out_uop_is_sfb : _slots_3_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_27 ? _slots_6_io_out_uop_br_mask : _GEN_26 ? _slots_5_io_out_uop_br_mask : _GEN_25 ? _slots_4_io_out_uop_br_mask : _slots_3_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_27 ? _slots_6_io_out_uop_br_tag : _GEN_26 ? _slots_5_io_out_uop_br_tag : _GEN_25 ? _slots_4_io_out_uop_br_tag : _slots_3_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_27 ? _slots_6_io_out_uop_ftq_idx : _GEN_26 ? _slots_5_io_out_uop_ftq_idx : _GEN_25 ? _slots_4_io_out_uop_ftq_idx : _slots_3_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_27 ? _slots_6_io_out_uop_edge_inst : _GEN_26 ? _slots_5_io_out_uop_edge_inst : _GEN_25 ? _slots_4_io_out_uop_edge_inst : _slots_3_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_27 ? _slots_6_io_out_uop_pc_lob : _GEN_26 ? _slots_5_io_out_uop_pc_lob : _GEN_25 ? _slots_4_io_out_uop_pc_lob : _slots_3_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_27 ? _slots_6_io_out_uop_taken : _GEN_26 ? _slots_5_io_out_uop_taken : _GEN_25 ? _slots_4_io_out_uop_taken : _slots_3_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_27 ? _slots_6_io_out_uop_imm_packed : _GEN_26 ? _slots_5_io_out_uop_imm_packed : _GEN_25 ? _slots_4_io_out_uop_imm_packed : _slots_3_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_27 ? _slots_6_io_out_uop_csr_addr : _GEN_26 ? _slots_5_io_out_uop_csr_addr : _GEN_25 ? _slots_4_io_out_uop_csr_addr : _slots_3_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_27 ? _slots_6_io_out_uop_rob_idx : _GEN_26 ? _slots_5_io_out_uop_rob_idx : _GEN_25 ? _slots_4_io_out_uop_rob_idx : _slots_3_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_27 ? _slots_6_io_out_uop_ldq_idx : _GEN_26 ? _slots_5_io_out_uop_ldq_idx : _GEN_25 ? _slots_4_io_out_uop_ldq_idx : _slots_3_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_27 ? _slots_6_io_out_uop_stq_idx : _GEN_26 ? _slots_5_io_out_uop_stq_idx : _GEN_25 ? _slots_4_io_out_uop_stq_idx : _slots_3_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_27 ? _slots_6_io_out_uop_rxq_idx : _GEN_26 ? _slots_5_io_out_uop_rxq_idx : _GEN_25 ? _slots_4_io_out_uop_rxq_idx : _slots_3_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_27 ? _slots_6_io_out_uop_pdst : _GEN_26 ? _slots_5_io_out_uop_pdst : _GEN_25 ? _slots_4_io_out_uop_pdst : _slots_3_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_27 ? _slots_6_io_out_uop_prs1 : _GEN_26 ? _slots_5_io_out_uop_prs1 : _GEN_25 ? _slots_4_io_out_uop_prs1 : _slots_3_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_27 ? _slots_6_io_out_uop_prs2 : _GEN_26 ? _slots_5_io_out_uop_prs2 : _GEN_25 ? _slots_4_io_out_uop_prs2 : _slots_3_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_27 ? _slots_6_io_out_uop_prs3 : _GEN_26 ? _slots_5_io_out_uop_prs3 : _GEN_25 ? _slots_4_io_out_uop_prs3 : _slots_3_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_27 ? _slots_6_io_out_uop_ppred : _GEN_26 ? _slots_5_io_out_uop_ppred : _GEN_25 ? _slots_4_io_out_uop_ppred : _slots_3_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_27 ? _slots_6_io_out_uop_prs1_busy : _GEN_26 ? _slots_5_io_out_uop_prs1_busy : _GEN_25 ? _slots_4_io_out_uop_prs1_busy : _slots_3_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_27 ? _slots_6_io_out_uop_prs2_busy : _GEN_26 ? _slots_5_io_out_uop_prs2_busy : _GEN_25 ? _slots_4_io_out_uop_prs2_busy : _slots_3_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_27 ? _slots_6_io_out_uop_prs3_busy : _GEN_26 ? _slots_5_io_out_uop_prs3_busy : _GEN_25 ? _slots_4_io_out_uop_prs3_busy : _slots_3_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_27 ? _slots_6_io_out_uop_ppred_busy : _GEN_26 ? _slots_5_io_out_uop_ppred_busy : _GEN_25 ? _slots_4_io_out_uop_ppred_busy : _slots_3_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_27 ? _slots_6_io_out_uop_stale_pdst : _GEN_26 ? _slots_5_io_out_uop_stale_pdst : _GEN_25 ? _slots_4_io_out_uop_stale_pdst : _slots_3_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_27 ? _slots_6_io_out_uop_exception : _GEN_26 ? _slots_5_io_out_uop_exception : _GEN_25 ? _slots_4_io_out_uop_exception : _slots_3_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_27 ? _slots_6_io_out_uop_exc_cause : _GEN_26 ? _slots_5_io_out_uop_exc_cause : _GEN_25 ? _slots_4_io_out_uop_exc_cause : _slots_3_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_27 ? _slots_6_io_out_uop_bypassable : _GEN_26 ? _slots_5_io_out_uop_bypassable : _GEN_25 ? _slots_4_io_out_uop_bypassable : _slots_3_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_27 ? _slots_6_io_out_uop_mem_cmd : _GEN_26 ? _slots_5_io_out_uop_mem_cmd : _GEN_25 ? _slots_4_io_out_uop_mem_cmd : _slots_3_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_27 ? _slots_6_io_out_uop_mem_size : _GEN_26 ? _slots_5_io_out_uop_mem_size : _GEN_25 ? _slots_4_io_out_uop_mem_size : _slots_3_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_27 ? _slots_6_io_out_uop_mem_signed : _GEN_26 ? _slots_5_io_out_uop_mem_signed : _GEN_25 ? _slots_4_io_out_uop_mem_signed : _slots_3_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_27 ? _slots_6_io_out_uop_is_fence : _GEN_26 ? _slots_5_io_out_uop_is_fence : _GEN_25 ? _slots_4_io_out_uop_is_fence : _slots_3_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_27 ? _slots_6_io_out_uop_is_fencei : _GEN_26 ? _slots_5_io_out_uop_is_fencei : _GEN_25 ? _slots_4_io_out_uop_is_fencei : _slots_3_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_27 ? _slots_6_io_out_uop_is_amo : _GEN_26 ? _slots_5_io_out_uop_is_amo : _GEN_25 ? _slots_4_io_out_uop_is_amo : _slots_3_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_27 ? _slots_6_io_out_uop_uses_ldq : _GEN_26 ? _slots_5_io_out_uop_uses_ldq : _GEN_25 ? _slots_4_io_out_uop_uses_ldq : _slots_3_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_27 ? _slots_6_io_out_uop_uses_stq : _GEN_26 ? _slots_5_io_out_uop_uses_stq : _GEN_25 ? _slots_4_io_out_uop_uses_stq : _slots_3_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_27 ? _slots_6_io_out_uop_is_sys_pc2epc : _GEN_26 ? _slots_5_io_out_uop_is_sys_pc2epc : _GEN_25 ? _slots_4_io_out_uop_is_sys_pc2epc : _slots_3_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_27 ? _slots_6_io_out_uop_is_unique : _GEN_26 ? _slots_5_io_out_uop_is_unique : _GEN_25 ? _slots_4_io_out_uop_is_unique : _slots_3_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_27 ? _slots_6_io_out_uop_flush_on_commit : _GEN_26 ? _slots_5_io_out_uop_flush_on_commit : _GEN_25 ? _slots_4_io_out_uop_flush_on_commit : _slots_3_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_27 ? _slots_6_io_out_uop_ldst_is_rs1 : _GEN_26 ? _slots_5_io_out_uop_ldst_is_rs1 : _GEN_25 ? _slots_4_io_out_uop_ldst_is_rs1 : _slots_3_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_27 ? _slots_6_io_out_uop_ldst : _GEN_26 ? _slots_5_io_out_uop_ldst : _GEN_25 ? _slots_4_io_out_uop_ldst : _slots_3_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_27 ? _slots_6_io_out_uop_lrs1 : _GEN_26 ? _slots_5_io_out_uop_lrs1 : _GEN_25 ? _slots_4_io_out_uop_lrs1 : _slots_3_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_27 ? _slots_6_io_out_uop_lrs2 : _GEN_26 ? _slots_5_io_out_uop_lrs2 : _GEN_25 ? _slots_4_io_out_uop_lrs2 : _slots_3_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_27 ? _slots_6_io_out_uop_lrs3 : _GEN_26 ? _slots_5_io_out_uop_lrs3 : _GEN_25 ? _slots_4_io_out_uop_lrs3 : _slots_3_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_27 ? _slots_6_io_out_uop_ldst_val : _GEN_26 ? _slots_5_io_out_uop_ldst_val : _GEN_25 ? _slots_4_io_out_uop_ldst_val : _slots_3_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_27 ? _slots_6_io_out_uop_dst_rtype : _GEN_26 ? _slots_5_io_out_uop_dst_rtype : _GEN_25 ? _slots_4_io_out_uop_dst_rtype : _slots_3_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_27 ? _slots_6_io_out_uop_lrs1_rtype : _GEN_26 ? _slots_5_io_out_uop_lrs1_rtype : _GEN_25 ? _slots_4_io_out_uop_lrs1_rtype : _slots_3_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_27 ? _slots_6_io_out_uop_lrs2_rtype : _GEN_26 ? _slots_5_io_out_uop_lrs2_rtype : _GEN_25 ? _slots_4_io_out_uop_lrs2_rtype : _slots_3_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_27 ? _slots_6_io_out_uop_frs3_en : _GEN_26 ? _slots_5_io_out_uop_frs3_en : _GEN_25 ? _slots_4_io_out_uop_frs3_en : _slots_3_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_27 ? _slots_6_io_out_uop_fp_val : _GEN_26 ? _slots_5_io_out_uop_fp_val : _GEN_25 ? _slots_4_io_out_uop_fp_val : _slots_3_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_27 ? _slots_6_io_out_uop_fp_single : _GEN_26 ? _slots_5_io_out_uop_fp_single : _GEN_25 ? _slots_4_io_out_uop_fp_single : _slots_3_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_27 ? _slots_6_io_out_uop_xcpt_pf_if : _GEN_26 ? _slots_5_io_out_uop_xcpt_pf_if : _GEN_25 ? _slots_4_io_out_uop_xcpt_pf_if : _slots_3_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_27 ? _slots_6_io_out_uop_xcpt_ae_if : _GEN_26 ? _slots_5_io_out_uop_xcpt_ae_if : _GEN_25 ? _slots_4_io_out_uop_xcpt_ae_if : _slots_3_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_27 ? _slots_6_io_out_uop_xcpt_ma_if : _GEN_26 ? _slots_5_io_out_uop_xcpt_ma_if : _GEN_25 ? _slots_4_io_out_uop_xcpt_ma_if : _slots_3_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_27 ? _slots_6_io_out_uop_bp_debug_if : _GEN_26 ? _slots_5_io_out_uop_bp_debug_if : _GEN_25 ? _slots_4_io_out_uop_bp_debug_if : _slots_3_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_27 ? _slots_6_io_out_uop_bp_xcpt_if : _GEN_26 ? _slots_5_io_out_uop_bp_xcpt_if : _GEN_25 ? _slots_4_io_out_uop_bp_xcpt_if : _slots_3_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_27 ? _slots_6_io_out_uop_debug_fsrc : _GEN_26 ? _slots_5_io_out_uop_debug_fsrc : _GEN_25 ? _slots_4_io_out_uop_debug_fsrc : _slots_3_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_27 ? _slots_6_io_out_uop_debug_tsrc : _GEN_26 ? _slots_5_io_out_uop_debug_tsrc : _GEN_25 ? _slots_4_io_out_uop_debug_tsrc : _slots_3_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_2_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_2_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_2_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_2_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_2_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_2_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_2_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_2_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_2_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_2_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_2_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_2_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_2_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_2_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_2_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_2_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_2_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_2_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_2_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_2_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_2_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_2_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_2_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_2_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_2_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_2_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_2_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_2_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_2_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_2_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_2_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_2_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_2_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_2_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_2_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_2_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_2_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_2_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_2_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_2_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_2_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_2_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_2_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_2_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_2_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_2_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_2_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_2_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_2_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_2_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_2_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_2_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_2_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_2_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_2_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_2_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_2_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_2_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_2_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_2_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_2_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_2_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_2_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_2_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_2_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_2_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_2_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_2_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_2_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_2_io_uop_uopc),
    .io_uop_inst                    (_slots_2_io_uop_inst),
    .io_uop_debug_inst              (_slots_2_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_2_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_2_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_2_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_2_io_uop_fu_code),
    .io_uop_iw_state                (_slots_2_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_2_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_2_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_2_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_2_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_2_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_2_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_2_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_2_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_2_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_2_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_2_io_uop_pc_lob),
    .io_uop_taken                   (_slots_2_io_uop_taken),
    .io_uop_imm_packed              (_slots_2_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_2_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_2_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_2_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_2_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_2_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_2_io_uop_pdst),
    .io_uop_prs1                    (_slots_2_io_uop_prs1),
    .io_uop_prs2                    (_slots_2_io_uop_prs2),
    .io_uop_prs3                    (_slots_2_io_uop_prs3),
    .io_uop_ppred                   (_slots_2_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_2_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_2_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_2_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_2_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_2_io_uop_stale_pdst),
    .io_uop_exception               (_slots_2_io_uop_exception),
    .io_uop_exc_cause               (_slots_2_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_2_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_2_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_2_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_2_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_2_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_2_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_2_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_2_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_2_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_2_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_2_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_2_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_2_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_2_io_uop_ldst),
    .io_uop_lrs1                    (_slots_2_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_2_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_2_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_2_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_2_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_2_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_2_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_2_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_2_io_uop_fp_val),
    .io_uop_fp_single               (_slots_2_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_2_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_2_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_2_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_2_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_2_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_2_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_2_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_3 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_3_io_valid),
    .io_will_be_valid               (_slots_3_io_will_be_valid),
    .io_request                     (_slots_3_io_request),
    .io_grant                       (issue_slots_3_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_2),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_3_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_30 ? _slots_7_io_out_uop_uopc : _GEN_29 ? _slots_6_io_out_uop_uopc : _GEN_28 ? _slots_5_io_out_uop_uopc : _slots_4_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_30 ? _slots_7_io_out_uop_inst : _GEN_29 ? _slots_6_io_out_uop_inst : _GEN_28 ? _slots_5_io_out_uop_inst : _slots_4_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_30 ? _slots_7_io_out_uop_debug_inst : _GEN_29 ? _slots_6_io_out_uop_debug_inst : _GEN_28 ? _slots_5_io_out_uop_debug_inst : _slots_4_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_30 ? _slots_7_io_out_uop_is_rvc : _GEN_29 ? _slots_6_io_out_uop_is_rvc : _GEN_28 ? _slots_5_io_out_uop_is_rvc : _slots_4_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_30 ? _slots_7_io_out_uop_debug_pc : _GEN_29 ? _slots_6_io_out_uop_debug_pc : _GEN_28 ? _slots_5_io_out_uop_debug_pc : _slots_4_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_30 ? _slots_7_io_out_uop_iq_type : _GEN_29 ? _slots_6_io_out_uop_iq_type : _GEN_28 ? _slots_5_io_out_uop_iq_type : _slots_4_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_30 ? _slots_7_io_out_uop_fu_code : _GEN_29 ? _slots_6_io_out_uop_fu_code : _GEN_28 ? _slots_5_io_out_uop_fu_code : _slots_4_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_30 ? _slots_7_io_out_uop_iw_state : _GEN_29 ? _slots_6_io_out_uop_iw_state : _GEN_28 ? _slots_5_io_out_uop_iw_state : _slots_4_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_30 ? _slots_7_io_out_uop_iw_p1_poisoned : _GEN_29 ? _slots_6_io_out_uop_iw_p1_poisoned : _GEN_28 ? _slots_5_io_out_uop_iw_p1_poisoned : _slots_4_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_30 ? _slots_7_io_out_uop_iw_p2_poisoned : _GEN_29 ? _slots_6_io_out_uop_iw_p2_poisoned : _GEN_28 ? _slots_5_io_out_uop_iw_p2_poisoned : _slots_4_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_30 ? _slots_7_io_out_uop_is_br : _GEN_29 ? _slots_6_io_out_uop_is_br : _GEN_28 ? _slots_5_io_out_uop_is_br : _slots_4_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_30 ? _slots_7_io_out_uop_is_jalr : _GEN_29 ? _slots_6_io_out_uop_is_jalr : _GEN_28 ? _slots_5_io_out_uop_is_jalr : _slots_4_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_30 ? _slots_7_io_out_uop_is_jal : _GEN_29 ? _slots_6_io_out_uop_is_jal : _GEN_28 ? _slots_5_io_out_uop_is_jal : _slots_4_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_30 ? _slots_7_io_out_uop_is_sfb : _GEN_29 ? _slots_6_io_out_uop_is_sfb : _GEN_28 ? _slots_5_io_out_uop_is_sfb : _slots_4_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_30 ? _slots_7_io_out_uop_br_mask : _GEN_29 ? _slots_6_io_out_uop_br_mask : _GEN_28 ? _slots_5_io_out_uop_br_mask : _slots_4_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_30 ? _slots_7_io_out_uop_br_tag : _GEN_29 ? _slots_6_io_out_uop_br_tag : _GEN_28 ? _slots_5_io_out_uop_br_tag : _slots_4_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_30 ? _slots_7_io_out_uop_ftq_idx : _GEN_29 ? _slots_6_io_out_uop_ftq_idx : _GEN_28 ? _slots_5_io_out_uop_ftq_idx : _slots_4_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_30 ? _slots_7_io_out_uop_edge_inst : _GEN_29 ? _slots_6_io_out_uop_edge_inst : _GEN_28 ? _slots_5_io_out_uop_edge_inst : _slots_4_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_30 ? _slots_7_io_out_uop_pc_lob : _GEN_29 ? _slots_6_io_out_uop_pc_lob : _GEN_28 ? _slots_5_io_out_uop_pc_lob : _slots_4_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_30 ? _slots_7_io_out_uop_taken : _GEN_29 ? _slots_6_io_out_uop_taken : _GEN_28 ? _slots_5_io_out_uop_taken : _slots_4_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_30 ? _slots_7_io_out_uop_imm_packed : _GEN_29 ? _slots_6_io_out_uop_imm_packed : _GEN_28 ? _slots_5_io_out_uop_imm_packed : _slots_4_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_30 ? _slots_7_io_out_uop_csr_addr : _GEN_29 ? _slots_6_io_out_uop_csr_addr : _GEN_28 ? _slots_5_io_out_uop_csr_addr : _slots_4_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_30 ? _slots_7_io_out_uop_rob_idx : _GEN_29 ? _slots_6_io_out_uop_rob_idx : _GEN_28 ? _slots_5_io_out_uop_rob_idx : _slots_4_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_30 ? _slots_7_io_out_uop_ldq_idx : _GEN_29 ? _slots_6_io_out_uop_ldq_idx : _GEN_28 ? _slots_5_io_out_uop_ldq_idx : _slots_4_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_30 ? _slots_7_io_out_uop_stq_idx : _GEN_29 ? _slots_6_io_out_uop_stq_idx : _GEN_28 ? _slots_5_io_out_uop_stq_idx : _slots_4_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_30 ? _slots_7_io_out_uop_rxq_idx : _GEN_29 ? _slots_6_io_out_uop_rxq_idx : _GEN_28 ? _slots_5_io_out_uop_rxq_idx : _slots_4_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_30 ? _slots_7_io_out_uop_pdst : _GEN_29 ? _slots_6_io_out_uop_pdst : _GEN_28 ? _slots_5_io_out_uop_pdst : _slots_4_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_30 ? _slots_7_io_out_uop_prs1 : _GEN_29 ? _slots_6_io_out_uop_prs1 : _GEN_28 ? _slots_5_io_out_uop_prs1 : _slots_4_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_30 ? _slots_7_io_out_uop_prs2 : _GEN_29 ? _slots_6_io_out_uop_prs2 : _GEN_28 ? _slots_5_io_out_uop_prs2 : _slots_4_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_30 ? _slots_7_io_out_uop_prs3 : _GEN_29 ? _slots_6_io_out_uop_prs3 : _GEN_28 ? _slots_5_io_out_uop_prs3 : _slots_4_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_30 ? _slots_7_io_out_uop_ppred : _GEN_29 ? _slots_6_io_out_uop_ppred : _GEN_28 ? _slots_5_io_out_uop_ppred : _slots_4_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_30 ? _slots_7_io_out_uop_prs1_busy : _GEN_29 ? _slots_6_io_out_uop_prs1_busy : _GEN_28 ? _slots_5_io_out_uop_prs1_busy : _slots_4_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_30 ? _slots_7_io_out_uop_prs2_busy : _GEN_29 ? _slots_6_io_out_uop_prs2_busy : _GEN_28 ? _slots_5_io_out_uop_prs2_busy : _slots_4_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_30 ? _slots_7_io_out_uop_prs3_busy : _GEN_29 ? _slots_6_io_out_uop_prs3_busy : _GEN_28 ? _slots_5_io_out_uop_prs3_busy : _slots_4_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_30 ? _slots_7_io_out_uop_ppred_busy : _GEN_29 ? _slots_6_io_out_uop_ppred_busy : _GEN_28 ? _slots_5_io_out_uop_ppred_busy : _slots_4_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_30 ? _slots_7_io_out_uop_stale_pdst : _GEN_29 ? _slots_6_io_out_uop_stale_pdst : _GEN_28 ? _slots_5_io_out_uop_stale_pdst : _slots_4_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_30 ? _slots_7_io_out_uop_exception : _GEN_29 ? _slots_6_io_out_uop_exception : _GEN_28 ? _slots_5_io_out_uop_exception : _slots_4_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_30 ? _slots_7_io_out_uop_exc_cause : _GEN_29 ? _slots_6_io_out_uop_exc_cause : _GEN_28 ? _slots_5_io_out_uop_exc_cause : _slots_4_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_30 ? _slots_7_io_out_uop_bypassable : _GEN_29 ? _slots_6_io_out_uop_bypassable : _GEN_28 ? _slots_5_io_out_uop_bypassable : _slots_4_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_30 ? _slots_7_io_out_uop_mem_cmd : _GEN_29 ? _slots_6_io_out_uop_mem_cmd : _GEN_28 ? _slots_5_io_out_uop_mem_cmd : _slots_4_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_30 ? _slots_7_io_out_uop_mem_size : _GEN_29 ? _slots_6_io_out_uop_mem_size : _GEN_28 ? _slots_5_io_out_uop_mem_size : _slots_4_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_30 ? _slots_7_io_out_uop_mem_signed : _GEN_29 ? _slots_6_io_out_uop_mem_signed : _GEN_28 ? _slots_5_io_out_uop_mem_signed : _slots_4_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_30 ? _slots_7_io_out_uop_is_fence : _GEN_29 ? _slots_6_io_out_uop_is_fence : _GEN_28 ? _slots_5_io_out_uop_is_fence : _slots_4_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_30 ? _slots_7_io_out_uop_is_fencei : _GEN_29 ? _slots_6_io_out_uop_is_fencei : _GEN_28 ? _slots_5_io_out_uop_is_fencei : _slots_4_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_30 ? _slots_7_io_out_uop_is_amo : _GEN_29 ? _slots_6_io_out_uop_is_amo : _GEN_28 ? _slots_5_io_out_uop_is_amo : _slots_4_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_30 ? _slots_7_io_out_uop_uses_ldq : _GEN_29 ? _slots_6_io_out_uop_uses_ldq : _GEN_28 ? _slots_5_io_out_uop_uses_ldq : _slots_4_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_30 ? _slots_7_io_out_uop_uses_stq : _GEN_29 ? _slots_6_io_out_uop_uses_stq : _GEN_28 ? _slots_5_io_out_uop_uses_stq : _slots_4_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_30 ? _slots_7_io_out_uop_is_sys_pc2epc : _GEN_29 ? _slots_6_io_out_uop_is_sys_pc2epc : _GEN_28 ? _slots_5_io_out_uop_is_sys_pc2epc : _slots_4_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_30 ? _slots_7_io_out_uop_is_unique : _GEN_29 ? _slots_6_io_out_uop_is_unique : _GEN_28 ? _slots_5_io_out_uop_is_unique : _slots_4_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_30 ? _slots_7_io_out_uop_flush_on_commit : _GEN_29 ? _slots_6_io_out_uop_flush_on_commit : _GEN_28 ? _slots_5_io_out_uop_flush_on_commit : _slots_4_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_30 ? _slots_7_io_out_uop_ldst_is_rs1 : _GEN_29 ? _slots_6_io_out_uop_ldst_is_rs1 : _GEN_28 ? _slots_5_io_out_uop_ldst_is_rs1 : _slots_4_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_30 ? _slots_7_io_out_uop_ldst : _GEN_29 ? _slots_6_io_out_uop_ldst : _GEN_28 ? _slots_5_io_out_uop_ldst : _slots_4_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_30 ? _slots_7_io_out_uop_lrs1 : _GEN_29 ? _slots_6_io_out_uop_lrs1 : _GEN_28 ? _slots_5_io_out_uop_lrs1 : _slots_4_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_30 ? _slots_7_io_out_uop_lrs2 : _GEN_29 ? _slots_6_io_out_uop_lrs2 : _GEN_28 ? _slots_5_io_out_uop_lrs2 : _slots_4_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_30 ? _slots_7_io_out_uop_lrs3 : _GEN_29 ? _slots_6_io_out_uop_lrs3 : _GEN_28 ? _slots_5_io_out_uop_lrs3 : _slots_4_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_30 ? _slots_7_io_out_uop_ldst_val : _GEN_29 ? _slots_6_io_out_uop_ldst_val : _GEN_28 ? _slots_5_io_out_uop_ldst_val : _slots_4_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_30 ? _slots_7_io_out_uop_dst_rtype : _GEN_29 ? _slots_6_io_out_uop_dst_rtype : _GEN_28 ? _slots_5_io_out_uop_dst_rtype : _slots_4_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_30 ? _slots_7_io_out_uop_lrs1_rtype : _GEN_29 ? _slots_6_io_out_uop_lrs1_rtype : _GEN_28 ? _slots_5_io_out_uop_lrs1_rtype : _slots_4_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_30 ? _slots_7_io_out_uop_lrs2_rtype : _GEN_29 ? _slots_6_io_out_uop_lrs2_rtype : _GEN_28 ? _slots_5_io_out_uop_lrs2_rtype : _slots_4_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_30 ? _slots_7_io_out_uop_frs3_en : _GEN_29 ? _slots_6_io_out_uop_frs3_en : _GEN_28 ? _slots_5_io_out_uop_frs3_en : _slots_4_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_30 ? _slots_7_io_out_uop_fp_val : _GEN_29 ? _slots_6_io_out_uop_fp_val : _GEN_28 ? _slots_5_io_out_uop_fp_val : _slots_4_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_30 ? _slots_7_io_out_uop_fp_single : _GEN_29 ? _slots_6_io_out_uop_fp_single : _GEN_28 ? _slots_5_io_out_uop_fp_single : _slots_4_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_30 ? _slots_7_io_out_uop_xcpt_pf_if : _GEN_29 ? _slots_6_io_out_uop_xcpt_pf_if : _GEN_28 ? _slots_5_io_out_uop_xcpt_pf_if : _slots_4_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_30 ? _slots_7_io_out_uop_xcpt_ae_if : _GEN_29 ? _slots_6_io_out_uop_xcpt_ae_if : _GEN_28 ? _slots_5_io_out_uop_xcpt_ae_if : _slots_4_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_30 ? _slots_7_io_out_uop_xcpt_ma_if : _GEN_29 ? _slots_6_io_out_uop_xcpt_ma_if : _GEN_28 ? _slots_5_io_out_uop_xcpt_ma_if : _slots_4_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_30 ? _slots_7_io_out_uop_bp_debug_if : _GEN_29 ? _slots_6_io_out_uop_bp_debug_if : _GEN_28 ? _slots_5_io_out_uop_bp_debug_if : _slots_4_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_30 ? _slots_7_io_out_uop_bp_xcpt_if : _GEN_29 ? _slots_6_io_out_uop_bp_xcpt_if : _GEN_28 ? _slots_5_io_out_uop_bp_xcpt_if : _slots_4_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_30 ? _slots_7_io_out_uop_debug_fsrc : _GEN_29 ? _slots_6_io_out_uop_debug_fsrc : _GEN_28 ? _slots_5_io_out_uop_debug_fsrc : _slots_4_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_30 ? _slots_7_io_out_uop_debug_tsrc : _GEN_29 ? _slots_6_io_out_uop_debug_tsrc : _GEN_28 ? _slots_5_io_out_uop_debug_tsrc : _slots_4_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_3_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_3_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_3_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_3_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_3_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_3_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_3_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_3_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_3_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_3_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_3_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_3_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_3_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_3_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_3_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_3_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_3_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_3_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_3_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_3_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_3_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_3_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_3_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_3_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_3_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_3_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_3_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_3_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_3_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_3_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_3_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_3_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_3_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_3_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_3_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_3_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_3_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_3_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_3_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_3_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_3_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_3_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_3_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_3_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_3_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_3_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_3_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_3_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_3_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_3_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_3_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_3_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_3_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_3_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_3_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_3_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_3_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_3_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_3_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_3_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_3_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_3_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_3_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_3_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_3_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_3_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_3_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_3_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_3_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_3_io_uop_uopc),
    .io_uop_inst                    (_slots_3_io_uop_inst),
    .io_uop_debug_inst              (_slots_3_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_3_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_3_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_3_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_3_io_uop_fu_code),
    .io_uop_iw_state                (_slots_3_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_3_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_3_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_3_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_3_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_3_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_3_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_3_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_3_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_3_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_3_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_3_io_uop_pc_lob),
    .io_uop_taken                   (_slots_3_io_uop_taken),
    .io_uop_imm_packed              (_slots_3_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_3_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_3_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_3_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_3_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_3_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_3_io_uop_pdst),
    .io_uop_prs1                    (_slots_3_io_uop_prs1),
    .io_uop_prs2                    (_slots_3_io_uop_prs2),
    .io_uop_prs3                    (_slots_3_io_uop_prs3),
    .io_uop_ppred                   (_slots_3_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_3_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_3_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_3_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_3_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_3_io_uop_stale_pdst),
    .io_uop_exception               (_slots_3_io_uop_exception),
    .io_uop_exc_cause               (_slots_3_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_3_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_3_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_3_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_3_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_3_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_3_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_3_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_3_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_3_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_3_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_3_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_3_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_3_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_3_io_uop_ldst),
    .io_uop_lrs1                    (_slots_3_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_3_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_3_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_3_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_3_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_3_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_3_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_3_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_3_io_uop_fp_val),
    .io_uop_fp_single               (_slots_3_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_3_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_3_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_3_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_3_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_3_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_3_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_3_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_4 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_4_io_valid),
    .io_will_be_valid               (_slots_4_io_will_be_valid),
    .io_request                     (_slots_4_io_request),
    .io_grant                       (issue_slots_4_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_3),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_4_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_33 ? _slots_8_io_out_uop_uopc : _GEN_32 ? _slots_7_io_out_uop_uopc : _GEN_31 ? _slots_6_io_out_uop_uopc : _slots_5_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_33 ? _slots_8_io_out_uop_inst : _GEN_32 ? _slots_7_io_out_uop_inst : _GEN_31 ? _slots_6_io_out_uop_inst : _slots_5_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_33 ? _slots_8_io_out_uop_debug_inst : _GEN_32 ? _slots_7_io_out_uop_debug_inst : _GEN_31 ? _slots_6_io_out_uop_debug_inst : _slots_5_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_33 ? _slots_8_io_out_uop_is_rvc : _GEN_32 ? _slots_7_io_out_uop_is_rvc : _GEN_31 ? _slots_6_io_out_uop_is_rvc : _slots_5_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_33 ? _slots_8_io_out_uop_debug_pc : _GEN_32 ? _slots_7_io_out_uop_debug_pc : _GEN_31 ? _slots_6_io_out_uop_debug_pc : _slots_5_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_33 ? _slots_8_io_out_uop_iq_type : _GEN_32 ? _slots_7_io_out_uop_iq_type : _GEN_31 ? _slots_6_io_out_uop_iq_type : _slots_5_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_33 ? _slots_8_io_out_uop_fu_code : _GEN_32 ? _slots_7_io_out_uop_fu_code : _GEN_31 ? _slots_6_io_out_uop_fu_code : _slots_5_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_33 ? _slots_8_io_out_uop_iw_state : _GEN_32 ? _slots_7_io_out_uop_iw_state : _GEN_31 ? _slots_6_io_out_uop_iw_state : _slots_5_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_33 ? _slots_8_io_out_uop_iw_p1_poisoned : _GEN_32 ? _slots_7_io_out_uop_iw_p1_poisoned : _GEN_31 ? _slots_6_io_out_uop_iw_p1_poisoned : _slots_5_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_33 ? _slots_8_io_out_uop_iw_p2_poisoned : _GEN_32 ? _slots_7_io_out_uop_iw_p2_poisoned : _GEN_31 ? _slots_6_io_out_uop_iw_p2_poisoned : _slots_5_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_33 ? _slots_8_io_out_uop_is_br : _GEN_32 ? _slots_7_io_out_uop_is_br : _GEN_31 ? _slots_6_io_out_uop_is_br : _slots_5_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_33 ? _slots_8_io_out_uop_is_jalr : _GEN_32 ? _slots_7_io_out_uop_is_jalr : _GEN_31 ? _slots_6_io_out_uop_is_jalr : _slots_5_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_33 ? _slots_8_io_out_uop_is_jal : _GEN_32 ? _slots_7_io_out_uop_is_jal : _GEN_31 ? _slots_6_io_out_uop_is_jal : _slots_5_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_33 ? _slots_8_io_out_uop_is_sfb : _GEN_32 ? _slots_7_io_out_uop_is_sfb : _GEN_31 ? _slots_6_io_out_uop_is_sfb : _slots_5_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_33 ? _slots_8_io_out_uop_br_mask : _GEN_32 ? _slots_7_io_out_uop_br_mask : _GEN_31 ? _slots_6_io_out_uop_br_mask : _slots_5_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_33 ? _slots_8_io_out_uop_br_tag : _GEN_32 ? _slots_7_io_out_uop_br_tag : _GEN_31 ? _slots_6_io_out_uop_br_tag : _slots_5_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_33 ? _slots_8_io_out_uop_ftq_idx : _GEN_32 ? _slots_7_io_out_uop_ftq_idx : _GEN_31 ? _slots_6_io_out_uop_ftq_idx : _slots_5_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_33 ? _slots_8_io_out_uop_edge_inst : _GEN_32 ? _slots_7_io_out_uop_edge_inst : _GEN_31 ? _slots_6_io_out_uop_edge_inst : _slots_5_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_33 ? _slots_8_io_out_uop_pc_lob : _GEN_32 ? _slots_7_io_out_uop_pc_lob : _GEN_31 ? _slots_6_io_out_uop_pc_lob : _slots_5_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_33 ? _slots_8_io_out_uop_taken : _GEN_32 ? _slots_7_io_out_uop_taken : _GEN_31 ? _slots_6_io_out_uop_taken : _slots_5_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_33 ? _slots_8_io_out_uop_imm_packed : _GEN_32 ? _slots_7_io_out_uop_imm_packed : _GEN_31 ? _slots_6_io_out_uop_imm_packed : _slots_5_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_33 ? _slots_8_io_out_uop_csr_addr : _GEN_32 ? _slots_7_io_out_uop_csr_addr : _GEN_31 ? _slots_6_io_out_uop_csr_addr : _slots_5_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_33 ? _slots_8_io_out_uop_rob_idx : _GEN_32 ? _slots_7_io_out_uop_rob_idx : _GEN_31 ? _slots_6_io_out_uop_rob_idx : _slots_5_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_33 ? _slots_8_io_out_uop_ldq_idx : _GEN_32 ? _slots_7_io_out_uop_ldq_idx : _GEN_31 ? _slots_6_io_out_uop_ldq_idx : _slots_5_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_33 ? _slots_8_io_out_uop_stq_idx : _GEN_32 ? _slots_7_io_out_uop_stq_idx : _GEN_31 ? _slots_6_io_out_uop_stq_idx : _slots_5_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_33 ? _slots_8_io_out_uop_rxq_idx : _GEN_32 ? _slots_7_io_out_uop_rxq_idx : _GEN_31 ? _slots_6_io_out_uop_rxq_idx : _slots_5_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_33 ? _slots_8_io_out_uop_pdst : _GEN_32 ? _slots_7_io_out_uop_pdst : _GEN_31 ? _slots_6_io_out_uop_pdst : _slots_5_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_33 ? _slots_8_io_out_uop_prs1 : _GEN_32 ? _slots_7_io_out_uop_prs1 : _GEN_31 ? _slots_6_io_out_uop_prs1 : _slots_5_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_33 ? _slots_8_io_out_uop_prs2 : _GEN_32 ? _slots_7_io_out_uop_prs2 : _GEN_31 ? _slots_6_io_out_uop_prs2 : _slots_5_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_33 ? _slots_8_io_out_uop_prs3 : _GEN_32 ? _slots_7_io_out_uop_prs3 : _GEN_31 ? _slots_6_io_out_uop_prs3 : _slots_5_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_33 ? _slots_8_io_out_uop_ppred : _GEN_32 ? _slots_7_io_out_uop_ppred : _GEN_31 ? _slots_6_io_out_uop_ppred : _slots_5_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_33 ? _slots_8_io_out_uop_prs1_busy : _GEN_32 ? _slots_7_io_out_uop_prs1_busy : _GEN_31 ? _slots_6_io_out_uop_prs1_busy : _slots_5_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_33 ? _slots_8_io_out_uop_prs2_busy : _GEN_32 ? _slots_7_io_out_uop_prs2_busy : _GEN_31 ? _slots_6_io_out_uop_prs2_busy : _slots_5_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_33 ? _slots_8_io_out_uop_prs3_busy : _GEN_32 ? _slots_7_io_out_uop_prs3_busy : _GEN_31 ? _slots_6_io_out_uop_prs3_busy : _slots_5_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_33 ? _slots_8_io_out_uop_ppred_busy : _GEN_32 ? _slots_7_io_out_uop_ppred_busy : _GEN_31 ? _slots_6_io_out_uop_ppred_busy : _slots_5_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_33 ? _slots_8_io_out_uop_stale_pdst : _GEN_32 ? _slots_7_io_out_uop_stale_pdst : _GEN_31 ? _slots_6_io_out_uop_stale_pdst : _slots_5_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_33 ? _slots_8_io_out_uop_exception : _GEN_32 ? _slots_7_io_out_uop_exception : _GEN_31 ? _slots_6_io_out_uop_exception : _slots_5_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_33 ? _slots_8_io_out_uop_exc_cause : _GEN_32 ? _slots_7_io_out_uop_exc_cause : _GEN_31 ? _slots_6_io_out_uop_exc_cause : _slots_5_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_33 ? _slots_8_io_out_uop_bypassable : _GEN_32 ? _slots_7_io_out_uop_bypassable : _GEN_31 ? _slots_6_io_out_uop_bypassable : _slots_5_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_33 ? _slots_8_io_out_uop_mem_cmd : _GEN_32 ? _slots_7_io_out_uop_mem_cmd : _GEN_31 ? _slots_6_io_out_uop_mem_cmd : _slots_5_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_33 ? _slots_8_io_out_uop_mem_size : _GEN_32 ? _slots_7_io_out_uop_mem_size : _GEN_31 ? _slots_6_io_out_uop_mem_size : _slots_5_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_33 ? _slots_8_io_out_uop_mem_signed : _GEN_32 ? _slots_7_io_out_uop_mem_signed : _GEN_31 ? _slots_6_io_out_uop_mem_signed : _slots_5_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_33 ? _slots_8_io_out_uop_is_fence : _GEN_32 ? _slots_7_io_out_uop_is_fence : _GEN_31 ? _slots_6_io_out_uop_is_fence : _slots_5_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_33 ? _slots_8_io_out_uop_is_fencei : _GEN_32 ? _slots_7_io_out_uop_is_fencei : _GEN_31 ? _slots_6_io_out_uop_is_fencei : _slots_5_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_33 ? _slots_8_io_out_uop_is_amo : _GEN_32 ? _slots_7_io_out_uop_is_amo : _GEN_31 ? _slots_6_io_out_uop_is_amo : _slots_5_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_33 ? _slots_8_io_out_uop_uses_ldq : _GEN_32 ? _slots_7_io_out_uop_uses_ldq : _GEN_31 ? _slots_6_io_out_uop_uses_ldq : _slots_5_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_33 ? _slots_8_io_out_uop_uses_stq : _GEN_32 ? _slots_7_io_out_uop_uses_stq : _GEN_31 ? _slots_6_io_out_uop_uses_stq : _slots_5_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_33 ? _slots_8_io_out_uop_is_sys_pc2epc : _GEN_32 ? _slots_7_io_out_uop_is_sys_pc2epc : _GEN_31 ? _slots_6_io_out_uop_is_sys_pc2epc : _slots_5_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_33 ? _slots_8_io_out_uop_is_unique : _GEN_32 ? _slots_7_io_out_uop_is_unique : _GEN_31 ? _slots_6_io_out_uop_is_unique : _slots_5_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_33 ? _slots_8_io_out_uop_flush_on_commit : _GEN_32 ? _slots_7_io_out_uop_flush_on_commit : _GEN_31 ? _slots_6_io_out_uop_flush_on_commit : _slots_5_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_33 ? _slots_8_io_out_uop_ldst_is_rs1 : _GEN_32 ? _slots_7_io_out_uop_ldst_is_rs1 : _GEN_31 ? _slots_6_io_out_uop_ldst_is_rs1 : _slots_5_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_33 ? _slots_8_io_out_uop_ldst : _GEN_32 ? _slots_7_io_out_uop_ldst : _GEN_31 ? _slots_6_io_out_uop_ldst : _slots_5_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_33 ? _slots_8_io_out_uop_lrs1 : _GEN_32 ? _slots_7_io_out_uop_lrs1 : _GEN_31 ? _slots_6_io_out_uop_lrs1 : _slots_5_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_33 ? _slots_8_io_out_uop_lrs2 : _GEN_32 ? _slots_7_io_out_uop_lrs2 : _GEN_31 ? _slots_6_io_out_uop_lrs2 : _slots_5_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_33 ? _slots_8_io_out_uop_lrs3 : _GEN_32 ? _slots_7_io_out_uop_lrs3 : _GEN_31 ? _slots_6_io_out_uop_lrs3 : _slots_5_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_33 ? _slots_8_io_out_uop_ldst_val : _GEN_32 ? _slots_7_io_out_uop_ldst_val : _GEN_31 ? _slots_6_io_out_uop_ldst_val : _slots_5_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_33 ? _slots_8_io_out_uop_dst_rtype : _GEN_32 ? _slots_7_io_out_uop_dst_rtype : _GEN_31 ? _slots_6_io_out_uop_dst_rtype : _slots_5_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_33 ? _slots_8_io_out_uop_lrs1_rtype : _GEN_32 ? _slots_7_io_out_uop_lrs1_rtype : _GEN_31 ? _slots_6_io_out_uop_lrs1_rtype : _slots_5_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_33 ? _slots_8_io_out_uop_lrs2_rtype : _GEN_32 ? _slots_7_io_out_uop_lrs2_rtype : _GEN_31 ? _slots_6_io_out_uop_lrs2_rtype : _slots_5_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_33 ? _slots_8_io_out_uop_frs3_en : _GEN_32 ? _slots_7_io_out_uop_frs3_en : _GEN_31 ? _slots_6_io_out_uop_frs3_en : _slots_5_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_33 ? _slots_8_io_out_uop_fp_val : _GEN_32 ? _slots_7_io_out_uop_fp_val : _GEN_31 ? _slots_6_io_out_uop_fp_val : _slots_5_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_33 ? _slots_8_io_out_uop_fp_single : _GEN_32 ? _slots_7_io_out_uop_fp_single : _GEN_31 ? _slots_6_io_out_uop_fp_single : _slots_5_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_33 ? _slots_8_io_out_uop_xcpt_pf_if : _GEN_32 ? _slots_7_io_out_uop_xcpt_pf_if : _GEN_31 ? _slots_6_io_out_uop_xcpt_pf_if : _slots_5_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_33 ? _slots_8_io_out_uop_xcpt_ae_if : _GEN_32 ? _slots_7_io_out_uop_xcpt_ae_if : _GEN_31 ? _slots_6_io_out_uop_xcpt_ae_if : _slots_5_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_33 ? _slots_8_io_out_uop_xcpt_ma_if : _GEN_32 ? _slots_7_io_out_uop_xcpt_ma_if : _GEN_31 ? _slots_6_io_out_uop_xcpt_ma_if : _slots_5_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_33 ? _slots_8_io_out_uop_bp_debug_if : _GEN_32 ? _slots_7_io_out_uop_bp_debug_if : _GEN_31 ? _slots_6_io_out_uop_bp_debug_if : _slots_5_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_33 ? _slots_8_io_out_uop_bp_xcpt_if : _GEN_32 ? _slots_7_io_out_uop_bp_xcpt_if : _GEN_31 ? _slots_6_io_out_uop_bp_xcpt_if : _slots_5_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_33 ? _slots_8_io_out_uop_debug_fsrc : _GEN_32 ? _slots_7_io_out_uop_debug_fsrc : _GEN_31 ? _slots_6_io_out_uop_debug_fsrc : _slots_5_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_33 ? _slots_8_io_out_uop_debug_tsrc : _GEN_32 ? _slots_7_io_out_uop_debug_tsrc : _GEN_31 ? _slots_6_io_out_uop_debug_tsrc : _slots_5_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_4_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_4_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_4_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_4_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_4_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_4_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_4_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_4_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_4_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_4_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_4_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_4_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_4_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_4_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_4_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_4_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_4_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_4_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_4_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_4_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_4_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_4_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_4_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_4_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_4_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_4_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_4_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_4_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_4_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_4_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_4_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_4_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_4_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_4_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_4_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_4_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_4_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_4_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_4_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_4_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_4_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_4_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_4_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_4_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_4_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_4_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_4_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_4_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_4_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_4_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_4_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_4_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_4_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_4_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_4_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_4_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_4_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_4_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_4_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_4_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_4_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_4_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_4_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_4_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_4_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_4_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_4_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_4_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_4_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_4_io_uop_uopc),
    .io_uop_inst                    (_slots_4_io_uop_inst),
    .io_uop_debug_inst              (_slots_4_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_4_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_4_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_4_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_4_io_uop_fu_code),
    .io_uop_iw_state                (_slots_4_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_4_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_4_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_4_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_4_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_4_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_4_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_4_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_4_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_4_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_4_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_4_io_uop_pc_lob),
    .io_uop_taken                   (_slots_4_io_uop_taken),
    .io_uop_imm_packed              (_slots_4_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_4_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_4_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_4_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_4_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_4_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_4_io_uop_pdst),
    .io_uop_prs1                    (_slots_4_io_uop_prs1),
    .io_uop_prs2                    (_slots_4_io_uop_prs2),
    .io_uop_prs3                    (_slots_4_io_uop_prs3),
    .io_uop_ppred                   (_slots_4_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_4_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_4_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_4_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_4_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_4_io_uop_stale_pdst),
    .io_uop_exception               (_slots_4_io_uop_exception),
    .io_uop_exc_cause               (_slots_4_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_4_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_4_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_4_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_4_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_4_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_4_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_4_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_4_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_4_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_4_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_4_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_4_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_4_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_4_io_uop_ldst),
    .io_uop_lrs1                    (_slots_4_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_4_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_4_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_4_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_4_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_4_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_4_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_4_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_4_io_uop_fp_val),
    .io_uop_fp_single               (_slots_4_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_4_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_4_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_4_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_4_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_4_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_4_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_4_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_5 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_5_io_valid),
    .io_will_be_valid               (_slots_5_io_will_be_valid),
    .io_request                     (_slots_5_io_request),
    .io_grant                       (issue_slots_5_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_4),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_5_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_36 ? _slots_9_io_out_uop_uopc : _GEN_35 ? _slots_8_io_out_uop_uopc : _GEN_34 ? _slots_7_io_out_uop_uopc : _slots_6_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_36 ? _slots_9_io_out_uop_inst : _GEN_35 ? _slots_8_io_out_uop_inst : _GEN_34 ? _slots_7_io_out_uop_inst : _slots_6_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_36 ? _slots_9_io_out_uop_debug_inst : _GEN_35 ? _slots_8_io_out_uop_debug_inst : _GEN_34 ? _slots_7_io_out_uop_debug_inst : _slots_6_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_36 ? _slots_9_io_out_uop_is_rvc : _GEN_35 ? _slots_8_io_out_uop_is_rvc : _GEN_34 ? _slots_7_io_out_uop_is_rvc : _slots_6_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_36 ? _slots_9_io_out_uop_debug_pc : _GEN_35 ? _slots_8_io_out_uop_debug_pc : _GEN_34 ? _slots_7_io_out_uop_debug_pc : _slots_6_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_36 ? _slots_9_io_out_uop_iq_type : _GEN_35 ? _slots_8_io_out_uop_iq_type : _GEN_34 ? _slots_7_io_out_uop_iq_type : _slots_6_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_36 ? _slots_9_io_out_uop_fu_code : _GEN_35 ? _slots_8_io_out_uop_fu_code : _GEN_34 ? _slots_7_io_out_uop_fu_code : _slots_6_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_36 ? _slots_9_io_out_uop_iw_state : _GEN_35 ? _slots_8_io_out_uop_iw_state : _GEN_34 ? _slots_7_io_out_uop_iw_state : _slots_6_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_36 ? _slots_9_io_out_uop_iw_p1_poisoned : _GEN_35 ? _slots_8_io_out_uop_iw_p1_poisoned : _GEN_34 ? _slots_7_io_out_uop_iw_p1_poisoned : _slots_6_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_36 ? _slots_9_io_out_uop_iw_p2_poisoned : _GEN_35 ? _slots_8_io_out_uop_iw_p2_poisoned : _GEN_34 ? _slots_7_io_out_uop_iw_p2_poisoned : _slots_6_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_36 ? _slots_9_io_out_uop_is_br : _GEN_35 ? _slots_8_io_out_uop_is_br : _GEN_34 ? _slots_7_io_out_uop_is_br : _slots_6_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_36 ? _slots_9_io_out_uop_is_jalr : _GEN_35 ? _slots_8_io_out_uop_is_jalr : _GEN_34 ? _slots_7_io_out_uop_is_jalr : _slots_6_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_36 ? _slots_9_io_out_uop_is_jal : _GEN_35 ? _slots_8_io_out_uop_is_jal : _GEN_34 ? _slots_7_io_out_uop_is_jal : _slots_6_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_36 ? _slots_9_io_out_uop_is_sfb : _GEN_35 ? _slots_8_io_out_uop_is_sfb : _GEN_34 ? _slots_7_io_out_uop_is_sfb : _slots_6_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_36 ? _slots_9_io_out_uop_br_mask : _GEN_35 ? _slots_8_io_out_uop_br_mask : _GEN_34 ? _slots_7_io_out_uop_br_mask : _slots_6_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_36 ? _slots_9_io_out_uop_br_tag : _GEN_35 ? _slots_8_io_out_uop_br_tag : _GEN_34 ? _slots_7_io_out_uop_br_tag : _slots_6_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_36 ? _slots_9_io_out_uop_ftq_idx : _GEN_35 ? _slots_8_io_out_uop_ftq_idx : _GEN_34 ? _slots_7_io_out_uop_ftq_idx : _slots_6_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_36 ? _slots_9_io_out_uop_edge_inst : _GEN_35 ? _slots_8_io_out_uop_edge_inst : _GEN_34 ? _slots_7_io_out_uop_edge_inst : _slots_6_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_36 ? _slots_9_io_out_uop_pc_lob : _GEN_35 ? _slots_8_io_out_uop_pc_lob : _GEN_34 ? _slots_7_io_out_uop_pc_lob : _slots_6_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_36 ? _slots_9_io_out_uop_taken : _GEN_35 ? _slots_8_io_out_uop_taken : _GEN_34 ? _slots_7_io_out_uop_taken : _slots_6_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_36 ? _slots_9_io_out_uop_imm_packed : _GEN_35 ? _slots_8_io_out_uop_imm_packed : _GEN_34 ? _slots_7_io_out_uop_imm_packed : _slots_6_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_36 ? _slots_9_io_out_uop_csr_addr : _GEN_35 ? _slots_8_io_out_uop_csr_addr : _GEN_34 ? _slots_7_io_out_uop_csr_addr : _slots_6_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_36 ? _slots_9_io_out_uop_rob_idx : _GEN_35 ? _slots_8_io_out_uop_rob_idx : _GEN_34 ? _slots_7_io_out_uop_rob_idx : _slots_6_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_36 ? _slots_9_io_out_uop_ldq_idx : _GEN_35 ? _slots_8_io_out_uop_ldq_idx : _GEN_34 ? _slots_7_io_out_uop_ldq_idx : _slots_6_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_36 ? _slots_9_io_out_uop_stq_idx : _GEN_35 ? _slots_8_io_out_uop_stq_idx : _GEN_34 ? _slots_7_io_out_uop_stq_idx : _slots_6_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_36 ? _slots_9_io_out_uop_rxq_idx : _GEN_35 ? _slots_8_io_out_uop_rxq_idx : _GEN_34 ? _slots_7_io_out_uop_rxq_idx : _slots_6_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_36 ? _slots_9_io_out_uop_pdst : _GEN_35 ? _slots_8_io_out_uop_pdst : _GEN_34 ? _slots_7_io_out_uop_pdst : _slots_6_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_36 ? _slots_9_io_out_uop_prs1 : _GEN_35 ? _slots_8_io_out_uop_prs1 : _GEN_34 ? _slots_7_io_out_uop_prs1 : _slots_6_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_36 ? _slots_9_io_out_uop_prs2 : _GEN_35 ? _slots_8_io_out_uop_prs2 : _GEN_34 ? _slots_7_io_out_uop_prs2 : _slots_6_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_36 ? _slots_9_io_out_uop_prs3 : _GEN_35 ? _slots_8_io_out_uop_prs3 : _GEN_34 ? _slots_7_io_out_uop_prs3 : _slots_6_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_36 ? _slots_9_io_out_uop_ppred : _GEN_35 ? _slots_8_io_out_uop_ppred : _GEN_34 ? _slots_7_io_out_uop_ppred : _slots_6_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_36 ? _slots_9_io_out_uop_prs1_busy : _GEN_35 ? _slots_8_io_out_uop_prs1_busy : _GEN_34 ? _slots_7_io_out_uop_prs1_busy : _slots_6_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_36 ? _slots_9_io_out_uop_prs2_busy : _GEN_35 ? _slots_8_io_out_uop_prs2_busy : _GEN_34 ? _slots_7_io_out_uop_prs2_busy : _slots_6_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_36 ? _slots_9_io_out_uop_prs3_busy : _GEN_35 ? _slots_8_io_out_uop_prs3_busy : _GEN_34 ? _slots_7_io_out_uop_prs3_busy : _slots_6_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_36 ? _slots_9_io_out_uop_ppred_busy : _GEN_35 ? _slots_8_io_out_uop_ppred_busy : _GEN_34 ? _slots_7_io_out_uop_ppred_busy : _slots_6_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_36 ? _slots_9_io_out_uop_stale_pdst : _GEN_35 ? _slots_8_io_out_uop_stale_pdst : _GEN_34 ? _slots_7_io_out_uop_stale_pdst : _slots_6_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_36 ? _slots_9_io_out_uop_exception : _GEN_35 ? _slots_8_io_out_uop_exception : _GEN_34 ? _slots_7_io_out_uop_exception : _slots_6_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_36 ? _slots_9_io_out_uop_exc_cause : _GEN_35 ? _slots_8_io_out_uop_exc_cause : _GEN_34 ? _slots_7_io_out_uop_exc_cause : _slots_6_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_36 ? _slots_9_io_out_uop_bypassable : _GEN_35 ? _slots_8_io_out_uop_bypassable : _GEN_34 ? _slots_7_io_out_uop_bypassable : _slots_6_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_36 ? _slots_9_io_out_uop_mem_cmd : _GEN_35 ? _slots_8_io_out_uop_mem_cmd : _GEN_34 ? _slots_7_io_out_uop_mem_cmd : _slots_6_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_36 ? _slots_9_io_out_uop_mem_size : _GEN_35 ? _slots_8_io_out_uop_mem_size : _GEN_34 ? _slots_7_io_out_uop_mem_size : _slots_6_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_36 ? _slots_9_io_out_uop_mem_signed : _GEN_35 ? _slots_8_io_out_uop_mem_signed : _GEN_34 ? _slots_7_io_out_uop_mem_signed : _slots_6_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_36 ? _slots_9_io_out_uop_is_fence : _GEN_35 ? _slots_8_io_out_uop_is_fence : _GEN_34 ? _slots_7_io_out_uop_is_fence : _slots_6_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_36 ? _slots_9_io_out_uop_is_fencei : _GEN_35 ? _slots_8_io_out_uop_is_fencei : _GEN_34 ? _slots_7_io_out_uop_is_fencei : _slots_6_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_36 ? _slots_9_io_out_uop_is_amo : _GEN_35 ? _slots_8_io_out_uop_is_amo : _GEN_34 ? _slots_7_io_out_uop_is_amo : _slots_6_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_36 ? _slots_9_io_out_uop_uses_ldq : _GEN_35 ? _slots_8_io_out_uop_uses_ldq : _GEN_34 ? _slots_7_io_out_uop_uses_ldq : _slots_6_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_36 ? _slots_9_io_out_uop_uses_stq : _GEN_35 ? _slots_8_io_out_uop_uses_stq : _GEN_34 ? _slots_7_io_out_uop_uses_stq : _slots_6_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_36 ? _slots_9_io_out_uop_is_sys_pc2epc : _GEN_35 ? _slots_8_io_out_uop_is_sys_pc2epc : _GEN_34 ? _slots_7_io_out_uop_is_sys_pc2epc : _slots_6_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_36 ? _slots_9_io_out_uop_is_unique : _GEN_35 ? _slots_8_io_out_uop_is_unique : _GEN_34 ? _slots_7_io_out_uop_is_unique : _slots_6_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_36 ? _slots_9_io_out_uop_flush_on_commit : _GEN_35 ? _slots_8_io_out_uop_flush_on_commit : _GEN_34 ? _slots_7_io_out_uop_flush_on_commit : _slots_6_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_36 ? _slots_9_io_out_uop_ldst_is_rs1 : _GEN_35 ? _slots_8_io_out_uop_ldst_is_rs1 : _GEN_34 ? _slots_7_io_out_uop_ldst_is_rs1 : _slots_6_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_36 ? _slots_9_io_out_uop_ldst : _GEN_35 ? _slots_8_io_out_uop_ldst : _GEN_34 ? _slots_7_io_out_uop_ldst : _slots_6_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_36 ? _slots_9_io_out_uop_lrs1 : _GEN_35 ? _slots_8_io_out_uop_lrs1 : _GEN_34 ? _slots_7_io_out_uop_lrs1 : _slots_6_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_36 ? _slots_9_io_out_uop_lrs2 : _GEN_35 ? _slots_8_io_out_uop_lrs2 : _GEN_34 ? _slots_7_io_out_uop_lrs2 : _slots_6_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_36 ? _slots_9_io_out_uop_lrs3 : _GEN_35 ? _slots_8_io_out_uop_lrs3 : _GEN_34 ? _slots_7_io_out_uop_lrs3 : _slots_6_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_36 ? _slots_9_io_out_uop_ldst_val : _GEN_35 ? _slots_8_io_out_uop_ldst_val : _GEN_34 ? _slots_7_io_out_uop_ldst_val : _slots_6_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_36 ? _slots_9_io_out_uop_dst_rtype : _GEN_35 ? _slots_8_io_out_uop_dst_rtype : _GEN_34 ? _slots_7_io_out_uop_dst_rtype : _slots_6_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_36 ? _slots_9_io_out_uop_lrs1_rtype : _GEN_35 ? _slots_8_io_out_uop_lrs1_rtype : _GEN_34 ? _slots_7_io_out_uop_lrs1_rtype : _slots_6_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_36 ? _slots_9_io_out_uop_lrs2_rtype : _GEN_35 ? _slots_8_io_out_uop_lrs2_rtype : _GEN_34 ? _slots_7_io_out_uop_lrs2_rtype : _slots_6_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_36 ? _slots_9_io_out_uop_frs3_en : _GEN_35 ? _slots_8_io_out_uop_frs3_en : _GEN_34 ? _slots_7_io_out_uop_frs3_en : _slots_6_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_36 ? _slots_9_io_out_uop_fp_val : _GEN_35 ? _slots_8_io_out_uop_fp_val : _GEN_34 ? _slots_7_io_out_uop_fp_val : _slots_6_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_36 ? _slots_9_io_out_uop_fp_single : _GEN_35 ? _slots_8_io_out_uop_fp_single : _GEN_34 ? _slots_7_io_out_uop_fp_single : _slots_6_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_36 ? _slots_9_io_out_uop_xcpt_pf_if : _GEN_35 ? _slots_8_io_out_uop_xcpt_pf_if : _GEN_34 ? _slots_7_io_out_uop_xcpt_pf_if : _slots_6_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_36 ? _slots_9_io_out_uop_xcpt_ae_if : _GEN_35 ? _slots_8_io_out_uop_xcpt_ae_if : _GEN_34 ? _slots_7_io_out_uop_xcpt_ae_if : _slots_6_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_36 ? _slots_9_io_out_uop_xcpt_ma_if : _GEN_35 ? _slots_8_io_out_uop_xcpt_ma_if : _GEN_34 ? _slots_7_io_out_uop_xcpt_ma_if : _slots_6_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_36 ? _slots_9_io_out_uop_bp_debug_if : _GEN_35 ? _slots_8_io_out_uop_bp_debug_if : _GEN_34 ? _slots_7_io_out_uop_bp_debug_if : _slots_6_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_36 ? _slots_9_io_out_uop_bp_xcpt_if : _GEN_35 ? _slots_8_io_out_uop_bp_xcpt_if : _GEN_34 ? _slots_7_io_out_uop_bp_xcpt_if : _slots_6_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_36 ? _slots_9_io_out_uop_debug_fsrc : _GEN_35 ? _slots_8_io_out_uop_debug_fsrc : _GEN_34 ? _slots_7_io_out_uop_debug_fsrc : _slots_6_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_36 ? _slots_9_io_out_uop_debug_tsrc : _GEN_35 ? _slots_8_io_out_uop_debug_tsrc : _GEN_34 ? _slots_7_io_out_uop_debug_tsrc : _slots_6_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_5_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_5_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_5_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_5_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_5_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_5_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_5_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_5_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_5_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_5_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_5_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_5_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_5_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_5_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_5_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_5_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_5_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_5_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_5_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_5_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_5_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_5_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_5_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_5_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_5_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_5_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_5_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_5_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_5_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_5_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_5_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_5_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_5_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_5_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_5_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_5_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_5_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_5_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_5_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_5_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_5_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_5_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_5_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_5_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_5_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_5_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_5_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_5_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_5_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_5_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_5_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_5_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_5_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_5_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_5_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_5_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_5_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_5_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_5_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_5_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_5_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_5_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_5_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_5_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_5_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_5_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_5_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_5_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_5_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_5_io_uop_uopc),
    .io_uop_inst                    (_slots_5_io_uop_inst),
    .io_uop_debug_inst              (_slots_5_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_5_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_5_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_5_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_5_io_uop_fu_code),
    .io_uop_iw_state                (_slots_5_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_5_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_5_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_5_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_5_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_5_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_5_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_5_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_5_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_5_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_5_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_5_io_uop_pc_lob),
    .io_uop_taken                   (_slots_5_io_uop_taken),
    .io_uop_imm_packed              (_slots_5_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_5_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_5_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_5_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_5_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_5_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_5_io_uop_pdst),
    .io_uop_prs1                    (_slots_5_io_uop_prs1),
    .io_uop_prs2                    (_slots_5_io_uop_prs2),
    .io_uop_prs3                    (_slots_5_io_uop_prs3),
    .io_uop_ppred                   (_slots_5_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_5_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_5_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_5_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_5_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_5_io_uop_stale_pdst),
    .io_uop_exception               (_slots_5_io_uop_exception),
    .io_uop_exc_cause               (_slots_5_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_5_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_5_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_5_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_5_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_5_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_5_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_5_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_5_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_5_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_5_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_5_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_5_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_5_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_5_io_uop_ldst),
    .io_uop_lrs1                    (_slots_5_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_5_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_5_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_5_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_5_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_5_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_5_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_5_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_5_io_uop_fp_val),
    .io_uop_fp_single               (_slots_5_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_5_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_5_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_5_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_5_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_5_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_5_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_5_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_6 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_6_io_valid),
    .io_will_be_valid               (_slots_6_io_will_be_valid),
    .io_request                     (_slots_6_io_request),
    .io_grant                       (issue_slots_6_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_5),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_6_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_39 ? _slots_10_io_out_uop_uopc : _GEN_38 ? _slots_9_io_out_uop_uopc : _GEN_37 ? _slots_8_io_out_uop_uopc : _slots_7_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_39 ? _slots_10_io_out_uop_inst : _GEN_38 ? _slots_9_io_out_uop_inst : _GEN_37 ? _slots_8_io_out_uop_inst : _slots_7_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_39 ? _slots_10_io_out_uop_debug_inst : _GEN_38 ? _slots_9_io_out_uop_debug_inst : _GEN_37 ? _slots_8_io_out_uop_debug_inst : _slots_7_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_39 ? _slots_10_io_out_uop_is_rvc : _GEN_38 ? _slots_9_io_out_uop_is_rvc : _GEN_37 ? _slots_8_io_out_uop_is_rvc : _slots_7_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_39 ? _slots_10_io_out_uop_debug_pc : _GEN_38 ? _slots_9_io_out_uop_debug_pc : _GEN_37 ? _slots_8_io_out_uop_debug_pc : _slots_7_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_39 ? _slots_10_io_out_uop_iq_type : _GEN_38 ? _slots_9_io_out_uop_iq_type : _GEN_37 ? _slots_8_io_out_uop_iq_type : _slots_7_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_39 ? _slots_10_io_out_uop_fu_code : _GEN_38 ? _slots_9_io_out_uop_fu_code : _GEN_37 ? _slots_8_io_out_uop_fu_code : _slots_7_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_39 ? _slots_10_io_out_uop_iw_state : _GEN_38 ? _slots_9_io_out_uop_iw_state : _GEN_37 ? _slots_8_io_out_uop_iw_state : _slots_7_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_39 ? _slots_10_io_out_uop_iw_p1_poisoned : _GEN_38 ? _slots_9_io_out_uop_iw_p1_poisoned : _GEN_37 ? _slots_8_io_out_uop_iw_p1_poisoned : _slots_7_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_39 ? _slots_10_io_out_uop_iw_p2_poisoned : _GEN_38 ? _slots_9_io_out_uop_iw_p2_poisoned : _GEN_37 ? _slots_8_io_out_uop_iw_p2_poisoned : _slots_7_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_39 ? _slots_10_io_out_uop_is_br : _GEN_38 ? _slots_9_io_out_uop_is_br : _GEN_37 ? _slots_8_io_out_uop_is_br : _slots_7_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_39 ? _slots_10_io_out_uop_is_jalr : _GEN_38 ? _slots_9_io_out_uop_is_jalr : _GEN_37 ? _slots_8_io_out_uop_is_jalr : _slots_7_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_39 ? _slots_10_io_out_uop_is_jal : _GEN_38 ? _slots_9_io_out_uop_is_jal : _GEN_37 ? _slots_8_io_out_uop_is_jal : _slots_7_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_39 ? _slots_10_io_out_uop_is_sfb : _GEN_38 ? _slots_9_io_out_uop_is_sfb : _GEN_37 ? _slots_8_io_out_uop_is_sfb : _slots_7_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_39 ? _slots_10_io_out_uop_br_mask : _GEN_38 ? _slots_9_io_out_uop_br_mask : _GEN_37 ? _slots_8_io_out_uop_br_mask : _slots_7_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_39 ? _slots_10_io_out_uop_br_tag : _GEN_38 ? _slots_9_io_out_uop_br_tag : _GEN_37 ? _slots_8_io_out_uop_br_tag : _slots_7_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_39 ? _slots_10_io_out_uop_ftq_idx : _GEN_38 ? _slots_9_io_out_uop_ftq_idx : _GEN_37 ? _slots_8_io_out_uop_ftq_idx : _slots_7_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_39 ? _slots_10_io_out_uop_edge_inst : _GEN_38 ? _slots_9_io_out_uop_edge_inst : _GEN_37 ? _slots_8_io_out_uop_edge_inst : _slots_7_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_39 ? _slots_10_io_out_uop_pc_lob : _GEN_38 ? _slots_9_io_out_uop_pc_lob : _GEN_37 ? _slots_8_io_out_uop_pc_lob : _slots_7_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_39 ? _slots_10_io_out_uop_taken : _GEN_38 ? _slots_9_io_out_uop_taken : _GEN_37 ? _slots_8_io_out_uop_taken : _slots_7_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_39 ? _slots_10_io_out_uop_imm_packed : _GEN_38 ? _slots_9_io_out_uop_imm_packed : _GEN_37 ? _slots_8_io_out_uop_imm_packed : _slots_7_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_39 ? _slots_10_io_out_uop_csr_addr : _GEN_38 ? _slots_9_io_out_uop_csr_addr : _GEN_37 ? _slots_8_io_out_uop_csr_addr : _slots_7_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_39 ? _slots_10_io_out_uop_rob_idx : _GEN_38 ? _slots_9_io_out_uop_rob_idx : _GEN_37 ? _slots_8_io_out_uop_rob_idx : _slots_7_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_39 ? _slots_10_io_out_uop_ldq_idx : _GEN_38 ? _slots_9_io_out_uop_ldq_idx : _GEN_37 ? _slots_8_io_out_uop_ldq_idx : _slots_7_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_39 ? _slots_10_io_out_uop_stq_idx : _GEN_38 ? _slots_9_io_out_uop_stq_idx : _GEN_37 ? _slots_8_io_out_uop_stq_idx : _slots_7_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_39 ? _slots_10_io_out_uop_rxq_idx : _GEN_38 ? _slots_9_io_out_uop_rxq_idx : _GEN_37 ? _slots_8_io_out_uop_rxq_idx : _slots_7_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_39 ? _slots_10_io_out_uop_pdst : _GEN_38 ? _slots_9_io_out_uop_pdst : _GEN_37 ? _slots_8_io_out_uop_pdst : _slots_7_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_39 ? _slots_10_io_out_uop_prs1 : _GEN_38 ? _slots_9_io_out_uop_prs1 : _GEN_37 ? _slots_8_io_out_uop_prs1 : _slots_7_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_39 ? _slots_10_io_out_uop_prs2 : _GEN_38 ? _slots_9_io_out_uop_prs2 : _GEN_37 ? _slots_8_io_out_uop_prs2 : _slots_7_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_39 ? _slots_10_io_out_uop_prs3 : _GEN_38 ? _slots_9_io_out_uop_prs3 : _GEN_37 ? _slots_8_io_out_uop_prs3 : _slots_7_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_39 ? _slots_10_io_out_uop_ppred : _GEN_38 ? _slots_9_io_out_uop_ppred : _GEN_37 ? _slots_8_io_out_uop_ppred : _slots_7_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_39 ? _slots_10_io_out_uop_prs1_busy : _GEN_38 ? _slots_9_io_out_uop_prs1_busy : _GEN_37 ? _slots_8_io_out_uop_prs1_busy : _slots_7_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_39 ? _slots_10_io_out_uop_prs2_busy : _GEN_38 ? _slots_9_io_out_uop_prs2_busy : _GEN_37 ? _slots_8_io_out_uop_prs2_busy : _slots_7_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_39 ? _slots_10_io_out_uop_prs3_busy : _GEN_38 ? _slots_9_io_out_uop_prs3_busy : _GEN_37 ? _slots_8_io_out_uop_prs3_busy : _slots_7_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_39 ? _slots_10_io_out_uop_ppred_busy : _GEN_38 ? _slots_9_io_out_uop_ppred_busy : _GEN_37 ? _slots_8_io_out_uop_ppred_busy : _slots_7_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_39 ? _slots_10_io_out_uop_stale_pdst : _GEN_38 ? _slots_9_io_out_uop_stale_pdst : _GEN_37 ? _slots_8_io_out_uop_stale_pdst : _slots_7_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_39 ? _slots_10_io_out_uop_exception : _GEN_38 ? _slots_9_io_out_uop_exception : _GEN_37 ? _slots_8_io_out_uop_exception : _slots_7_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_39 ? _slots_10_io_out_uop_exc_cause : _GEN_38 ? _slots_9_io_out_uop_exc_cause : _GEN_37 ? _slots_8_io_out_uop_exc_cause : _slots_7_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_39 ? _slots_10_io_out_uop_bypassable : _GEN_38 ? _slots_9_io_out_uop_bypassable : _GEN_37 ? _slots_8_io_out_uop_bypassable : _slots_7_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_39 ? _slots_10_io_out_uop_mem_cmd : _GEN_38 ? _slots_9_io_out_uop_mem_cmd : _GEN_37 ? _slots_8_io_out_uop_mem_cmd : _slots_7_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_39 ? _slots_10_io_out_uop_mem_size : _GEN_38 ? _slots_9_io_out_uop_mem_size : _GEN_37 ? _slots_8_io_out_uop_mem_size : _slots_7_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_39 ? _slots_10_io_out_uop_mem_signed : _GEN_38 ? _slots_9_io_out_uop_mem_signed : _GEN_37 ? _slots_8_io_out_uop_mem_signed : _slots_7_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_39 ? _slots_10_io_out_uop_is_fence : _GEN_38 ? _slots_9_io_out_uop_is_fence : _GEN_37 ? _slots_8_io_out_uop_is_fence : _slots_7_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_39 ? _slots_10_io_out_uop_is_fencei : _GEN_38 ? _slots_9_io_out_uop_is_fencei : _GEN_37 ? _slots_8_io_out_uop_is_fencei : _slots_7_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_39 ? _slots_10_io_out_uop_is_amo : _GEN_38 ? _slots_9_io_out_uop_is_amo : _GEN_37 ? _slots_8_io_out_uop_is_amo : _slots_7_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_39 ? _slots_10_io_out_uop_uses_ldq : _GEN_38 ? _slots_9_io_out_uop_uses_ldq : _GEN_37 ? _slots_8_io_out_uop_uses_ldq : _slots_7_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_39 ? _slots_10_io_out_uop_uses_stq : _GEN_38 ? _slots_9_io_out_uop_uses_stq : _GEN_37 ? _slots_8_io_out_uop_uses_stq : _slots_7_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_39 ? _slots_10_io_out_uop_is_sys_pc2epc : _GEN_38 ? _slots_9_io_out_uop_is_sys_pc2epc : _GEN_37 ? _slots_8_io_out_uop_is_sys_pc2epc : _slots_7_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_39 ? _slots_10_io_out_uop_is_unique : _GEN_38 ? _slots_9_io_out_uop_is_unique : _GEN_37 ? _slots_8_io_out_uop_is_unique : _slots_7_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_39 ? _slots_10_io_out_uop_flush_on_commit : _GEN_38 ? _slots_9_io_out_uop_flush_on_commit : _GEN_37 ? _slots_8_io_out_uop_flush_on_commit : _slots_7_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_39 ? _slots_10_io_out_uop_ldst_is_rs1 : _GEN_38 ? _slots_9_io_out_uop_ldst_is_rs1 : _GEN_37 ? _slots_8_io_out_uop_ldst_is_rs1 : _slots_7_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_39 ? _slots_10_io_out_uop_ldst : _GEN_38 ? _slots_9_io_out_uop_ldst : _GEN_37 ? _slots_8_io_out_uop_ldst : _slots_7_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_39 ? _slots_10_io_out_uop_lrs1 : _GEN_38 ? _slots_9_io_out_uop_lrs1 : _GEN_37 ? _slots_8_io_out_uop_lrs1 : _slots_7_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_39 ? _slots_10_io_out_uop_lrs2 : _GEN_38 ? _slots_9_io_out_uop_lrs2 : _GEN_37 ? _slots_8_io_out_uop_lrs2 : _slots_7_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_39 ? _slots_10_io_out_uop_lrs3 : _GEN_38 ? _slots_9_io_out_uop_lrs3 : _GEN_37 ? _slots_8_io_out_uop_lrs3 : _slots_7_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_39 ? _slots_10_io_out_uop_ldst_val : _GEN_38 ? _slots_9_io_out_uop_ldst_val : _GEN_37 ? _slots_8_io_out_uop_ldst_val : _slots_7_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_39 ? _slots_10_io_out_uop_dst_rtype : _GEN_38 ? _slots_9_io_out_uop_dst_rtype : _GEN_37 ? _slots_8_io_out_uop_dst_rtype : _slots_7_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_39 ? _slots_10_io_out_uop_lrs1_rtype : _GEN_38 ? _slots_9_io_out_uop_lrs1_rtype : _GEN_37 ? _slots_8_io_out_uop_lrs1_rtype : _slots_7_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_39 ? _slots_10_io_out_uop_lrs2_rtype : _GEN_38 ? _slots_9_io_out_uop_lrs2_rtype : _GEN_37 ? _slots_8_io_out_uop_lrs2_rtype : _slots_7_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_39 ? _slots_10_io_out_uop_frs3_en : _GEN_38 ? _slots_9_io_out_uop_frs3_en : _GEN_37 ? _slots_8_io_out_uop_frs3_en : _slots_7_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_39 ? _slots_10_io_out_uop_fp_val : _GEN_38 ? _slots_9_io_out_uop_fp_val : _GEN_37 ? _slots_8_io_out_uop_fp_val : _slots_7_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_39 ? _slots_10_io_out_uop_fp_single : _GEN_38 ? _slots_9_io_out_uop_fp_single : _GEN_37 ? _slots_8_io_out_uop_fp_single : _slots_7_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_39 ? _slots_10_io_out_uop_xcpt_pf_if : _GEN_38 ? _slots_9_io_out_uop_xcpt_pf_if : _GEN_37 ? _slots_8_io_out_uop_xcpt_pf_if : _slots_7_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_39 ? _slots_10_io_out_uop_xcpt_ae_if : _GEN_38 ? _slots_9_io_out_uop_xcpt_ae_if : _GEN_37 ? _slots_8_io_out_uop_xcpt_ae_if : _slots_7_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_39 ? _slots_10_io_out_uop_xcpt_ma_if : _GEN_38 ? _slots_9_io_out_uop_xcpt_ma_if : _GEN_37 ? _slots_8_io_out_uop_xcpt_ma_if : _slots_7_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_39 ? _slots_10_io_out_uop_bp_debug_if : _GEN_38 ? _slots_9_io_out_uop_bp_debug_if : _GEN_37 ? _slots_8_io_out_uop_bp_debug_if : _slots_7_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_39 ? _slots_10_io_out_uop_bp_xcpt_if : _GEN_38 ? _slots_9_io_out_uop_bp_xcpt_if : _GEN_37 ? _slots_8_io_out_uop_bp_xcpt_if : _slots_7_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_39 ? _slots_10_io_out_uop_debug_fsrc : _GEN_38 ? _slots_9_io_out_uop_debug_fsrc : _GEN_37 ? _slots_8_io_out_uop_debug_fsrc : _slots_7_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_39 ? _slots_10_io_out_uop_debug_tsrc : _GEN_38 ? _slots_9_io_out_uop_debug_tsrc : _GEN_37 ? _slots_8_io_out_uop_debug_tsrc : _slots_7_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_6_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_6_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_6_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_6_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_6_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_6_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_6_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_6_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_6_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_6_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_6_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_6_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_6_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_6_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_6_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_6_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_6_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_6_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_6_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_6_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_6_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_6_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_6_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_6_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_6_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_6_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_6_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_6_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_6_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_6_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_6_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_6_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_6_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_6_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_6_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_6_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_6_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_6_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_6_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_6_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_6_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_6_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_6_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_6_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_6_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_6_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_6_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_6_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_6_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_6_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_6_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_6_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_6_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_6_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_6_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_6_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_6_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_6_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_6_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_6_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_6_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_6_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_6_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_6_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_6_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_6_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_6_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_6_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_6_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_6_io_uop_uopc),
    .io_uop_inst                    (_slots_6_io_uop_inst),
    .io_uop_debug_inst              (_slots_6_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_6_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_6_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_6_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_6_io_uop_fu_code),
    .io_uop_iw_state                (_slots_6_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_6_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_6_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_6_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_6_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_6_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_6_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_6_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_6_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_6_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_6_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_6_io_uop_pc_lob),
    .io_uop_taken                   (_slots_6_io_uop_taken),
    .io_uop_imm_packed              (_slots_6_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_6_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_6_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_6_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_6_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_6_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_6_io_uop_pdst),
    .io_uop_prs1                    (_slots_6_io_uop_prs1),
    .io_uop_prs2                    (_slots_6_io_uop_prs2),
    .io_uop_prs3                    (_slots_6_io_uop_prs3),
    .io_uop_ppred                   (_slots_6_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_6_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_6_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_6_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_6_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_6_io_uop_stale_pdst),
    .io_uop_exception               (_slots_6_io_uop_exception),
    .io_uop_exc_cause               (_slots_6_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_6_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_6_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_6_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_6_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_6_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_6_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_6_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_6_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_6_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_6_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_6_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_6_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_6_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_6_io_uop_ldst),
    .io_uop_lrs1                    (_slots_6_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_6_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_6_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_6_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_6_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_6_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_6_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_6_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_6_io_uop_fp_val),
    .io_uop_fp_single               (_slots_6_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_6_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_6_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_6_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_6_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_6_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_6_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_6_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_7 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_7_io_valid),
    .io_will_be_valid               (_slots_7_io_will_be_valid),
    .io_request                     (_slots_7_io_request),
    .io_grant                       (issue_slots_7_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_6),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_7_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_42 ? _slots_11_io_out_uop_uopc : _GEN_41 ? _slots_10_io_out_uop_uopc : _GEN_40 ? _slots_9_io_out_uop_uopc : _slots_8_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_42 ? _slots_11_io_out_uop_inst : _GEN_41 ? _slots_10_io_out_uop_inst : _GEN_40 ? _slots_9_io_out_uop_inst : _slots_8_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_42 ? _slots_11_io_out_uop_debug_inst : _GEN_41 ? _slots_10_io_out_uop_debug_inst : _GEN_40 ? _slots_9_io_out_uop_debug_inst : _slots_8_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_42 ? _slots_11_io_out_uop_is_rvc : _GEN_41 ? _slots_10_io_out_uop_is_rvc : _GEN_40 ? _slots_9_io_out_uop_is_rvc : _slots_8_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_42 ? _slots_11_io_out_uop_debug_pc : _GEN_41 ? _slots_10_io_out_uop_debug_pc : _GEN_40 ? _slots_9_io_out_uop_debug_pc : _slots_8_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_42 ? _slots_11_io_out_uop_iq_type : _GEN_41 ? _slots_10_io_out_uop_iq_type : _GEN_40 ? _slots_9_io_out_uop_iq_type : _slots_8_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_42 ? _slots_11_io_out_uop_fu_code : _GEN_41 ? _slots_10_io_out_uop_fu_code : _GEN_40 ? _slots_9_io_out_uop_fu_code : _slots_8_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_42 ? _slots_11_io_out_uop_iw_state : _GEN_41 ? _slots_10_io_out_uop_iw_state : _GEN_40 ? _slots_9_io_out_uop_iw_state : _slots_8_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_42 ? _slots_11_io_out_uop_iw_p1_poisoned : _GEN_41 ? _slots_10_io_out_uop_iw_p1_poisoned : _GEN_40 ? _slots_9_io_out_uop_iw_p1_poisoned : _slots_8_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_42 ? _slots_11_io_out_uop_iw_p2_poisoned : _GEN_41 ? _slots_10_io_out_uop_iw_p2_poisoned : _GEN_40 ? _slots_9_io_out_uop_iw_p2_poisoned : _slots_8_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_42 ? _slots_11_io_out_uop_is_br : _GEN_41 ? _slots_10_io_out_uop_is_br : _GEN_40 ? _slots_9_io_out_uop_is_br : _slots_8_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_42 ? _slots_11_io_out_uop_is_jalr : _GEN_41 ? _slots_10_io_out_uop_is_jalr : _GEN_40 ? _slots_9_io_out_uop_is_jalr : _slots_8_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_42 ? _slots_11_io_out_uop_is_jal : _GEN_41 ? _slots_10_io_out_uop_is_jal : _GEN_40 ? _slots_9_io_out_uop_is_jal : _slots_8_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_42 ? _slots_11_io_out_uop_is_sfb : _GEN_41 ? _slots_10_io_out_uop_is_sfb : _GEN_40 ? _slots_9_io_out_uop_is_sfb : _slots_8_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_42 ? _slots_11_io_out_uop_br_mask : _GEN_41 ? _slots_10_io_out_uop_br_mask : _GEN_40 ? _slots_9_io_out_uop_br_mask : _slots_8_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_42 ? _slots_11_io_out_uop_br_tag : _GEN_41 ? _slots_10_io_out_uop_br_tag : _GEN_40 ? _slots_9_io_out_uop_br_tag : _slots_8_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_42 ? _slots_11_io_out_uop_ftq_idx : _GEN_41 ? _slots_10_io_out_uop_ftq_idx : _GEN_40 ? _slots_9_io_out_uop_ftq_idx : _slots_8_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_42 ? _slots_11_io_out_uop_edge_inst : _GEN_41 ? _slots_10_io_out_uop_edge_inst : _GEN_40 ? _slots_9_io_out_uop_edge_inst : _slots_8_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_42 ? _slots_11_io_out_uop_pc_lob : _GEN_41 ? _slots_10_io_out_uop_pc_lob : _GEN_40 ? _slots_9_io_out_uop_pc_lob : _slots_8_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_42 ? _slots_11_io_out_uop_taken : _GEN_41 ? _slots_10_io_out_uop_taken : _GEN_40 ? _slots_9_io_out_uop_taken : _slots_8_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_42 ? _slots_11_io_out_uop_imm_packed : _GEN_41 ? _slots_10_io_out_uop_imm_packed : _GEN_40 ? _slots_9_io_out_uop_imm_packed : _slots_8_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_42 ? _slots_11_io_out_uop_csr_addr : _GEN_41 ? _slots_10_io_out_uop_csr_addr : _GEN_40 ? _slots_9_io_out_uop_csr_addr : _slots_8_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_42 ? _slots_11_io_out_uop_rob_idx : _GEN_41 ? _slots_10_io_out_uop_rob_idx : _GEN_40 ? _slots_9_io_out_uop_rob_idx : _slots_8_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_42 ? _slots_11_io_out_uop_ldq_idx : _GEN_41 ? _slots_10_io_out_uop_ldq_idx : _GEN_40 ? _slots_9_io_out_uop_ldq_idx : _slots_8_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_42 ? _slots_11_io_out_uop_stq_idx : _GEN_41 ? _slots_10_io_out_uop_stq_idx : _GEN_40 ? _slots_9_io_out_uop_stq_idx : _slots_8_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_42 ? _slots_11_io_out_uop_rxq_idx : _GEN_41 ? _slots_10_io_out_uop_rxq_idx : _GEN_40 ? _slots_9_io_out_uop_rxq_idx : _slots_8_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_42 ? _slots_11_io_out_uop_pdst : _GEN_41 ? _slots_10_io_out_uop_pdst : _GEN_40 ? _slots_9_io_out_uop_pdst : _slots_8_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_42 ? _slots_11_io_out_uop_prs1 : _GEN_41 ? _slots_10_io_out_uop_prs1 : _GEN_40 ? _slots_9_io_out_uop_prs1 : _slots_8_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_42 ? _slots_11_io_out_uop_prs2 : _GEN_41 ? _slots_10_io_out_uop_prs2 : _GEN_40 ? _slots_9_io_out_uop_prs2 : _slots_8_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_42 ? _slots_11_io_out_uop_prs3 : _GEN_41 ? _slots_10_io_out_uop_prs3 : _GEN_40 ? _slots_9_io_out_uop_prs3 : _slots_8_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_42 ? _slots_11_io_out_uop_ppred : _GEN_41 ? _slots_10_io_out_uop_ppred : _GEN_40 ? _slots_9_io_out_uop_ppred : _slots_8_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_42 ? _slots_11_io_out_uop_prs1_busy : _GEN_41 ? _slots_10_io_out_uop_prs1_busy : _GEN_40 ? _slots_9_io_out_uop_prs1_busy : _slots_8_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_42 ? _slots_11_io_out_uop_prs2_busy : _GEN_41 ? _slots_10_io_out_uop_prs2_busy : _GEN_40 ? _slots_9_io_out_uop_prs2_busy : _slots_8_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_42 ? _slots_11_io_out_uop_prs3_busy : _GEN_41 ? _slots_10_io_out_uop_prs3_busy : _GEN_40 ? _slots_9_io_out_uop_prs3_busy : _slots_8_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_42 ? _slots_11_io_out_uop_ppred_busy : _GEN_41 ? _slots_10_io_out_uop_ppred_busy : _GEN_40 ? _slots_9_io_out_uop_ppred_busy : _slots_8_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_42 ? _slots_11_io_out_uop_stale_pdst : _GEN_41 ? _slots_10_io_out_uop_stale_pdst : _GEN_40 ? _slots_9_io_out_uop_stale_pdst : _slots_8_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_42 ? _slots_11_io_out_uop_exception : _GEN_41 ? _slots_10_io_out_uop_exception : _GEN_40 ? _slots_9_io_out_uop_exception : _slots_8_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_42 ? _slots_11_io_out_uop_exc_cause : _GEN_41 ? _slots_10_io_out_uop_exc_cause : _GEN_40 ? _slots_9_io_out_uop_exc_cause : _slots_8_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_42 ? _slots_11_io_out_uop_bypassable : _GEN_41 ? _slots_10_io_out_uop_bypassable : _GEN_40 ? _slots_9_io_out_uop_bypassable : _slots_8_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_42 ? _slots_11_io_out_uop_mem_cmd : _GEN_41 ? _slots_10_io_out_uop_mem_cmd : _GEN_40 ? _slots_9_io_out_uop_mem_cmd : _slots_8_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_42 ? _slots_11_io_out_uop_mem_size : _GEN_41 ? _slots_10_io_out_uop_mem_size : _GEN_40 ? _slots_9_io_out_uop_mem_size : _slots_8_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_42 ? _slots_11_io_out_uop_mem_signed : _GEN_41 ? _slots_10_io_out_uop_mem_signed : _GEN_40 ? _slots_9_io_out_uop_mem_signed : _slots_8_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_42 ? _slots_11_io_out_uop_is_fence : _GEN_41 ? _slots_10_io_out_uop_is_fence : _GEN_40 ? _slots_9_io_out_uop_is_fence : _slots_8_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_42 ? _slots_11_io_out_uop_is_fencei : _GEN_41 ? _slots_10_io_out_uop_is_fencei : _GEN_40 ? _slots_9_io_out_uop_is_fencei : _slots_8_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_42 ? _slots_11_io_out_uop_is_amo : _GEN_41 ? _slots_10_io_out_uop_is_amo : _GEN_40 ? _slots_9_io_out_uop_is_amo : _slots_8_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_42 ? _slots_11_io_out_uop_uses_ldq : _GEN_41 ? _slots_10_io_out_uop_uses_ldq : _GEN_40 ? _slots_9_io_out_uop_uses_ldq : _slots_8_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_42 ? _slots_11_io_out_uop_uses_stq : _GEN_41 ? _slots_10_io_out_uop_uses_stq : _GEN_40 ? _slots_9_io_out_uop_uses_stq : _slots_8_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_42 ? _slots_11_io_out_uop_is_sys_pc2epc : _GEN_41 ? _slots_10_io_out_uop_is_sys_pc2epc : _GEN_40 ? _slots_9_io_out_uop_is_sys_pc2epc : _slots_8_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_42 ? _slots_11_io_out_uop_is_unique : _GEN_41 ? _slots_10_io_out_uop_is_unique : _GEN_40 ? _slots_9_io_out_uop_is_unique : _slots_8_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_42 ? _slots_11_io_out_uop_flush_on_commit : _GEN_41 ? _slots_10_io_out_uop_flush_on_commit : _GEN_40 ? _slots_9_io_out_uop_flush_on_commit : _slots_8_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_42 ? _slots_11_io_out_uop_ldst_is_rs1 : _GEN_41 ? _slots_10_io_out_uop_ldst_is_rs1 : _GEN_40 ? _slots_9_io_out_uop_ldst_is_rs1 : _slots_8_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_42 ? _slots_11_io_out_uop_ldst : _GEN_41 ? _slots_10_io_out_uop_ldst : _GEN_40 ? _slots_9_io_out_uop_ldst : _slots_8_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_42 ? _slots_11_io_out_uop_lrs1 : _GEN_41 ? _slots_10_io_out_uop_lrs1 : _GEN_40 ? _slots_9_io_out_uop_lrs1 : _slots_8_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_42 ? _slots_11_io_out_uop_lrs2 : _GEN_41 ? _slots_10_io_out_uop_lrs2 : _GEN_40 ? _slots_9_io_out_uop_lrs2 : _slots_8_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_42 ? _slots_11_io_out_uop_lrs3 : _GEN_41 ? _slots_10_io_out_uop_lrs3 : _GEN_40 ? _slots_9_io_out_uop_lrs3 : _slots_8_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_42 ? _slots_11_io_out_uop_ldst_val : _GEN_41 ? _slots_10_io_out_uop_ldst_val : _GEN_40 ? _slots_9_io_out_uop_ldst_val : _slots_8_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_42 ? _slots_11_io_out_uop_dst_rtype : _GEN_41 ? _slots_10_io_out_uop_dst_rtype : _GEN_40 ? _slots_9_io_out_uop_dst_rtype : _slots_8_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_42 ? _slots_11_io_out_uop_lrs1_rtype : _GEN_41 ? _slots_10_io_out_uop_lrs1_rtype : _GEN_40 ? _slots_9_io_out_uop_lrs1_rtype : _slots_8_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_42 ? _slots_11_io_out_uop_lrs2_rtype : _GEN_41 ? _slots_10_io_out_uop_lrs2_rtype : _GEN_40 ? _slots_9_io_out_uop_lrs2_rtype : _slots_8_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_42 ? _slots_11_io_out_uop_frs3_en : _GEN_41 ? _slots_10_io_out_uop_frs3_en : _GEN_40 ? _slots_9_io_out_uop_frs3_en : _slots_8_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_42 ? _slots_11_io_out_uop_fp_val : _GEN_41 ? _slots_10_io_out_uop_fp_val : _GEN_40 ? _slots_9_io_out_uop_fp_val : _slots_8_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_42 ? _slots_11_io_out_uop_fp_single : _GEN_41 ? _slots_10_io_out_uop_fp_single : _GEN_40 ? _slots_9_io_out_uop_fp_single : _slots_8_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_42 ? _slots_11_io_out_uop_xcpt_pf_if : _GEN_41 ? _slots_10_io_out_uop_xcpt_pf_if : _GEN_40 ? _slots_9_io_out_uop_xcpt_pf_if : _slots_8_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_42 ? _slots_11_io_out_uop_xcpt_ae_if : _GEN_41 ? _slots_10_io_out_uop_xcpt_ae_if : _GEN_40 ? _slots_9_io_out_uop_xcpt_ae_if : _slots_8_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_42 ? _slots_11_io_out_uop_xcpt_ma_if : _GEN_41 ? _slots_10_io_out_uop_xcpt_ma_if : _GEN_40 ? _slots_9_io_out_uop_xcpt_ma_if : _slots_8_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_42 ? _slots_11_io_out_uop_bp_debug_if : _GEN_41 ? _slots_10_io_out_uop_bp_debug_if : _GEN_40 ? _slots_9_io_out_uop_bp_debug_if : _slots_8_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_42 ? _slots_11_io_out_uop_bp_xcpt_if : _GEN_41 ? _slots_10_io_out_uop_bp_xcpt_if : _GEN_40 ? _slots_9_io_out_uop_bp_xcpt_if : _slots_8_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_42 ? _slots_11_io_out_uop_debug_fsrc : _GEN_41 ? _slots_10_io_out_uop_debug_fsrc : _GEN_40 ? _slots_9_io_out_uop_debug_fsrc : _slots_8_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_42 ? _slots_11_io_out_uop_debug_tsrc : _GEN_41 ? _slots_10_io_out_uop_debug_tsrc : _GEN_40 ? _slots_9_io_out_uop_debug_tsrc : _slots_8_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_7_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_7_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_7_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_7_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_7_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_7_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_7_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_7_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_7_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_7_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_7_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_7_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_7_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_7_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_7_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_7_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_7_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_7_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_7_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_7_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_7_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_7_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_7_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_7_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_7_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_7_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_7_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_7_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_7_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_7_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_7_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_7_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_7_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_7_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_7_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_7_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_7_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_7_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_7_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_7_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_7_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_7_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_7_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_7_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_7_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_7_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_7_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_7_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_7_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_7_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_7_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_7_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_7_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_7_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_7_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_7_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_7_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_7_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_7_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_7_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_7_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_7_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_7_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_7_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_7_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_7_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_7_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_7_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_7_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_7_io_uop_uopc),
    .io_uop_inst                    (_slots_7_io_uop_inst),
    .io_uop_debug_inst              (_slots_7_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_7_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_7_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_7_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_7_io_uop_fu_code),
    .io_uop_iw_state                (_slots_7_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_7_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_7_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_7_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_7_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_7_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_7_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_7_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_7_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_7_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_7_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_7_io_uop_pc_lob),
    .io_uop_taken                   (_slots_7_io_uop_taken),
    .io_uop_imm_packed              (_slots_7_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_7_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_7_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_7_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_7_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_7_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_7_io_uop_pdst),
    .io_uop_prs1                    (_slots_7_io_uop_prs1),
    .io_uop_prs2                    (_slots_7_io_uop_prs2),
    .io_uop_prs3                    (_slots_7_io_uop_prs3),
    .io_uop_ppred                   (_slots_7_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_7_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_7_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_7_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_7_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_7_io_uop_stale_pdst),
    .io_uop_exception               (_slots_7_io_uop_exception),
    .io_uop_exc_cause               (_slots_7_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_7_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_7_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_7_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_7_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_7_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_7_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_7_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_7_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_7_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_7_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_7_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_7_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_7_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_7_io_uop_ldst),
    .io_uop_lrs1                    (_slots_7_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_7_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_7_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_7_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_7_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_7_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_7_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_7_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_7_io_uop_fp_val),
    .io_uop_fp_single               (_slots_7_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_7_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_7_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_7_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_7_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_7_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_7_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_7_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_8 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_8_io_valid),
    .io_will_be_valid               (_slots_8_io_will_be_valid),
    .io_request                     (_slots_8_io_request),
    .io_grant                       (issue_slots_8_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_7),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_8_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_45 ? _slots_12_io_out_uop_uopc : _GEN_44 ? _slots_11_io_out_uop_uopc : _GEN_43 ? _slots_10_io_out_uop_uopc : _slots_9_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_45 ? _slots_12_io_out_uop_inst : _GEN_44 ? _slots_11_io_out_uop_inst : _GEN_43 ? _slots_10_io_out_uop_inst : _slots_9_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_45 ? _slots_12_io_out_uop_debug_inst : _GEN_44 ? _slots_11_io_out_uop_debug_inst : _GEN_43 ? _slots_10_io_out_uop_debug_inst : _slots_9_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_45 ? _slots_12_io_out_uop_is_rvc : _GEN_44 ? _slots_11_io_out_uop_is_rvc : _GEN_43 ? _slots_10_io_out_uop_is_rvc : _slots_9_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_45 ? _slots_12_io_out_uop_debug_pc : _GEN_44 ? _slots_11_io_out_uop_debug_pc : _GEN_43 ? _slots_10_io_out_uop_debug_pc : _slots_9_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_45 ? _slots_12_io_out_uop_iq_type : _GEN_44 ? _slots_11_io_out_uop_iq_type : _GEN_43 ? _slots_10_io_out_uop_iq_type : _slots_9_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_45 ? _slots_12_io_out_uop_fu_code : _GEN_44 ? _slots_11_io_out_uop_fu_code : _GEN_43 ? _slots_10_io_out_uop_fu_code : _slots_9_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_45 ? _slots_12_io_out_uop_iw_state : _GEN_44 ? _slots_11_io_out_uop_iw_state : _GEN_43 ? _slots_10_io_out_uop_iw_state : _slots_9_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_45 ? _slots_12_io_out_uop_iw_p1_poisoned : _GEN_44 ? _slots_11_io_out_uop_iw_p1_poisoned : _GEN_43 ? _slots_10_io_out_uop_iw_p1_poisoned : _slots_9_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_45 ? _slots_12_io_out_uop_iw_p2_poisoned : _GEN_44 ? _slots_11_io_out_uop_iw_p2_poisoned : _GEN_43 ? _slots_10_io_out_uop_iw_p2_poisoned : _slots_9_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_45 ? _slots_12_io_out_uop_is_br : _GEN_44 ? _slots_11_io_out_uop_is_br : _GEN_43 ? _slots_10_io_out_uop_is_br : _slots_9_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_45 ? _slots_12_io_out_uop_is_jalr : _GEN_44 ? _slots_11_io_out_uop_is_jalr : _GEN_43 ? _slots_10_io_out_uop_is_jalr : _slots_9_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_45 ? _slots_12_io_out_uop_is_jal : _GEN_44 ? _slots_11_io_out_uop_is_jal : _GEN_43 ? _slots_10_io_out_uop_is_jal : _slots_9_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_45 ? _slots_12_io_out_uop_is_sfb : _GEN_44 ? _slots_11_io_out_uop_is_sfb : _GEN_43 ? _slots_10_io_out_uop_is_sfb : _slots_9_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_45 ? _slots_12_io_out_uop_br_mask : _GEN_44 ? _slots_11_io_out_uop_br_mask : _GEN_43 ? _slots_10_io_out_uop_br_mask : _slots_9_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_45 ? _slots_12_io_out_uop_br_tag : _GEN_44 ? _slots_11_io_out_uop_br_tag : _GEN_43 ? _slots_10_io_out_uop_br_tag : _slots_9_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_45 ? _slots_12_io_out_uop_ftq_idx : _GEN_44 ? _slots_11_io_out_uop_ftq_idx : _GEN_43 ? _slots_10_io_out_uop_ftq_idx : _slots_9_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_45 ? _slots_12_io_out_uop_edge_inst : _GEN_44 ? _slots_11_io_out_uop_edge_inst : _GEN_43 ? _slots_10_io_out_uop_edge_inst : _slots_9_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_45 ? _slots_12_io_out_uop_pc_lob : _GEN_44 ? _slots_11_io_out_uop_pc_lob : _GEN_43 ? _slots_10_io_out_uop_pc_lob : _slots_9_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_45 ? _slots_12_io_out_uop_taken : _GEN_44 ? _slots_11_io_out_uop_taken : _GEN_43 ? _slots_10_io_out_uop_taken : _slots_9_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_45 ? _slots_12_io_out_uop_imm_packed : _GEN_44 ? _slots_11_io_out_uop_imm_packed : _GEN_43 ? _slots_10_io_out_uop_imm_packed : _slots_9_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_45 ? _slots_12_io_out_uop_csr_addr : _GEN_44 ? _slots_11_io_out_uop_csr_addr : _GEN_43 ? _slots_10_io_out_uop_csr_addr : _slots_9_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_45 ? _slots_12_io_out_uop_rob_idx : _GEN_44 ? _slots_11_io_out_uop_rob_idx : _GEN_43 ? _slots_10_io_out_uop_rob_idx : _slots_9_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_45 ? _slots_12_io_out_uop_ldq_idx : _GEN_44 ? _slots_11_io_out_uop_ldq_idx : _GEN_43 ? _slots_10_io_out_uop_ldq_idx : _slots_9_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_45 ? _slots_12_io_out_uop_stq_idx : _GEN_44 ? _slots_11_io_out_uop_stq_idx : _GEN_43 ? _slots_10_io_out_uop_stq_idx : _slots_9_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_45 ? _slots_12_io_out_uop_rxq_idx : _GEN_44 ? _slots_11_io_out_uop_rxq_idx : _GEN_43 ? _slots_10_io_out_uop_rxq_idx : _slots_9_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_45 ? _slots_12_io_out_uop_pdst : _GEN_44 ? _slots_11_io_out_uop_pdst : _GEN_43 ? _slots_10_io_out_uop_pdst : _slots_9_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_45 ? _slots_12_io_out_uop_prs1 : _GEN_44 ? _slots_11_io_out_uop_prs1 : _GEN_43 ? _slots_10_io_out_uop_prs1 : _slots_9_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_45 ? _slots_12_io_out_uop_prs2 : _GEN_44 ? _slots_11_io_out_uop_prs2 : _GEN_43 ? _slots_10_io_out_uop_prs2 : _slots_9_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_45 ? _slots_12_io_out_uop_prs3 : _GEN_44 ? _slots_11_io_out_uop_prs3 : _GEN_43 ? _slots_10_io_out_uop_prs3 : _slots_9_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_45 ? _slots_12_io_out_uop_ppred : _GEN_44 ? _slots_11_io_out_uop_ppred : _GEN_43 ? _slots_10_io_out_uop_ppred : _slots_9_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_45 ? _slots_12_io_out_uop_prs1_busy : _GEN_44 ? _slots_11_io_out_uop_prs1_busy : _GEN_43 ? _slots_10_io_out_uop_prs1_busy : _slots_9_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_45 ? _slots_12_io_out_uop_prs2_busy : _GEN_44 ? _slots_11_io_out_uop_prs2_busy : _GEN_43 ? _slots_10_io_out_uop_prs2_busy : _slots_9_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_45 ? _slots_12_io_out_uop_prs3_busy : _GEN_44 ? _slots_11_io_out_uop_prs3_busy : _GEN_43 ? _slots_10_io_out_uop_prs3_busy : _slots_9_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_45 ? _slots_12_io_out_uop_ppred_busy : _GEN_44 ? _slots_11_io_out_uop_ppred_busy : _GEN_43 ? _slots_10_io_out_uop_ppred_busy : _slots_9_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_45 ? _slots_12_io_out_uop_stale_pdst : _GEN_44 ? _slots_11_io_out_uop_stale_pdst : _GEN_43 ? _slots_10_io_out_uop_stale_pdst : _slots_9_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_45 ? _slots_12_io_out_uop_exception : _GEN_44 ? _slots_11_io_out_uop_exception : _GEN_43 ? _slots_10_io_out_uop_exception : _slots_9_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_45 ? _slots_12_io_out_uop_exc_cause : _GEN_44 ? _slots_11_io_out_uop_exc_cause : _GEN_43 ? _slots_10_io_out_uop_exc_cause : _slots_9_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_45 ? _slots_12_io_out_uop_bypassable : _GEN_44 ? _slots_11_io_out_uop_bypassable : _GEN_43 ? _slots_10_io_out_uop_bypassable : _slots_9_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_45 ? _slots_12_io_out_uop_mem_cmd : _GEN_44 ? _slots_11_io_out_uop_mem_cmd : _GEN_43 ? _slots_10_io_out_uop_mem_cmd : _slots_9_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_45 ? _slots_12_io_out_uop_mem_size : _GEN_44 ? _slots_11_io_out_uop_mem_size : _GEN_43 ? _slots_10_io_out_uop_mem_size : _slots_9_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_45 ? _slots_12_io_out_uop_mem_signed : _GEN_44 ? _slots_11_io_out_uop_mem_signed : _GEN_43 ? _slots_10_io_out_uop_mem_signed : _slots_9_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_45 ? _slots_12_io_out_uop_is_fence : _GEN_44 ? _slots_11_io_out_uop_is_fence : _GEN_43 ? _slots_10_io_out_uop_is_fence : _slots_9_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_45 ? _slots_12_io_out_uop_is_fencei : _GEN_44 ? _slots_11_io_out_uop_is_fencei : _GEN_43 ? _slots_10_io_out_uop_is_fencei : _slots_9_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_45 ? _slots_12_io_out_uop_is_amo : _GEN_44 ? _slots_11_io_out_uop_is_amo : _GEN_43 ? _slots_10_io_out_uop_is_amo : _slots_9_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_45 ? _slots_12_io_out_uop_uses_ldq : _GEN_44 ? _slots_11_io_out_uop_uses_ldq : _GEN_43 ? _slots_10_io_out_uop_uses_ldq : _slots_9_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_45 ? _slots_12_io_out_uop_uses_stq : _GEN_44 ? _slots_11_io_out_uop_uses_stq : _GEN_43 ? _slots_10_io_out_uop_uses_stq : _slots_9_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_45 ? _slots_12_io_out_uop_is_sys_pc2epc : _GEN_44 ? _slots_11_io_out_uop_is_sys_pc2epc : _GEN_43 ? _slots_10_io_out_uop_is_sys_pc2epc : _slots_9_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_45 ? _slots_12_io_out_uop_is_unique : _GEN_44 ? _slots_11_io_out_uop_is_unique : _GEN_43 ? _slots_10_io_out_uop_is_unique : _slots_9_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_45 ? _slots_12_io_out_uop_flush_on_commit : _GEN_44 ? _slots_11_io_out_uop_flush_on_commit : _GEN_43 ? _slots_10_io_out_uop_flush_on_commit : _slots_9_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_45 ? _slots_12_io_out_uop_ldst_is_rs1 : _GEN_44 ? _slots_11_io_out_uop_ldst_is_rs1 : _GEN_43 ? _slots_10_io_out_uop_ldst_is_rs1 : _slots_9_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_45 ? _slots_12_io_out_uop_ldst : _GEN_44 ? _slots_11_io_out_uop_ldst : _GEN_43 ? _slots_10_io_out_uop_ldst : _slots_9_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_45 ? _slots_12_io_out_uop_lrs1 : _GEN_44 ? _slots_11_io_out_uop_lrs1 : _GEN_43 ? _slots_10_io_out_uop_lrs1 : _slots_9_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_45 ? _slots_12_io_out_uop_lrs2 : _GEN_44 ? _slots_11_io_out_uop_lrs2 : _GEN_43 ? _slots_10_io_out_uop_lrs2 : _slots_9_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_45 ? _slots_12_io_out_uop_lrs3 : _GEN_44 ? _slots_11_io_out_uop_lrs3 : _GEN_43 ? _slots_10_io_out_uop_lrs3 : _slots_9_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_45 ? _slots_12_io_out_uop_ldst_val : _GEN_44 ? _slots_11_io_out_uop_ldst_val : _GEN_43 ? _slots_10_io_out_uop_ldst_val : _slots_9_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_45 ? _slots_12_io_out_uop_dst_rtype : _GEN_44 ? _slots_11_io_out_uop_dst_rtype : _GEN_43 ? _slots_10_io_out_uop_dst_rtype : _slots_9_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_45 ? _slots_12_io_out_uop_lrs1_rtype : _GEN_44 ? _slots_11_io_out_uop_lrs1_rtype : _GEN_43 ? _slots_10_io_out_uop_lrs1_rtype : _slots_9_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_45 ? _slots_12_io_out_uop_lrs2_rtype : _GEN_44 ? _slots_11_io_out_uop_lrs2_rtype : _GEN_43 ? _slots_10_io_out_uop_lrs2_rtype : _slots_9_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_45 ? _slots_12_io_out_uop_frs3_en : _GEN_44 ? _slots_11_io_out_uop_frs3_en : _GEN_43 ? _slots_10_io_out_uop_frs3_en : _slots_9_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_45 ? _slots_12_io_out_uop_fp_val : _GEN_44 ? _slots_11_io_out_uop_fp_val : _GEN_43 ? _slots_10_io_out_uop_fp_val : _slots_9_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_45 ? _slots_12_io_out_uop_fp_single : _GEN_44 ? _slots_11_io_out_uop_fp_single : _GEN_43 ? _slots_10_io_out_uop_fp_single : _slots_9_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_45 ? _slots_12_io_out_uop_xcpt_pf_if : _GEN_44 ? _slots_11_io_out_uop_xcpt_pf_if : _GEN_43 ? _slots_10_io_out_uop_xcpt_pf_if : _slots_9_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_45 ? _slots_12_io_out_uop_xcpt_ae_if : _GEN_44 ? _slots_11_io_out_uop_xcpt_ae_if : _GEN_43 ? _slots_10_io_out_uop_xcpt_ae_if : _slots_9_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_45 ? _slots_12_io_out_uop_xcpt_ma_if : _GEN_44 ? _slots_11_io_out_uop_xcpt_ma_if : _GEN_43 ? _slots_10_io_out_uop_xcpt_ma_if : _slots_9_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_45 ? _slots_12_io_out_uop_bp_debug_if : _GEN_44 ? _slots_11_io_out_uop_bp_debug_if : _GEN_43 ? _slots_10_io_out_uop_bp_debug_if : _slots_9_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_45 ? _slots_12_io_out_uop_bp_xcpt_if : _GEN_44 ? _slots_11_io_out_uop_bp_xcpt_if : _GEN_43 ? _slots_10_io_out_uop_bp_xcpt_if : _slots_9_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_45 ? _slots_12_io_out_uop_debug_fsrc : _GEN_44 ? _slots_11_io_out_uop_debug_fsrc : _GEN_43 ? _slots_10_io_out_uop_debug_fsrc : _slots_9_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_45 ? _slots_12_io_out_uop_debug_tsrc : _GEN_44 ? _slots_11_io_out_uop_debug_tsrc : _GEN_43 ? _slots_10_io_out_uop_debug_tsrc : _slots_9_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_8_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_8_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_8_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_8_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_8_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_8_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_8_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_8_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_8_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_8_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_8_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_8_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_8_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_8_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_8_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_8_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_8_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_8_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_8_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_8_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_8_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_8_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_8_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_8_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_8_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_8_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_8_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_8_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_8_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_8_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_8_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_8_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_8_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_8_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_8_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_8_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_8_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_8_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_8_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_8_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_8_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_8_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_8_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_8_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_8_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_8_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_8_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_8_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_8_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_8_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_8_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_8_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_8_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_8_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_8_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_8_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_8_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_8_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_8_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_8_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_8_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_8_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_8_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_8_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_8_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_8_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_8_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_8_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_8_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_8_io_uop_uopc),
    .io_uop_inst                    (_slots_8_io_uop_inst),
    .io_uop_debug_inst              (_slots_8_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_8_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_8_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_8_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_8_io_uop_fu_code),
    .io_uop_iw_state                (_slots_8_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_8_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_8_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_8_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_8_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_8_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_8_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_8_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_8_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_8_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_8_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_8_io_uop_pc_lob),
    .io_uop_taken                   (_slots_8_io_uop_taken),
    .io_uop_imm_packed              (_slots_8_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_8_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_8_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_8_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_8_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_8_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_8_io_uop_pdst),
    .io_uop_prs1                    (_slots_8_io_uop_prs1),
    .io_uop_prs2                    (_slots_8_io_uop_prs2),
    .io_uop_prs3                    (_slots_8_io_uop_prs3),
    .io_uop_ppred                   (_slots_8_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_8_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_8_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_8_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_8_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_8_io_uop_stale_pdst),
    .io_uop_exception               (_slots_8_io_uop_exception),
    .io_uop_exc_cause               (_slots_8_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_8_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_8_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_8_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_8_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_8_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_8_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_8_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_8_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_8_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_8_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_8_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_8_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_8_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_8_io_uop_ldst),
    .io_uop_lrs1                    (_slots_8_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_8_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_8_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_8_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_8_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_8_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_8_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_8_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_8_io_uop_fp_val),
    .io_uop_fp_single               (_slots_8_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_8_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_8_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_8_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_8_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_8_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_8_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_8_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_9 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_9_io_valid),
    .io_will_be_valid               (_slots_9_io_will_be_valid),
    .io_request                     (_slots_9_io_request),
    .io_grant                       (issue_slots_9_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_8),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_9_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_48 ? _slots_13_io_out_uop_uopc : _GEN_47 ? _slots_12_io_out_uop_uopc : _GEN_46 ? _slots_11_io_out_uop_uopc : _slots_10_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_48 ? _slots_13_io_out_uop_inst : _GEN_47 ? _slots_12_io_out_uop_inst : _GEN_46 ? _slots_11_io_out_uop_inst : _slots_10_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_48 ? _slots_13_io_out_uop_debug_inst : _GEN_47 ? _slots_12_io_out_uop_debug_inst : _GEN_46 ? _slots_11_io_out_uop_debug_inst : _slots_10_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_48 ? _slots_13_io_out_uop_is_rvc : _GEN_47 ? _slots_12_io_out_uop_is_rvc : _GEN_46 ? _slots_11_io_out_uop_is_rvc : _slots_10_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_48 ? _slots_13_io_out_uop_debug_pc : _GEN_47 ? _slots_12_io_out_uop_debug_pc : _GEN_46 ? _slots_11_io_out_uop_debug_pc : _slots_10_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_48 ? _slots_13_io_out_uop_iq_type : _GEN_47 ? _slots_12_io_out_uop_iq_type : _GEN_46 ? _slots_11_io_out_uop_iq_type : _slots_10_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_48 ? _slots_13_io_out_uop_fu_code : _GEN_47 ? _slots_12_io_out_uop_fu_code : _GEN_46 ? _slots_11_io_out_uop_fu_code : _slots_10_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_48 ? _slots_13_io_out_uop_iw_state : _GEN_47 ? _slots_12_io_out_uop_iw_state : _GEN_46 ? _slots_11_io_out_uop_iw_state : _slots_10_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_48 ? _slots_13_io_out_uop_iw_p1_poisoned : _GEN_47 ? _slots_12_io_out_uop_iw_p1_poisoned : _GEN_46 ? _slots_11_io_out_uop_iw_p1_poisoned : _slots_10_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_48 ? _slots_13_io_out_uop_iw_p2_poisoned : _GEN_47 ? _slots_12_io_out_uop_iw_p2_poisoned : _GEN_46 ? _slots_11_io_out_uop_iw_p2_poisoned : _slots_10_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_48 ? _slots_13_io_out_uop_is_br : _GEN_47 ? _slots_12_io_out_uop_is_br : _GEN_46 ? _slots_11_io_out_uop_is_br : _slots_10_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_48 ? _slots_13_io_out_uop_is_jalr : _GEN_47 ? _slots_12_io_out_uop_is_jalr : _GEN_46 ? _slots_11_io_out_uop_is_jalr : _slots_10_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_48 ? _slots_13_io_out_uop_is_jal : _GEN_47 ? _slots_12_io_out_uop_is_jal : _GEN_46 ? _slots_11_io_out_uop_is_jal : _slots_10_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_48 ? _slots_13_io_out_uop_is_sfb : _GEN_47 ? _slots_12_io_out_uop_is_sfb : _GEN_46 ? _slots_11_io_out_uop_is_sfb : _slots_10_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_48 ? _slots_13_io_out_uop_br_mask : _GEN_47 ? _slots_12_io_out_uop_br_mask : _GEN_46 ? _slots_11_io_out_uop_br_mask : _slots_10_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_48 ? _slots_13_io_out_uop_br_tag : _GEN_47 ? _slots_12_io_out_uop_br_tag : _GEN_46 ? _slots_11_io_out_uop_br_tag : _slots_10_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_48 ? _slots_13_io_out_uop_ftq_idx : _GEN_47 ? _slots_12_io_out_uop_ftq_idx : _GEN_46 ? _slots_11_io_out_uop_ftq_idx : _slots_10_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_48 ? _slots_13_io_out_uop_edge_inst : _GEN_47 ? _slots_12_io_out_uop_edge_inst : _GEN_46 ? _slots_11_io_out_uop_edge_inst : _slots_10_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_48 ? _slots_13_io_out_uop_pc_lob : _GEN_47 ? _slots_12_io_out_uop_pc_lob : _GEN_46 ? _slots_11_io_out_uop_pc_lob : _slots_10_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_48 ? _slots_13_io_out_uop_taken : _GEN_47 ? _slots_12_io_out_uop_taken : _GEN_46 ? _slots_11_io_out_uop_taken : _slots_10_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_48 ? _slots_13_io_out_uop_imm_packed : _GEN_47 ? _slots_12_io_out_uop_imm_packed : _GEN_46 ? _slots_11_io_out_uop_imm_packed : _slots_10_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_48 ? _slots_13_io_out_uop_csr_addr : _GEN_47 ? _slots_12_io_out_uop_csr_addr : _GEN_46 ? _slots_11_io_out_uop_csr_addr : _slots_10_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_48 ? _slots_13_io_out_uop_rob_idx : _GEN_47 ? _slots_12_io_out_uop_rob_idx : _GEN_46 ? _slots_11_io_out_uop_rob_idx : _slots_10_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_48 ? _slots_13_io_out_uop_ldq_idx : _GEN_47 ? _slots_12_io_out_uop_ldq_idx : _GEN_46 ? _slots_11_io_out_uop_ldq_idx : _slots_10_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_48 ? _slots_13_io_out_uop_stq_idx : _GEN_47 ? _slots_12_io_out_uop_stq_idx : _GEN_46 ? _slots_11_io_out_uop_stq_idx : _slots_10_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_48 ? _slots_13_io_out_uop_rxq_idx : _GEN_47 ? _slots_12_io_out_uop_rxq_idx : _GEN_46 ? _slots_11_io_out_uop_rxq_idx : _slots_10_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_48 ? _slots_13_io_out_uop_pdst : _GEN_47 ? _slots_12_io_out_uop_pdst : _GEN_46 ? _slots_11_io_out_uop_pdst : _slots_10_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_48 ? _slots_13_io_out_uop_prs1 : _GEN_47 ? _slots_12_io_out_uop_prs1 : _GEN_46 ? _slots_11_io_out_uop_prs1 : _slots_10_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_48 ? _slots_13_io_out_uop_prs2 : _GEN_47 ? _slots_12_io_out_uop_prs2 : _GEN_46 ? _slots_11_io_out_uop_prs2 : _slots_10_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_48 ? _slots_13_io_out_uop_prs3 : _GEN_47 ? _slots_12_io_out_uop_prs3 : _GEN_46 ? _slots_11_io_out_uop_prs3 : _slots_10_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_48 ? _slots_13_io_out_uop_ppred : _GEN_47 ? _slots_12_io_out_uop_ppred : _GEN_46 ? _slots_11_io_out_uop_ppred : _slots_10_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_48 ? _slots_13_io_out_uop_prs1_busy : _GEN_47 ? _slots_12_io_out_uop_prs1_busy : _GEN_46 ? _slots_11_io_out_uop_prs1_busy : _slots_10_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_48 ? _slots_13_io_out_uop_prs2_busy : _GEN_47 ? _slots_12_io_out_uop_prs2_busy : _GEN_46 ? _slots_11_io_out_uop_prs2_busy : _slots_10_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_48 ? _slots_13_io_out_uop_prs3_busy : _GEN_47 ? _slots_12_io_out_uop_prs3_busy : _GEN_46 ? _slots_11_io_out_uop_prs3_busy : _slots_10_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_48 ? _slots_13_io_out_uop_ppred_busy : _GEN_47 ? _slots_12_io_out_uop_ppred_busy : _GEN_46 ? _slots_11_io_out_uop_ppred_busy : _slots_10_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_48 ? _slots_13_io_out_uop_stale_pdst : _GEN_47 ? _slots_12_io_out_uop_stale_pdst : _GEN_46 ? _slots_11_io_out_uop_stale_pdst : _slots_10_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_48 ? _slots_13_io_out_uop_exception : _GEN_47 ? _slots_12_io_out_uop_exception : _GEN_46 ? _slots_11_io_out_uop_exception : _slots_10_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_48 ? _slots_13_io_out_uop_exc_cause : _GEN_47 ? _slots_12_io_out_uop_exc_cause : _GEN_46 ? _slots_11_io_out_uop_exc_cause : _slots_10_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_48 ? _slots_13_io_out_uop_bypassable : _GEN_47 ? _slots_12_io_out_uop_bypassable : _GEN_46 ? _slots_11_io_out_uop_bypassable : _slots_10_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_48 ? _slots_13_io_out_uop_mem_cmd : _GEN_47 ? _slots_12_io_out_uop_mem_cmd : _GEN_46 ? _slots_11_io_out_uop_mem_cmd : _slots_10_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_48 ? _slots_13_io_out_uop_mem_size : _GEN_47 ? _slots_12_io_out_uop_mem_size : _GEN_46 ? _slots_11_io_out_uop_mem_size : _slots_10_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_48 ? _slots_13_io_out_uop_mem_signed : _GEN_47 ? _slots_12_io_out_uop_mem_signed : _GEN_46 ? _slots_11_io_out_uop_mem_signed : _slots_10_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_48 ? _slots_13_io_out_uop_is_fence : _GEN_47 ? _slots_12_io_out_uop_is_fence : _GEN_46 ? _slots_11_io_out_uop_is_fence : _slots_10_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_48 ? _slots_13_io_out_uop_is_fencei : _GEN_47 ? _slots_12_io_out_uop_is_fencei : _GEN_46 ? _slots_11_io_out_uop_is_fencei : _slots_10_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_48 ? _slots_13_io_out_uop_is_amo : _GEN_47 ? _slots_12_io_out_uop_is_amo : _GEN_46 ? _slots_11_io_out_uop_is_amo : _slots_10_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_48 ? _slots_13_io_out_uop_uses_ldq : _GEN_47 ? _slots_12_io_out_uop_uses_ldq : _GEN_46 ? _slots_11_io_out_uop_uses_ldq : _slots_10_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_48 ? _slots_13_io_out_uop_uses_stq : _GEN_47 ? _slots_12_io_out_uop_uses_stq : _GEN_46 ? _slots_11_io_out_uop_uses_stq : _slots_10_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_48 ? _slots_13_io_out_uop_is_sys_pc2epc : _GEN_47 ? _slots_12_io_out_uop_is_sys_pc2epc : _GEN_46 ? _slots_11_io_out_uop_is_sys_pc2epc : _slots_10_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_48 ? _slots_13_io_out_uop_is_unique : _GEN_47 ? _slots_12_io_out_uop_is_unique : _GEN_46 ? _slots_11_io_out_uop_is_unique : _slots_10_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_48 ? _slots_13_io_out_uop_flush_on_commit : _GEN_47 ? _slots_12_io_out_uop_flush_on_commit : _GEN_46 ? _slots_11_io_out_uop_flush_on_commit : _slots_10_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_48 ? _slots_13_io_out_uop_ldst_is_rs1 : _GEN_47 ? _slots_12_io_out_uop_ldst_is_rs1 : _GEN_46 ? _slots_11_io_out_uop_ldst_is_rs1 : _slots_10_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_48 ? _slots_13_io_out_uop_ldst : _GEN_47 ? _slots_12_io_out_uop_ldst : _GEN_46 ? _slots_11_io_out_uop_ldst : _slots_10_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_48 ? _slots_13_io_out_uop_lrs1 : _GEN_47 ? _slots_12_io_out_uop_lrs1 : _GEN_46 ? _slots_11_io_out_uop_lrs1 : _slots_10_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_48 ? _slots_13_io_out_uop_lrs2 : _GEN_47 ? _slots_12_io_out_uop_lrs2 : _GEN_46 ? _slots_11_io_out_uop_lrs2 : _slots_10_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_48 ? _slots_13_io_out_uop_lrs3 : _GEN_47 ? _slots_12_io_out_uop_lrs3 : _GEN_46 ? _slots_11_io_out_uop_lrs3 : _slots_10_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_48 ? _slots_13_io_out_uop_ldst_val : _GEN_47 ? _slots_12_io_out_uop_ldst_val : _GEN_46 ? _slots_11_io_out_uop_ldst_val : _slots_10_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_48 ? _slots_13_io_out_uop_dst_rtype : _GEN_47 ? _slots_12_io_out_uop_dst_rtype : _GEN_46 ? _slots_11_io_out_uop_dst_rtype : _slots_10_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_48 ? _slots_13_io_out_uop_lrs1_rtype : _GEN_47 ? _slots_12_io_out_uop_lrs1_rtype : _GEN_46 ? _slots_11_io_out_uop_lrs1_rtype : _slots_10_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_48 ? _slots_13_io_out_uop_lrs2_rtype : _GEN_47 ? _slots_12_io_out_uop_lrs2_rtype : _GEN_46 ? _slots_11_io_out_uop_lrs2_rtype : _slots_10_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_48 ? _slots_13_io_out_uop_frs3_en : _GEN_47 ? _slots_12_io_out_uop_frs3_en : _GEN_46 ? _slots_11_io_out_uop_frs3_en : _slots_10_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_48 ? _slots_13_io_out_uop_fp_val : _GEN_47 ? _slots_12_io_out_uop_fp_val : _GEN_46 ? _slots_11_io_out_uop_fp_val : _slots_10_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_48 ? _slots_13_io_out_uop_fp_single : _GEN_47 ? _slots_12_io_out_uop_fp_single : _GEN_46 ? _slots_11_io_out_uop_fp_single : _slots_10_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_48 ? _slots_13_io_out_uop_xcpt_pf_if : _GEN_47 ? _slots_12_io_out_uop_xcpt_pf_if : _GEN_46 ? _slots_11_io_out_uop_xcpt_pf_if : _slots_10_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_48 ? _slots_13_io_out_uop_xcpt_ae_if : _GEN_47 ? _slots_12_io_out_uop_xcpt_ae_if : _GEN_46 ? _slots_11_io_out_uop_xcpt_ae_if : _slots_10_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_48 ? _slots_13_io_out_uop_xcpt_ma_if : _GEN_47 ? _slots_12_io_out_uop_xcpt_ma_if : _GEN_46 ? _slots_11_io_out_uop_xcpt_ma_if : _slots_10_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_48 ? _slots_13_io_out_uop_bp_debug_if : _GEN_47 ? _slots_12_io_out_uop_bp_debug_if : _GEN_46 ? _slots_11_io_out_uop_bp_debug_if : _slots_10_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_48 ? _slots_13_io_out_uop_bp_xcpt_if : _GEN_47 ? _slots_12_io_out_uop_bp_xcpt_if : _GEN_46 ? _slots_11_io_out_uop_bp_xcpt_if : _slots_10_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_48 ? _slots_13_io_out_uop_debug_fsrc : _GEN_47 ? _slots_12_io_out_uop_debug_fsrc : _GEN_46 ? _slots_11_io_out_uop_debug_fsrc : _slots_10_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_48 ? _slots_13_io_out_uop_debug_tsrc : _GEN_47 ? _slots_12_io_out_uop_debug_tsrc : _GEN_46 ? _slots_11_io_out_uop_debug_tsrc : _slots_10_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_9_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_9_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_9_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_9_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_9_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_9_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_9_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_9_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_9_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_9_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_9_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_9_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_9_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_9_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_9_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_9_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_9_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_9_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_9_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_9_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_9_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_9_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_9_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_9_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_9_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_9_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_9_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_9_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_9_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_9_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_9_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_9_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_9_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_9_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_9_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_9_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_9_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_9_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_9_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_9_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_9_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_9_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_9_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_9_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_9_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_9_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_9_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_9_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_9_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_9_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_9_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_9_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_9_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_9_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_9_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_9_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_9_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_9_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_9_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_9_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_9_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_9_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_9_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_9_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_9_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_9_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_9_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_9_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_9_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_9_io_uop_uopc),
    .io_uop_inst                    (_slots_9_io_uop_inst),
    .io_uop_debug_inst              (_slots_9_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_9_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_9_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_9_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_9_io_uop_fu_code),
    .io_uop_iw_state                (_slots_9_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_9_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_9_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_9_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_9_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_9_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_9_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_9_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_9_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_9_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_9_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_9_io_uop_pc_lob),
    .io_uop_taken                   (_slots_9_io_uop_taken),
    .io_uop_imm_packed              (_slots_9_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_9_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_9_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_9_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_9_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_9_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_9_io_uop_pdst),
    .io_uop_prs1                    (_slots_9_io_uop_prs1),
    .io_uop_prs2                    (_slots_9_io_uop_prs2),
    .io_uop_prs3                    (_slots_9_io_uop_prs3),
    .io_uop_ppred                   (_slots_9_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_9_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_9_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_9_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_9_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_9_io_uop_stale_pdst),
    .io_uop_exception               (_slots_9_io_uop_exception),
    .io_uop_exc_cause               (_slots_9_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_9_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_9_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_9_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_9_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_9_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_9_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_9_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_9_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_9_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_9_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_9_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_9_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_9_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_9_io_uop_ldst),
    .io_uop_lrs1                    (_slots_9_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_9_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_9_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_9_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_9_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_9_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_9_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_9_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_9_io_uop_fp_val),
    .io_uop_fp_single               (_slots_9_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_9_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_9_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_9_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_9_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_9_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_9_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_9_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_10 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_10_io_valid),
    .io_will_be_valid               (_slots_10_io_will_be_valid),
    .io_request                     (_slots_10_io_request),
    .io_grant                       (issue_slots_10_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_9),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_10_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_51 ? _slots_14_io_out_uop_uopc : _GEN_50 ? _slots_13_io_out_uop_uopc : _GEN_49 ? _slots_12_io_out_uop_uopc : _slots_11_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_51 ? _slots_14_io_out_uop_inst : _GEN_50 ? _slots_13_io_out_uop_inst : _GEN_49 ? _slots_12_io_out_uop_inst : _slots_11_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_51 ? _slots_14_io_out_uop_debug_inst : _GEN_50 ? _slots_13_io_out_uop_debug_inst : _GEN_49 ? _slots_12_io_out_uop_debug_inst : _slots_11_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_51 ? _slots_14_io_out_uop_is_rvc : _GEN_50 ? _slots_13_io_out_uop_is_rvc : _GEN_49 ? _slots_12_io_out_uop_is_rvc : _slots_11_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_51 ? _slots_14_io_out_uop_debug_pc : _GEN_50 ? _slots_13_io_out_uop_debug_pc : _GEN_49 ? _slots_12_io_out_uop_debug_pc : _slots_11_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_51 ? _slots_14_io_out_uop_iq_type : _GEN_50 ? _slots_13_io_out_uop_iq_type : _GEN_49 ? _slots_12_io_out_uop_iq_type : _slots_11_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_51 ? _slots_14_io_out_uop_fu_code : _GEN_50 ? _slots_13_io_out_uop_fu_code : _GEN_49 ? _slots_12_io_out_uop_fu_code : _slots_11_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_51 ? _slots_14_io_out_uop_iw_state : _GEN_50 ? _slots_13_io_out_uop_iw_state : _GEN_49 ? _slots_12_io_out_uop_iw_state : _slots_11_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_51 ? _slots_14_io_out_uop_iw_p1_poisoned : _GEN_50 ? _slots_13_io_out_uop_iw_p1_poisoned : _GEN_49 ? _slots_12_io_out_uop_iw_p1_poisoned : _slots_11_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_51 ? _slots_14_io_out_uop_iw_p2_poisoned : _GEN_50 ? _slots_13_io_out_uop_iw_p2_poisoned : _GEN_49 ? _slots_12_io_out_uop_iw_p2_poisoned : _slots_11_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_51 ? _slots_14_io_out_uop_is_br : _GEN_50 ? _slots_13_io_out_uop_is_br : _GEN_49 ? _slots_12_io_out_uop_is_br : _slots_11_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_51 ? _slots_14_io_out_uop_is_jalr : _GEN_50 ? _slots_13_io_out_uop_is_jalr : _GEN_49 ? _slots_12_io_out_uop_is_jalr : _slots_11_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_51 ? _slots_14_io_out_uop_is_jal : _GEN_50 ? _slots_13_io_out_uop_is_jal : _GEN_49 ? _slots_12_io_out_uop_is_jal : _slots_11_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_51 ? _slots_14_io_out_uop_is_sfb : _GEN_50 ? _slots_13_io_out_uop_is_sfb : _GEN_49 ? _slots_12_io_out_uop_is_sfb : _slots_11_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_51 ? _slots_14_io_out_uop_br_mask : _GEN_50 ? _slots_13_io_out_uop_br_mask : _GEN_49 ? _slots_12_io_out_uop_br_mask : _slots_11_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_51 ? _slots_14_io_out_uop_br_tag : _GEN_50 ? _slots_13_io_out_uop_br_tag : _GEN_49 ? _slots_12_io_out_uop_br_tag : _slots_11_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_51 ? _slots_14_io_out_uop_ftq_idx : _GEN_50 ? _slots_13_io_out_uop_ftq_idx : _GEN_49 ? _slots_12_io_out_uop_ftq_idx : _slots_11_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_51 ? _slots_14_io_out_uop_edge_inst : _GEN_50 ? _slots_13_io_out_uop_edge_inst : _GEN_49 ? _slots_12_io_out_uop_edge_inst : _slots_11_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_51 ? _slots_14_io_out_uop_pc_lob : _GEN_50 ? _slots_13_io_out_uop_pc_lob : _GEN_49 ? _slots_12_io_out_uop_pc_lob : _slots_11_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_51 ? _slots_14_io_out_uop_taken : _GEN_50 ? _slots_13_io_out_uop_taken : _GEN_49 ? _slots_12_io_out_uop_taken : _slots_11_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_51 ? _slots_14_io_out_uop_imm_packed : _GEN_50 ? _slots_13_io_out_uop_imm_packed : _GEN_49 ? _slots_12_io_out_uop_imm_packed : _slots_11_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_51 ? _slots_14_io_out_uop_csr_addr : _GEN_50 ? _slots_13_io_out_uop_csr_addr : _GEN_49 ? _slots_12_io_out_uop_csr_addr : _slots_11_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_51 ? _slots_14_io_out_uop_rob_idx : _GEN_50 ? _slots_13_io_out_uop_rob_idx : _GEN_49 ? _slots_12_io_out_uop_rob_idx : _slots_11_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_51 ? _slots_14_io_out_uop_ldq_idx : _GEN_50 ? _slots_13_io_out_uop_ldq_idx : _GEN_49 ? _slots_12_io_out_uop_ldq_idx : _slots_11_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_51 ? _slots_14_io_out_uop_stq_idx : _GEN_50 ? _slots_13_io_out_uop_stq_idx : _GEN_49 ? _slots_12_io_out_uop_stq_idx : _slots_11_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_51 ? _slots_14_io_out_uop_rxq_idx : _GEN_50 ? _slots_13_io_out_uop_rxq_idx : _GEN_49 ? _slots_12_io_out_uop_rxq_idx : _slots_11_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_51 ? _slots_14_io_out_uop_pdst : _GEN_50 ? _slots_13_io_out_uop_pdst : _GEN_49 ? _slots_12_io_out_uop_pdst : _slots_11_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_51 ? _slots_14_io_out_uop_prs1 : _GEN_50 ? _slots_13_io_out_uop_prs1 : _GEN_49 ? _slots_12_io_out_uop_prs1 : _slots_11_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_51 ? _slots_14_io_out_uop_prs2 : _GEN_50 ? _slots_13_io_out_uop_prs2 : _GEN_49 ? _slots_12_io_out_uop_prs2 : _slots_11_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_51 ? _slots_14_io_out_uop_prs3 : _GEN_50 ? _slots_13_io_out_uop_prs3 : _GEN_49 ? _slots_12_io_out_uop_prs3 : _slots_11_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_51 ? _slots_14_io_out_uop_ppred : _GEN_50 ? _slots_13_io_out_uop_ppred : _GEN_49 ? _slots_12_io_out_uop_ppred : _slots_11_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_51 ? _slots_14_io_out_uop_prs1_busy : _GEN_50 ? _slots_13_io_out_uop_prs1_busy : _GEN_49 ? _slots_12_io_out_uop_prs1_busy : _slots_11_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_51 ? _slots_14_io_out_uop_prs2_busy : _GEN_50 ? _slots_13_io_out_uop_prs2_busy : _GEN_49 ? _slots_12_io_out_uop_prs2_busy : _slots_11_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_51 ? _slots_14_io_out_uop_prs3_busy : _GEN_50 ? _slots_13_io_out_uop_prs3_busy : _GEN_49 ? _slots_12_io_out_uop_prs3_busy : _slots_11_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_51 ? _slots_14_io_out_uop_ppred_busy : _GEN_50 ? _slots_13_io_out_uop_ppred_busy : _GEN_49 ? _slots_12_io_out_uop_ppred_busy : _slots_11_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_51 ? _slots_14_io_out_uop_stale_pdst : _GEN_50 ? _slots_13_io_out_uop_stale_pdst : _GEN_49 ? _slots_12_io_out_uop_stale_pdst : _slots_11_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_51 ? _slots_14_io_out_uop_exception : _GEN_50 ? _slots_13_io_out_uop_exception : _GEN_49 ? _slots_12_io_out_uop_exception : _slots_11_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_51 ? _slots_14_io_out_uop_exc_cause : _GEN_50 ? _slots_13_io_out_uop_exc_cause : _GEN_49 ? _slots_12_io_out_uop_exc_cause : _slots_11_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_51 ? _slots_14_io_out_uop_bypassable : _GEN_50 ? _slots_13_io_out_uop_bypassable : _GEN_49 ? _slots_12_io_out_uop_bypassable : _slots_11_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_51 ? _slots_14_io_out_uop_mem_cmd : _GEN_50 ? _slots_13_io_out_uop_mem_cmd : _GEN_49 ? _slots_12_io_out_uop_mem_cmd : _slots_11_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_51 ? _slots_14_io_out_uop_mem_size : _GEN_50 ? _slots_13_io_out_uop_mem_size : _GEN_49 ? _slots_12_io_out_uop_mem_size : _slots_11_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_51 ? _slots_14_io_out_uop_mem_signed : _GEN_50 ? _slots_13_io_out_uop_mem_signed : _GEN_49 ? _slots_12_io_out_uop_mem_signed : _slots_11_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_51 ? _slots_14_io_out_uop_is_fence : _GEN_50 ? _slots_13_io_out_uop_is_fence : _GEN_49 ? _slots_12_io_out_uop_is_fence : _slots_11_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_51 ? _slots_14_io_out_uop_is_fencei : _GEN_50 ? _slots_13_io_out_uop_is_fencei : _GEN_49 ? _slots_12_io_out_uop_is_fencei : _slots_11_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_51 ? _slots_14_io_out_uop_is_amo : _GEN_50 ? _slots_13_io_out_uop_is_amo : _GEN_49 ? _slots_12_io_out_uop_is_amo : _slots_11_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_51 ? _slots_14_io_out_uop_uses_ldq : _GEN_50 ? _slots_13_io_out_uop_uses_ldq : _GEN_49 ? _slots_12_io_out_uop_uses_ldq : _slots_11_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_51 ? _slots_14_io_out_uop_uses_stq : _GEN_50 ? _slots_13_io_out_uop_uses_stq : _GEN_49 ? _slots_12_io_out_uop_uses_stq : _slots_11_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_51 ? _slots_14_io_out_uop_is_sys_pc2epc : _GEN_50 ? _slots_13_io_out_uop_is_sys_pc2epc : _GEN_49 ? _slots_12_io_out_uop_is_sys_pc2epc : _slots_11_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_51 ? _slots_14_io_out_uop_is_unique : _GEN_50 ? _slots_13_io_out_uop_is_unique : _GEN_49 ? _slots_12_io_out_uop_is_unique : _slots_11_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_51 ? _slots_14_io_out_uop_flush_on_commit : _GEN_50 ? _slots_13_io_out_uop_flush_on_commit : _GEN_49 ? _slots_12_io_out_uop_flush_on_commit : _slots_11_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_51 ? _slots_14_io_out_uop_ldst_is_rs1 : _GEN_50 ? _slots_13_io_out_uop_ldst_is_rs1 : _GEN_49 ? _slots_12_io_out_uop_ldst_is_rs1 : _slots_11_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_51 ? _slots_14_io_out_uop_ldst : _GEN_50 ? _slots_13_io_out_uop_ldst : _GEN_49 ? _slots_12_io_out_uop_ldst : _slots_11_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_51 ? _slots_14_io_out_uop_lrs1 : _GEN_50 ? _slots_13_io_out_uop_lrs1 : _GEN_49 ? _slots_12_io_out_uop_lrs1 : _slots_11_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_51 ? _slots_14_io_out_uop_lrs2 : _GEN_50 ? _slots_13_io_out_uop_lrs2 : _GEN_49 ? _slots_12_io_out_uop_lrs2 : _slots_11_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_51 ? _slots_14_io_out_uop_lrs3 : _GEN_50 ? _slots_13_io_out_uop_lrs3 : _GEN_49 ? _slots_12_io_out_uop_lrs3 : _slots_11_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_51 ? _slots_14_io_out_uop_ldst_val : _GEN_50 ? _slots_13_io_out_uop_ldst_val : _GEN_49 ? _slots_12_io_out_uop_ldst_val : _slots_11_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_51 ? _slots_14_io_out_uop_dst_rtype : _GEN_50 ? _slots_13_io_out_uop_dst_rtype : _GEN_49 ? _slots_12_io_out_uop_dst_rtype : _slots_11_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_51 ? _slots_14_io_out_uop_lrs1_rtype : _GEN_50 ? _slots_13_io_out_uop_lrs1_rtype : _GEN_49 ? _slots_12_io_out_uop_lrs1_rtype : _slots_11_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_51 ? _slots_14_io_out_uop_lrs2_rtype : _GEN_50 ? _slots_13_io_out_uop_lrs2_rtype : _GEN_49 ? _slots_12_io_out_uop_lrs2_rtype : _slots_11_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_51 ? _slots_14_io_out_uop_frs3_en : _GEN_50 ? _slots_13_io_out_uop_frs3_en : _GEN_49 ? _slots_12_io_out_uop_frs3_en : _slots_11_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_51 ? _slots_14_io_out_uop_fp_val : _GEN_50 ? _slots_13_io_out_uop_fp_val : _GEN_49 ? _slots_12_io_out_uop_fp_val : _slots_11_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_51 ? _slots_14_io_out_uop_fp_single : _GEN_50 ? _slots_13_io_out_uop_fp_single : _GEN_49 ? _slots_12_io_out_uop_fp_single : _slots_11_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_51 ? _slots_14_io_out_uop_xcpt_pf_if : _GEN_50 ? _slots_13_io_out_uop_xcpt_pf_if : _GEN_49 ? _slots_12_io_out_uop_xcpt_pf_if : _slots_11_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_51 ? _slots_14_io_out_uop_xcpt_ae_if : _GEN_50 ? _slots_13_io_out_uop_xcpt_ae_if : _GEN_49 ? _slots_12_io_out_uop_xcpt_ae_if : _slots_11_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_51 ? _slots_14_io_out_uop_xcpt_ma_if : _GEN_50 ? _slots_13_io_out_uop_xcpt_ma_if : _GEN_49 ? _slots_12_io_out_uop_xcpt_ma_if : _slots_11_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_51 ? _slots_14_io_out_uop_bp_debug_if : _GEN_50 ? _slots_13_io_out_uop_bp_debug_if : _GEN_49 ? _slots_12_io_out_uop_bp_debug_if : _slots_11_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_51 ? _slots_14_io_out_uop_bp_xcpt_if : _GEN_50 ? _slots_13_io_out_uop_bp_xcpt_if : _GEN_49 ? _slots_12_io_out_uop_bp_xcpt_if : _slots_11_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_51 ? _slots_14_io_out_uop_debug_fsrc : _GEN_50 ? _slots_13_io_out_uop_debug_fsrc : _GEN_49 ? _slots_12_io_out_uop_debug_fsrc : _slots_11_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_51 ? _slots_14_io_out_uop_debug_tsrc : _GEN_50 ? _slots_13_io_out_uop_debug_tsrc : _GEN_49 ? _slots_12_io_out_uop_debug_tsrc : _slots_11_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_10_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_10_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_10_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_10_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_10_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_10_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_10_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_10_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_10_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_10_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_10_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_10_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_10_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_10_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_10_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_10_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_10_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_10_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_10_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_10_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_10_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_10_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_10_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_10_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_10_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_10_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_10_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_10_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_10_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_10_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_10_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_10_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_10_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_10_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_10_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_10_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_10_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_10_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_10_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_10_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_10_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_10_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_10_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_10_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_10_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_10_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_10_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_10_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_10_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_10_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_10_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_10_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_10_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_10_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_10_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_10_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_10_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_10_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_10_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_10_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_10_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_10_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_10_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_10_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_10_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_10_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_10_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_10_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_10_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_10_io_uop_uopc),
    .io_uop_inst                    (_slots_10_io_uop_inst),
    .io_uop_debug_inst              (_slots_10_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_10_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_10_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_10_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_10_io_uop_fu_code),
    .io_uop_iw_state                (_slots_10_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_10_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_10_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_10_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_10_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_10_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_10_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_10_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_10_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_10_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_10_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_10_io_uop_pc_lob),
    .io_uop_taken                   (_slots_10_io_uop_taken),
    .io_uop_imm_packed              (_slots_10_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_10_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_10_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_10_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_10_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_10_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_10_io_uop_pdst),
    .io_uop_prs1                    (_slots_10_io_uop_prs1),
    .io_uop_prs2                    (_slots_10_io_uop_prs2),
    .io_uop_prs3                    (_slots_10_io_uop_prs3),
    .io_uop_ppred                   (_slots_10_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_10_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_10_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_10_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_10_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_10_io_uop_stale_pdst),
    .io_uop_exception               (_slots_10_io_uop_exception),
    .io_uop_exc_cause               (_slots_10_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_10_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_10_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_10_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_10_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_10_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_10_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_10_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_10_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_10_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_10_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_10_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_10_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_10_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_10_io_uop_ldst),
    .io_uop_lrs1                    (_slots_10_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_10_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_10_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_10_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_10_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_10_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_10_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_10_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_10_io_uop_fp_val),
    .io_uop_fp_single               (_slots_10_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_10_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_10_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_10_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_10_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_10_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_10_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_10_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_11 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_11_io_valid),
    .io_will_be_valid               (_slots_11_io_will_be_valid),
    .io_request                     (_slots_11_io_request),
    .io_grant                       (issue_slots_11_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_10),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_11_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_54 ? _slots_15_io_out_uop_uopc : _GEN_53 ? _slots_14_io_out_uop_uopc : _GEN_52 ? _slots_13_io_out_uop_uopc : _slots_12_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_54 ? _slots_15_io_out_uop_inst : _GEN_53 ? _slots_14_io_out_uop_inst : _GEN_52 ? _slots_13_io_out_uop_inst : _slots_12_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_54 ? _slots_15_io_out_uop_debug_inst : _GEN_53 ? _slots_14_io_out_uop_debug_inst : _GEN_52 ? _slots_13_io_out_uop_debug_inst : _slots_12_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_54 ? _slots_15_io_out_uop_is_rvc : _GEN_53 ? _slots_14_io_out_uop_is_rvc : _GEN_52 ? _slots_13_io_out_uop_is_rvc : _slots_12_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_54 ? _slots_15_io_out_uop_debug_pc : _GEN_53 ? _slots_14_io_out_uop_debug_pc : _GEN_52 ? _slots_13_io_out_uop_debug_pc : _slots_12_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_54 ? _slots_15_io_out_uop_iq_type : _GEN_53 ? _slots_14_io_out_uop_iq_type : _GEN_52 ? _slots_13_io_out_uop_iq_type : _slots_12_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_54 ? _slots_15_io_out_uop_fu_code : _GEN_53 ? _slots_14_io_out_uop_fu_code : _GEN_52 ? _slots_13_io_out_uop_fu_code : _slots_12_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_54 ? _slots_15_io_out_uop_iw_state : _GEN_53 ? _slots_14_io_out_uop_iw_state : _GEN_52 ? _slots_13_io_out_uop_iw_state : _slots_12_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_54 ? _slots_15_io_out_uop_iw_p1_poisoned : _GEN_53 ? _slots_14_io_out_uop_iw_p1_poisoned : _GEN_52 ? _slots_13_io_out_uop_iw_p1_poisoned : _slots_12_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_54 ? _slots_15_io_out_uop_iw_p2_poisoned : _GEN_53 ? _slots_14_io_out_uop_iw_p2_poisoned : _GEN_52 ? _slots_13_io_out_uop_iw_p2_poisoned : _slots_12_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_54 ? _slots_15_io_out_uop_is_br : _GEN_53 ? _slots_14_io_out_uop_is_br : _GEN_52 ? _slots_13_io_out_uop_is_br : _slots_12_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_54 ? _slots_15_io_out_uop_is_jalr : _GEN_53 ? _slots_14_io_out_uop_is_jalr : _GEN_52 ? _slots_13_io_out_uop_is_jalr : _slots_12_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_54 ? _slots_15_io_out_uop_is_jal : _GEN_53 ? _slots_14_io_out_uop_is_jal : _GEN_52 ? _slots_13_io_out_uop_is_jal : _slots_12_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_54 ? _slots_15_io_out_uop_is_sfb : _GEN_53 ? _slots_14_io_out_uop_is_sfb : _GEN_52 ? _slots_13_io_out_uop_is_sfb : _slots_12_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_54 ? _slots_15_io_out_uop_br_mask : _GEN_53 ? _slots_14_io_out_uop_br_mask : _GEN_52 ? _slots_13_io_out_uop_br_mask : _slots_12_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_54 ? _slots_15_io_out_uop_br_tag : _GEN_53 ? _slots_14_io_out_uop_br_tag : _GEN_52 ? _slots_13_io_out_uop_br_tag : _slots_12_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_54 ? _slots_15_io_out_uop_ftq_idx : _GEN_53 ? _slots_14_io_out_uop_ftq_idx : _GEN_52 ? _slots_13_io_out_uop_ftq_idx : _slots_12_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_54 ? _slots_15_io_out_uop_edge_inst : _GEN_53 ? _slots_14_io_out_uop_edge_inst : _GEN_52 ? _slots_13_io_out_uop_edge_inst : _slots_12_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_54 ? _slots_15_io_out_uop_pc_lob : _GEN_53 ? _slots_14_io_out_uop_pc_lob : _GEN_52 ? _slots_13_io_out_uop_pc_lob : _slots_12_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_54 ? _slots_15_io_out_uop_taken : _GEN_53 ? _slots_14_io_out_uop_taken : _GEN_52 ? _slots_13_io_out_uop_taken : _slots_12_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_54 ? _slots_15_io_out_uop_imm_packed : _GEN_53 ? _slots_14_io_out_uop_imm_packed : _GEN_52 ? _slots_13_io_out_uop_imm_packed : _slots_12_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_54 ? _slots_15_io_out_uop_csr_addr : _GEN_53 ? _slots_14_io_out_uop_csr_addr : _GEN_52 ? _slots_13_io_out_uop_csr_addr : _slots_12_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_54 ? _slots_15_io_out_uop_rob_idx : _GEN_53 ? _slots_14_io_out_uop_rob_idx : _GEN_52 ? _slots_13_io_out_uop_rob_idx : _slots_12_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_54 ? _slots_15_io_out_uop_ldq_idx : _GEN_53 ? _slots_14_io_out_uop_ldq_idx : _GEN_52 ? _slots_13_io_out_uop_ldq_idx : _slots_12_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_54 ? _slots_15_io_out_uop_stq_idx : _GEN_53 ? _slots_14_io_out_uop_stq_idx : _GEN_52 ? _slots_13_io_out_uop_stq_idx : _slots_12_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_54 ? _slots_15_io_out_uop_rxq_idx : _GEN_53 ? _slots_14_io_out_uop_rxq_idx : _GEN_52 ? _slots_13_io_out_uop_rxq_idx : _slots_12_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_54 ? _slots_15_io_out_uop_pdst : _GEN_53 ? _slots_14_io_out_uop_pdst : _GEN_52 ? _slots_13_io_out_uop_pdst : _slots_12_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_54 ? _slots_15_io_out_uop_prs1 : _GEN_53 ? _slots_14_io_out_uop_prs1 : _GEN_52 ? _slots_13_io_out_uop_prs1 : _slots_12_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_54 ? _slots_15_io_out_uop_prs2 : _GEN_53 ? _slots_14_io_out_uop_prs2 : _GEN_52 ? _slots_13_io_out_uop_prs2 : _slots_12_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_54 ? _slots_15_io_out_uop_prs3 : _GEN_53 ? _slots_14_io_out_uop_prs3 : _GEN_52 ? _slots_13_io_out_uop_prs3 : _slots_12_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_54 ? _slots_15_io_out_uop_ppred : _GEN_53 ? _slots_14_io_out_uop_ppred : _GEN_52 ? _slots_13_io_out_uop_ppred : _slots_12_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_54 ? _slots_15_io_out_uop_prs1_busy : _GEN_53 ? _slots_14_io_out_uop_prs1_busy : _GEN_52 ? _slots_13_io_out_uop_prs1_busy : _slots_12_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_54 ? _slots_15_io_out_uop_prs2_busy : _GEN_53 ? _slots_14_io_out_uop_prs2_busy : _GEN_52 ? _slots_13_io_out_uop_prs2_busy : _slots_12_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_54 ? _slots_15_io_out_uop_prs3_busy : _GEN_53 ? _slots_14_io_out_uop_prs3_busy : _GEN_52 ? _slots_13_io_out_uop_prs3_busy : _slots_12_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_54 ? _slots_15_io_out_uop_ppred_busy : _GEN_53 ? _slots_14_io_out_uop_ppred_busy : _GEN_52 ? _slots_13_io_out_uop_ppred_busy : _slots_12_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_54 ? _slots_15_io_out_uop_stale_pdst : _GEN_53 ? _slots_14_io_out_uop_stale_pdst : _GEN_52 ? _slots_13_io_out_uop_stale_pdst : _slots_12_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_54 ? _slots_15_io_out_uop_exception : _GEN_53 ? _slots_14_io_out_uop_exception : _GEN_52 ? _slots_13_io_out_uop_exception : _slots_12_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_54 ? _slots_15_io_out_uop_exc_cause : _GEN_53 ? _slots_14_io_out_uop_exc_cause : _GEN_52 ? _slots_13_io_out_uop_exc_cause : _slots_12_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_54 ? _slots_15_io_out_uop_bypassable : _GEN_53 ? _slots_14_io_out_uop_bypassable : _GEN_52 ? _slots_13_io_out_uop_bypassable : _slots_12_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_54 ? _slots_15_io_out_uop_mem_cmd : _GEN_53 ? _slots_14_io_out_uop_mem_cmd : _GEN_52 ? _slots_13_io_out_uop_mem_cmd : _slots_12_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_54 ? _slots_15_io_out_uop_mem_size : _GEN_53 ? _slots_14_io_out_uop_mem_size : _GEN_52 ? _slots_13_io_out_uop_mem_size : _slots_12_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_54 ? _slots_15_io_out_uop_mem_signed : _GEN_53 ? _slots_14_io_out_uop_mem_signed : _GEN_52 ? _slots_13_io_out_uop_mem_signed : _slots_12_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_54 ? _slots_15_io_out_uop_is_fence : _GEN_53 ? _slots_14_io_out_uop_is_fence : _GEN_52 ? _slots_13_io_out_uop_is_fence : _slots_12_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_54 ? _slots_15_io_out_uop_is_fencei : _GEN_53 ? _slots_14_io_out_uop_is_fencei : _GEN_52 ? _slots_13_io_out_uop_is_fencei : _slots_12_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_54 ? _slots_15_io_out_uop_is_amo : _GEN_53 ? _slots_14_io_out_uop_is_amo : _GEN_52 ? _slots_13_io_out_uop_is_amo : _slots_12_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_54 ? _slots_15_io_out_uop_uses_ldq : _GEN_53 ? _slots_14_io_out_uop_uses_ldq : _GEN_52 ? _slots_13_io_out_uop_uses_ldq : _slots_12_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_54 ? _slots_15_io_out_uop_uses_stq : _GEN_53 ? _slots_14_io_out_uop_uses_stq : _GEN_52 ? _slots_13_io_out_uop_uses_stq : _slots_12_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_54 ? _slots_15_io_out_uop_is_sys_pc2epc : _GEN_53 ? _slots_14_io_out_uop_is_sys_pc2epc : _GEN_52 ? _slots_13_io_out_uop_is_sys_pc2epc : _slots_12_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_54 ? _slots_15_io_out_uop_is_unique : _GEN_53 ? _slots_14_io_out_uop_is_unique : _GEN_52 ? _slots_13_io_out_uop_is_unique : _slots_12_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_54 ? _slots_15_io_out_uop_flush_on_commit : _GEN_53 ? _slots_14_io_out_uop_flush_on_commit : _GEN_52 ? _slots_13_io_out_uop_flush_on_commit : _slots_12_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_54 ? _slots_15_io_out_uop_ldst_is_rs1 : _GEN_53 ? _slots_14_io_out_uop_ldst_is_rs1 : _GEN_52 ? _slots_13_io_out_uop_ldst_is_rs1 : _slots_12_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_54 ? _slots_15_io_out_uop_ldst : _GEN_53 ? _slots_14_io_out_uop_ldst : _GEN_52 ? _slots_13_io_out_uop_ldst : _slots_12_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_54 ? _slots_15_io_out_uop_lrs1 : _GEN_53 ? _slots_14_io_out_uop_lrs1 : _GEN_52 ? _slots_13_io_out_uop_lrs1 : _slots_12_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_54 ? _slots_15_io_out_uop_lrs2 : _GEN_53 ? _slots_14_io_out_uop_lrs2 : _GEN_52 ? _slots_13_io_out_uop_lrs2 : _slots_12_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_54 ? _slots_15_io_out_uop_lrs3 : _GEN_53 ? _slots_14_io_out_uop_lrs3 : _GEN_52 ? _slots_13_io_out_uop_lrs3 : _slots_12_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_54 ? _slots_15_io_out_uop_ldst_val : _GEN_53 ? _slots_14_io_out_uop_ldst_val : _GEN_52 ? _slots_13_io_out_uop_ldst_val : _slots_12_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_54 ? _slots_15_io_out_uop_dst_rtype : _GEN_53 ? _slots_14_io_out_uop_dst_rtype : _GEN_52 ? _slots_13_io_out_uop_dst_rtype : _slots_12_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_54 ? _slots_15_io_out_uop_lrs1_rtype : _GEN_53 ? _slots_14_io_out_uop_lrs1_rtype : _GEN_52 ? _slots_13_io_out_uop_lrs1_rtype : _slots_12_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_54 ? _slots_15_io_out_uop_lrs2_rtype : _GEN_53 ? _slots_14_io_out_uop_lrs2_rtype : _GEN_52 ? _slots_13_io_out_uop_lrs2_rtype : _slots_12_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_54 ? _slots_15_io_out_uop_frs3_en : _GEN_53 ? _slots_14_io_out_uop_frs3_en : _GEN_52 ? _slots_13_io_out_uop_frs3_en : _slots_12_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_54 ? _slots_15_io_out_uop_fp_val : _GEN_53 ? _slots_14_io_out_uop_fp_val : _GEN_52 ? _slots_13_io_out_uop_fp_val : _slots_12_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_54 ? _slots_15_io_out_uop_fp_single : _GEN_53 ? _slots_14_io_out_uop_fp_single : _GEN_52 ? _slots_13_io_out_uop_fp_single : _slots_12_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_54 ? _slots_15_io_out_uop_xcpt_pf_if : _GEN_53 ? _slots_14_io_out_uop_xcpt_pf_if : _GEN_52 ? _slots_13_io_out_uop_xcpt_pf_if : _slots_12_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_54 ? _slots_15_io_out_uop_xcpt_ae_if : _GEN_53 ? _slots_14_io_out_uop_xcpt_ae_if : _GEN_52 ? _slots_13_io_out_uop_xcpt_ae_if : _slots_12_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_54 ? _slots_15_io_out_uop_xcpt_ma_if : _GEN_53 ? _slots_14_io_out_uop_xcpt_ma_if : _GEN_52 ? _slots_13_io_out_uop_xcpt_ma_if : _slots_12_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_54 ? _slots_15_io_out_uop_bp_debug_if : _GEN_53 ? _slots_14_io_out_uop_bp_debug_if : _GEN_52 ? _slots_13_io_out_uop_bp_debug_if : _slots_12_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_54 ? _slots_15_io_out_uop_bp_xcpt_if : _GEN_53 ? _slots_14_io_out_uop_bp_xcpt_if : _GEN_52 ? _slots_13_io_out_uop_bp_xcpt_if : _slots_12_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_54 ? _slots_15_io_out_uop_debug_fsrc : _GEN_53 ? _slots_14_io_out_uop_debug_fsrc : _GEN_52 ? _slots_13_io_out_uop_debug_fsrc : _slots_12_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_54 ? _slots_15_io_out_uop_debug_tsrc : _GEN_53 ? _slots_14_io_out_uop_debug_tsrc : _GEN_52 ? _slots_13_io_out_uop_debug_tsrc : _slots_12_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_11_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_11_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_11_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_11_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_11_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_11_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_11_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_11_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_11_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_11_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_11_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_11_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_11_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_11_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_11_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_11_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_11_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_11_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_11_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_11_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_11_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_11_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_11_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_11_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_11_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_11_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_11_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_11_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_11_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_11_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_11_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_11_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_11_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_11_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_11_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_11_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_11_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_11_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_11_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_11_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_11_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_11_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_11_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_11_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_11_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_11_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_11_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_11_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_11_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_11_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_11_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_11_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_11_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_11_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_11_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_11_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_11_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_11_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_11_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_11_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_11_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_11_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_11_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_11_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_11_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_11_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_11_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_11_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_11_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_11_io_uop_uopc),
    .io_uop_inst                    (_slots_11_io_uop_inst),
    .io_uop_debug_inst              (_slots_11_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_11_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_11_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_11_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_11_io_uop_fu_code),
    .io_uop_iw_state                (_slots_11_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_11_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_11_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_11_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_11_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_11_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_11_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_11_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_11_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_11_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_11_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_11_io_uop_pc_lob),
    .io_uop_taken                   (_slots_11_io_uop_taken),
    .io_uop_imm_packed              (_slots_11_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_11_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_11_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_11_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_11_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_11_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_11_io_uop_pdst),
    .io_uop_prs1                    (_slots_11_io_uop_prs1),
    .io_uop_prs2                    (_slots_11_io_uop_prs2),
    .io_uop_prs3                    (_slots_11_io_uop_prs3),
    .io_uop_ppred                   (_slots_11_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_11_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_11_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_11_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_11_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_11_io_uop_stale_pdst),
    .io_uop_exception               (_slots_11_io_uop_exception),
    .io_uop_exc_cause               (_slots_11_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_11_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_11_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_11_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_11_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_11_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_11_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_11_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_11_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_11_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_11_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_11_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_11_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_11_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_11_io_uop_ldst),
    .io_uop_lrs1                    (_slots_11_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_11_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_11_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_11_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_11_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_11_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_11_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_11_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_11_io_uop_fp_val),
    .io_uop_fp_single               (_slots_11_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_11_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_11_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_11_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_11_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_11_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_11_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_11_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_12 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_12_io_valid),
    .io_will_be_valid               (_slots_12_io_will_be_valid),
    .io_request                     (_slots_12_io_request),
    .io_grant                       (issue_slots_12_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_11),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_12_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_57 ? _slots_16_io_out_uop_uopc : _GEN_56 ? _slots_15_io_out_uop_uopc : _GEN_55 ? _slots_14_io_out_uop_uopc : _slots_13_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_57 ? _slots_16_io_out_uop_inst : _GEN_56 ? _slots_15_io_out_uop_inst : _GEN_55 ? _slots_14_io_out_uop_inst : _slots_13_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_57 ? _slots_16_io_out_uop_debug_inst : _GEN_56 ? _slots_15_io_out_uop_debug_inst : _GEN_55 ? _slots_14_io_out_uop_debug_inst : _slots_13_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_57 ? _slots_16_io_out_uop_is_rvc : _GEN_56 ? _slots_15_io_out_uop_is_rvc : _GEN_55 ? _slots_14_io_out_uop_is_rvc : _slots_13_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_57 ? _slots_16_io_out_uop_debug_pc : _GEN_56 ? _slots_15_io_out_uop_debug_pc : _GEN_55 ? _slots_14_io_out_uop_debug_pc : _slots_13_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_57 ? _slots_16_io_out_uop_iq_type : _GEN_56 ? _slots_15_io_out_uop_iq_type : _GEN_55 ? _slots_14_io_out_uop_iq_type : _slots_13_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_57 ? _slots_16_io_out_uop_fu_code : _GEN_56 ? _slots_15_io_out_uop_fu_code : _GEN_55 ? _slots_14_io_out_uop_fu_code : _slots_13_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_57 ? _slots_16_io_out_uop_iw_state : _GEN_56 ? _slots_15_io_out_uop_iw_state : _GEN_55 ? _slots_14_io_out_uop_iw_state : _slots_13_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_57 ? _slots_16_io_out_uop_iw_p1_poisoned : _GEN_56 ? _slots_15_io_out_uop_iw_p1_poisoned : _GEN_55 ? _slots_14_io_out_uop_iw_p1_poisoned : _slots_13_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_57 ? _slots_16_io_out_uop_iw_p2_poisoned : _GEN_56 ? _slots_15_io_out_uop_iw_p2_poisoned : _GEN_55 ? _slots_14_io_out_uop_iw_p2_poisoned : _slots_13_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_57 ? _slots_16_io_out_uop_is_br : _GEN_56 ? _slots_15_io_out_uop_is_br : _GEN_55 ? _slots_14_io_out_uop_is_br : _slots_13_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_57 ? _slots_16_io_out_uop_is_jalr : _GEN_56 ? _slots_15_io_out_uop_is_jalr : _GEN_55 ? _slots_14_io_out_uop_is_jalr : _slots_13_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_57 ? _slots_16_io_out_uop_is_jal : _GEN_56 ? _slots_15_io_out_uop_is_jal : _GEN_55 ? _slots_14_io_out_uop_is_jal : _slots_13_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_57 ? _slots_16_io_out_uop_is_sfb : _GEN_56 ? _slots_15_io_out_uop_is_sfb : _GEN_55 ? _slots_14_io_out_uop_is_sfb : _slots_13_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_57 ? _slots_16_io_out_uop_br_mask : _GEN_56 ? _slots_15_io_out_uop_br_mask : _GEN_55 ? _slots_14_io_out_uop_br_mask : _slots_13_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_57 ? _slots_16_io_out_uop_br_tag : _GEN_56 ? _slots_15_io_out_uop_br_tag : _GEN_55 ? _slots_14_io_out_uop_br_tag : _slots_13_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_57 ? _slots_16_io_out_uop_ftq_idx : _GEN_56 ? _slots_15_io_out_uop_ftq_idx : _GEN_55 ? _slots_14_io_out_uop_ftq_idx : _slots_13_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_57 ? _slots_16_io_out_uop_edge_inst : _GEN_56 ? _slots_15_io_out_uop_edge_inst : _GEN_55 ? _slots_14_io_out_uop_edge_inst : _slots_13_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_57 ? _slots_16_io_out_uop_pc_lob : _GEN_56 ? _slots_15_io_out_uop_pc_lob : _GEN_55 ? _slots_14_io_out_uop_pc_lob : _slots_13_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_57 ? _slots_16_io_out_uop_taken : _GEN_56 ? _slots_15_io_out_uop_taken : _GEN_55 ? _slots_14_io_out_uop_taken : _slots_13_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_57 ? _slots_16_io_out_uop_imm_packed : _GEN_56 ? _slots_15_io_out_uop_imm_packed : _GEN_55 ? _slots_14_io_out_uop_imm_packed : _slots_13_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_57 ? _slots_16_io_out_uop_csr_addr : _GEN_56 ? _slots_15_io_out_uop_csr_addr : _GEN_55 ? _slots_14_io_out_uop_csr_addr : _slots_13_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_57 ? _slots_16_io_out_uop_rob_idx : _GEN_56 ? _slots_15_io_out_uop_rob_idx : _GEN_55 ? _slots_14_io_out_uop_rob_idx : _slots_13_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_57 ? _slots_16_io_out_uop_ldq_idx : _GEN_56 ? _slots_15_io_out_uop_ldq_idx : _GEN_55 ? _slots_14_io_out_uop_ldq_idx : _slots_13_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_57 ? _slots_16_io_out_uop_stq_idx : _GEN_56 ? _slots_15_io_out_uop_stq_idx : _GEN_55 ? _slots_14_io_out_uop_stq_idx : _slots_13_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_57 ? _slots_16_io_out_uop_rxq_idx : _GEN_56 ? _slots_15_io_out_uop_rxq_idx : _GEN_55 ? _slots_14_io_out_uop_rxq_idx : _slots_13_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_57 ? _slots_16_io_out_uop_pdst : _GEN_56 ? _slots_15_io_out_uop_pdst : _GEN_55 ? _slots_14_io_out_uop_pdst : _slots_13_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_57 ? _slots_16_io_out_uop_prs1 : _GEN_56 ? _slots_15_io_out_uop_prs1 : _GEN_55 ? _slots_14_io_out_uop_prs1 : _slots_13_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_57 ? _slots_16_io_out_uop_prs2 : _GEN_56 ? _slots_15_io_out_uop_prs2 : _GEN_55 ? _slots_14_io_out_uop_prs2 : _slots_13_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_57 ? _slots_16_io_out_uop_prs3 : _GEN_56 ? _slots_15_io_out_uop_prs3 : _GEN_55 ? _slots_14_io_out_uop_prs3 : _slots_13_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_57 ? _slots_16_io_out_uop_ppred : _GEN_56 ? _slots_15_io_out_uop_ppred : _GEN_55 ? _slots_14_io_out_uop_ppred : _slots_13_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_57 ? _slots_16_io_out_uop_prs1_busy : _GEN_56 ? _slots_15_io_out_uop_prs1_busy : _GEN_55 ? _slots_14_io_out_uop_prs1_busy : _slots_13_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_57 ? _slots_16_io_out_uop_prs2_busy : _GEN_56 ? _slots_15_io_out_uop_prs2_busy : _GEN_55 ? _slots_14_io_out_uop_prs2_busy : _slots_13_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_57 ? _slots_16_io_out_uop_prs3_busy : _GEN_56 ? _slots_15_io_out_uop_prs3_busy : _GEN_55 ? _slots_14_io_out_uop_prs3_busy : _slots_13_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_57 ? _slots_16_io_out_uop_ppred_busy : _GEN_56 ? _slots_15_io_out_uop_ppred_busy : _GEN_55 ? _slots_14_io_out_uop_ppred_busy : _slots_13_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_57 ? _slots_16_io_out_uop_stale_pdst : _GEN_56 ? _slots_15_io_out_uop_stale_pdst : _GEN_55 ? _slots_14_io_out_uop_stale_pdst : _slots_13_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_57 ? _slots_16_io_out_uop_exception : _GEN_56 ? _slots_15_io_out_uop_exception : _GEN_55 ? _slots_14_io_out_uop_exception : _slots_13_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_57 ? _slots_16_io_out_uop_exc_cause : _GEN_56 ? _slots_15_io_out_uop_exc_cause : _GEN_55 ? _slots_14_io_out_uop_exc_cause : _slots_13_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_57 ? _slots_16_io_out_uop_bypassable : _GEN_56 ? _slots_15_io_out_uop_bypassable : _GEN_55 ? _slots_14_io_out_uop_bypassable : _slots_13_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_57 ? _slots_16_io_out_uop_mem_cmd : _GEN_56 ? _slots_15_io_out_uop_mem_cmd : _GEN_55 ? _slots_14_io_out_uop_mem_cmd : _slots_13_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_57 ? _slots_16_io_out_uop_mem_size : _GEN_56 ? _slots_15_io_out_uop_mem_size : _GEN_55 ? _slots_14_io_out_uop_mem_size : _slots_13_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_57 ? _slots_16_io_out_uop_mem_signed : _GEN_56 ? _slots_15_io_out_uop_mem_signed : _GEN_55 ? _slots_14_io_out_uop_mem_signed : _slots_13_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_57 ? _slots_16_io_out_uop_is_fence : _GEN_56 ? _slots_15_io_out_uop_is_fence : _GEN_55 ? _slots_14_io_out_uop_is_fence : _slots_13_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_57 ? _slots_16_io_out_uop_is_fencei : _GEN_56 ? _slots_15_io_out_uop_is_fencei : _GEN_55 ? _slots_14_io_out_uop_is_fencei : _slots_13_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_57 ? _slots_16_io_out_uop_is_amo : _GEN_56 ? _slots_15_io_out_uop_is_amo : _GEN_55 ? _slots_14_io_out_uop_is_amo : _slots_13_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_57 ? _slots_16_io_out_uop_uses_ldq : _GEN_56 ? _slots_15_io_out_uop_uses_ldq : _GEN_55 ? _slots_14_io_out_uop_uses_ldq : _slots_13_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_57 ? _slots_16_io_out_uop_uses_stq : _GEN_56 ? _slots_15_io_out_uop_uses_stq : _GEN_55 ? _slots_14_io_out_uop_uses_stq : _slots_13_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_57 ? _slots_16_io_out_uop_is_sys_pc2epc : _GEN_56 ? _slots_15_io_out_uop_is_sys_pc2epc : _GEN_55 ? _slots_14_io_out_uop_is_sys_pc2epc : _slots_13_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_57 ? _slots_16_io_out_uop_is_unique : _GEN_56 ? _slots_15_io_out_uop_is_unique : _GEN_55 ? _slots_14_io_out_uop_is_unique : _slots_13_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_57 ? _slots_16_io_out_uop_flush_on_commit : _GEN_56 ? _slots_15_io_out_uop_flush_on_commit : _GEN_55 ? _slots_14_io_out_uop_flush_on_commit : _slots_13_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_57 ? _slots_16_io_out_uop_ldst_is_rs1 : _GEN_56 ? _slots_15_io_out_uop_ldst_is_rs1 : _GEN_55 ? _slots_14_io_out_uop_ldst_is_rs1 : _slots_13_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_57 ? _slots_16_io_out_uop_ldst : _GEN_56 ? _slots_15_io_out_uop_ldst : _GEN_55 ? _slots_14_io_out_uop_ldst : _slots_13_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_57 ? _slots_16_io_out_uop_lrs1 : _GEN_56 ? _slots_15_io_out_uop_lrs1 : _GEN_55 ? _slots_14_io_out_uop_lrs1 : _slots_13_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_57 ? _slots_16_io_out_uop_lrs2 : _GEN_56 ? _slots_15_io_out_uop_lrs2 : _GEN_55 ? _slots_14_io_out_uop_lrs2 : _slots_13_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_57 ? _slots_16_io_out_uop_lrs3 : _GEN_56 ? _slots_15_io_out_uop_lrs3 : _GEN_55 ? _slots_14_io_out_uop_lrs3 : _slots_13_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_57 ? _slots_16_io_out_uop_ldst_val : _GEN_56 ? _slots_15_io_out_uop_ldst_val : _GEN_55 ? _slots_14_io_out_uop_ldst_val : _slots_13_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_57 ? _slots_16_io_out_uop_dst_rtype : _GEN_56 ? _slots_15_io_out_uop_dst_rtype : _GEN_55 ? _slots_14_io_out_uop_dst_rtype : _slots_13_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_57 ? _slots_16_io_out_uop_lrs1_rtype : _GEN_56 ? _slots_15_io_out_uop_lrs1_rtype : _GEN_55 ? _slots_14_io_out_uop_lrs1_rtype : _slots_13_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_57 ? _slots_16_io_out_uop_lrs2_rtype : _GEN_56 ? _slots_15_io_out_uop_lrs2_rtype : _GEN_55 ? _slots_14_io_out_uop_lrs2_rtype : _slots_13_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_57 ? _slots_16_io_out_uop_frs3_en : _GEN_56 ? _slots_15_io_out_uop_frs3_en : _GEN_55 ? _slots_14_io_out_uop_frs3_en : _slots_13_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_57 ? _slots_16_io_out_uop_fp_val : _GEN_56 ? _slots_15_io_out_uop_fp_val : _GEN_55 ? _slots_14_io_out_uop_fp_val : _slots_13_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_57 ? _slots_16_io_out_uop_fp_single : _GEN_56 ? _slots_15_io_out_uop_fp_single : _GEN_55 ? _slots_14_io_out_uop_fp_single : _slots_13_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_57 ? _slots_16_io_out_uop_xcpt_pf_if : _GEN_56 ? _slots_15_io_out_uop_xcpt_pf_if : _GEN_55 ? _slots_14_io_out_uop_xcpt_pf_if : _slots_13_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_57 ? _slots_16_io_out_uop_xcpt_ae_if : _GEN_56 ? _slots_15_io_out_uop_xcpt_ae_if : _GEN_55 ? _slots_14_io_out_uop_xcpt_ae_if : _slots_13_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_57 ? _slots_16_io_out_uop_xcpt_ma_if : _GEN_56 ? _slots_15_io_out_uop_xcpt_ma_if : _GEN_55 ? _slots_14_io_out_uop_xcpt_ma_if : _slots_13_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_57 ? _slots_16_io_out_uop_bp_debug_if : _GEN_56 ? _slots_15_io_out_uop_bp_debug_if : _GEN_55 ? _slots_14_io_out_uop_bp_debug_if : _slots_13_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_57 ? _slots_16_io_out_uop_bp_xcpt_if : _GEN_56 ? _slots_15_io_out_uop_bp_xcpt_if : _GEN_55 ? _slots_14_io_out_uop_bp_xcpt_if : _slots_13_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_57 ? _slots_16_io_out_uop_debug_fsrc : _GEN_56 ? _slots_15_io_out_uop_debug_fsrc : _GEN_55 ? _slots_14_io_out_uop_debug_fsrc : _slots_13_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_57 ? _slots_16_io_out_uop_debug_tsrc : _GEN_56 ? _slots_15_io_out_uop_debug_tsrc : _GEN_55 ? _slots_14_io_out_uop_debug_tsrc : _slots_13_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_12_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_12_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_12_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_12_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_12_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_12_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_12_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_12_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_12_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_12_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_12_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_12_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_12_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_12_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_12_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_12_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_12_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_12_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_12_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_12_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_12_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_12_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_12_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_12_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_12_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_12_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_12_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_12_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_12_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_12_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_12_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_12_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_12_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_12_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_12_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_12_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_12_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_12_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_12_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_12_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_12_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_12_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_12_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_12_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_12_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_12_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_12_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_12_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_12_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_12_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_12_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_12_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_12_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_12_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_12_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_12_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_12_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_12_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_12_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_12_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_12_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_12_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_12_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_12_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_12_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_12_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_12_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_12_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_12_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_12_io_uop_uopc),
    .io_uop_inst                    (_slots_12_io_uop_inst),
    .io_uop_debug_inst              (_slots_12_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_12_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_12_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_12_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_12_io_uop_fu_code),
    .io_uop_iw_state                (_slots_12_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_12_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_12_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_12_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_12_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_12_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_12_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_12_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_12_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_12_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_12_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_12_io_uop_pc_lob),
    .io_uop_taken                   (_slots_12_io_uop_taken),
    .io_uop_imm_packed              (_slots_12_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_12_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_12_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_12_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_12_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_12_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_12_io_uop_pdst),
    .io_uop_prs1                    (_slots_12_io_uop_prs1),
    .io_uop_prs2                    (_slots_12_io_uop_prs2),
    .io_uop_prs3                    (_slots_12_io_uop_prs3),
    .io_uop_ppred                   (_slots_12_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_12_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_12_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_12_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_12_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_12_io_uop_stale_pdst),
    .io_uop_exception               (_slots_12_io_uop_exception),
    .io_uop_exc_cause               (_slots_12_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_12_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_12_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_12_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_12_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_12_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_12_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_12_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_12_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_12_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_12_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_12_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_12_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_12_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_12_io_uop_ldst),
    .io_uop_lrs1                    (_slots_12_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_12_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_12_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_12_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_12_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_12_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_12_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_12_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_12_io_uop_fp_val),
    .io_uop_fp_single               (_slots_12_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_12_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_12_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_12_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_12_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_12_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_12_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_12_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_13 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_13_io_valid),
    .io_will_be_valid               (_slots_13_io_will_be_valid),
    .io_request                     (_slots_13_io_request),
    .io_grant                       (issue_slots_13_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_12),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_13_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_60 ? _slots_17_io_out_uop_uopc : _GEN_59 ? _slots_16_io_out_uop_uopc : _GEN_58 ? _slots_15_io_out_uop_uopc : _slots_14_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_60 ? _slots_17_io_out_uop_inst : _GEN_59 ? _slots_16_io_out_uop_inst : _GEN_58 ? _slots_15_io_out_uop_inst : _slots_14_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_60 ? _slots_17_io_out_uop_debug_inst : _GEN_59 ? _slots_16_io_out_uop_debug_inst : _GEN_58 ? _slots_15_io_out_uop_debug_inst : _slots_14_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_60 ? _slots_17_io_out_uop_is_rvc : _GEN_59 ? _slots_16_io_out_uop_is_rvc : _GEN_58 ? _slots_15_io_out_uop_is_rvc : _slots_14_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_60 ? _slots_17_io_out_uop_debug_pc : _GEN_59 ? _slots_16_io_out_uop_debug_pc : _GEN_58 ? _slots_15_io_out_uop_debug_pc : _slots_14_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_60 ? _slots_17_io_out_uop_iq_type : _GEN_59 ? _slots_16_io_out_uop_iq_type : _GEN_58 ? _slots_15_io_out_uop_iq_type : _slots_14_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_60 ? _slots_17_io_out_uop_fu_code : _GEN_59 ? _slots_16_io_out_uop_fu_code : _GEN_58 ? _slots_15_io_out_uop_fu_code : _slots_14_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_60 ? _slots_17_io_out_uop_iw_state : _GEN_59 ? _slots_16_io_out_uop_iw_state : _GEN_58 ? _slots_15_io_out_uop_iw_state : _slots_14_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_60 ? _slots_17_io_out_uop_iw_p1_poisoned : _GEN_59 ? _slots_16_io_out_uop_iw_p1_poisoned : _GEN_58 ? _slots_15_io_out_uop_iw_p1_poisoned : _slots_14_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_60 ? _slots_17_io_out_uop_iw_p2_poisoned : _GEN_59 ? _slots_16_io_out_uop_iw_p2_poisoned : _GEN_58 ? _slots_15_io_out_uop_iw_p2_poisoned : _slots_14_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_60 ? _slots_17_io_out_uop_is_br : _GEN_59 ? _slots_16_io_out_uop_is_br : _GEN_58 ? _slots_15_io_out_uop_is_br : _slots_14_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_60 ? _slots_17_io_out_uop_is_jalr : _GEN_59 ? _slots_16_io_out_uop_is_jalr : _GEN_58 ? _slots_15_io_out_uop_is_jalr : _slots_14_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_60 ? _slots_17_io_out_uop_is_jal : _GEN_59 ? _slots_16_io_out_uop_is_jal : _GEN_58 ? _slots_15_io_out_uop_is_jal : _slots_14_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_60 ? _slots_17_io_out_uop_is_sfb : _GEN_59 ? _slots_16_io_out_uop_is_sfb : _GEN_58 ? _slots_15_io_out_uop_is_sfb : _slots_14_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_60 ? _slots_17_io_out_uop_br_mask : _GEN_59 ? _slots_16_io_out_uop_br_mask : _GEN_58 ? _slots_15_io_out_uop_br_mask : _slots_14_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_60 ? _slots_17_io_out_uop_br_tag : _GEN_59 ? _slots_16_io_out_uop_br_tag : _GEN_58 ? _slots_15_io_out_uop_br_tag : _slots_14_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_60 ? _slots_17_io_out_uop_ftq_idx : _GEN_59 ? _slots_16_io_out_uop_ftq_idx : _GEN_58 ? _slots_15_io_out_uop_ftq_idx : _slots_14_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_60 ? _slots_17_io_out_uop_edge_inst : _GEN_59 ? _slots_16_io_out_uop_edge_inst : _GEN_58 ? _slots_15_io_out_uop_edge_inst : _slots_14_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_60 ? _slots_17_io_out_uop_pc_lob : _GEN_59 ? _slots_16_io_out_uop_pc_lob : _GEN_58 ? _slots_15_io_out_uop_pc_lob : _slots_14_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_60 ? _slots_17_io_out_uop_taken : _GEN_59 ? _slots_16_io_out_uop_taken : _GEN_58 ? _slots_15_io_out_uop_taken : _slots_14_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_60 ? _slots_17_io_out_uop_imm_packed : _GEN_59 ? _slots_16_io_out_uop_imm_packed : _GEN_58 ? _slots_15_io_out_uop_imm_packed : _slots_14_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_60 ? _slots_17_io_out_uop_csr_addr : _GEN_59 ? _slots_16_io_out_uop_csr_addr : _GEN_58 ? _slots_15_io_out_uop_csr_addr : _slots_14_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_60 ? _slots_17_io_out_uop_rob_idx : _GEN_59 ? _slots_16_io_out_uop_rob_idx : _GEN_58 ? _slots_15_io_out_uop_rob_idx : _slots_14_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_60 ? _slots_17_io_out_uop_ldq_idx : _GEN_59 ? _slots_16_io_out_uop_ldq_idx : _GEN_58 ? _slots_15_io_out_uop_ldq_idx : _slots_14_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_60 ? _slots_17_io_out_uop_stq_idx : _GEN_59 ? _slots_16_io_out_uop_stq_idx : _GEN_58 ? _slots_15_io_out_uop_stq_idx : _slots_14_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_60 ? _slots_17_io_out_uop_rxq_idx : _GEN_59 ? _slots_16_io_out_uop_rxq_idx : _GEN_58 ? _slots_15_io_out_uop_rxq_idx : _slots_14_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_60 ? _slots_17_io_out_uop_pdst : _GEN_59 ? _slots_16_io_out_uop_pdst : _GEN_58 ? _slots_15_io_out_uop_pdst : _slots_14_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_60 ? _slots_17_io_out_uop_prs1 : _GEN_59 ? _slots_16_io_out_uop_prs1 : _GEN_58 ? _slots_15_io_out_uop_prs1 : _slots_14_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_60 ? _slots_17_io_out_uop_prs2 : _GEN_59 ? _slots_16_io_out_uop_prs2 : _GEN_58 ? _slots_15_io_out_uop_prs2 : _slots_14_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_60 ? _slots_17_io_out_uop_prs3 : _GEN_59 ? _slots_16_io_out_uop_prs3 : _GEN_58 ? _slots_15_io_out_uop_prs3 : _slots_14_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_60 ? _slots_17_io_out_uop_ppred : _GEN_59 ? _slots_16_io_out_uop_ppred : _GEN_58 ? _slots_15_io_out_uop_ppred : _slots_14_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_60 ? _slots_17_io_out_uop_prs1_busy : _GEN_59 ? _slots_16_io_out_uop_prs1_busy : _GEN_58 ? _slots_15_io_out_uop_prs1_busy : _slots_14_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_60 ? _slots_17_io_out_uop_prs2_busy : _GEN_59 ? _slots_16_io_out_uop_prs2_busy : _GEN_58 ? _slots_15_io_out_uop_prs2_busy : _slots_14_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_60 ? _slots_17_io_out_uop_prs3_busy : _GEN_59 ? _slots_16_io_out_uop_prs3_busy : _GEN_58 ? _slots_15_io_out_uop_prs3_busy : _slots_14_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_60 ? _slots_17_io_out_uop_ppred_busy : _GEN_59 ? _slots_16_io_out_uop_ppred_busy : _GEN_58 ? _slots_15_io_out_uop_ppred_busy : _slots_14_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_60 ? _slots_17_io_out_uop_stale_pdst : _GEN_59 ? _slots_16_io_out_uop_stale_pdst : _GEN_58 ? _slots_15_io_out_uop_stale_pdst : _slots_14_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_60 ? _slots_17_io_out_uop_exception : _GEN_59 ? _slots_16_io_out_uop_exception : _GEN_58 ? _slots_15_io_out_uop_exception : _slots_14_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_60 ? _slots_17_io_out_uop_exc_cause : _GEN_59 ? _slots_16_io_out_uop_exc_cause : _GEN_58 ? _slots_15_io_out_uop_exc_cause : _slots_14_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_60 ? _slots_17_io_out_uop_bypassable : _GEN_59 ? _slots_16_io_out_uop_bypassable : _GEN_58 ? _slots_15_io_out_uop_bypassable : _slots_14_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_60 ? _slots_17_io_out_uop_mem_cmd : _GEN_59 ? _slots_16_io_out_uop_mem_cmd : _GEN_58 ? _slots_15_io_out_uop_mem_cmd : _slots_14_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_60 ? _slots_17_io_out_uop_mem_size : _GEN_59 ? _slots_16_io_out_uop_mem_size : _GEN_58 ? _slots_15_io_out_uop_mem_size : _slots_14_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_60 ? _slots_17_io_out_uop_mem_signed : _GEN_59 ? _slots_16_io_out_uop_mem_signed : _GEN_58 ? _slots_15_io_out_uop_mem_signed : _slots_14_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_60 ? _slots_17_io_out_uop_is_fence : _GEN_59 ? _slots_16_io_out_uop_is_fence : _GEN_58 ? _slots_15_io_out_uop_is_fence : _slots_14_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_60 ? _slots_17_io_out_uop_is_fencei : _GEN_59 ? _slots_16_io_out_uop_is_fencei : _GEN_58 ? _slots_15_io_out_uop_is_fencei : _slots_14_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_60 ? _slots_17_io_out_uop_is_amo : _GEN_59 ? _slots_16_io_out_uop_is_amo : _GEN_58 ? _slots_15_io_out_uop_is_amo : _slots_14_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_60 ? _slots_17_io_out_uop_uses_ldq : _GEN_59 ? _slots_16_io_out_uop_uses_ldq : _GEN_58 ? _slots_15_io_out_uop_uses_ldq : _slots_14_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_60 ? _slots_17_io_out_uop_uses_stq : _GEN_59 ? _slots_16_io_out_uop_uses_stq : _GEN_58 ? _slots_15_io_out_uop_uses_stq : _slots_14_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_60 ? _slots_17_io_out_uop_is_sys_pc2epc : _GEN_59 ? _slots_16_io_out_uop_is_sys_pc2epc : _GEN_58 ? _slots_15_io_out_uop_is_sys_pc2epc : _slots_14_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_60 ? _slots_17_io_out_uop_is_unique : _GEN_59 ? _slots_16_io_out_uop_is_unique : _GEN_58 ? _slots_15_io_out_uop_is_unique : _slots_14_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_60 ? _slots_17_io_out_uop_flush_on_commit : _GEN_59 ? _slots_16_io_out_uop_flush_on_commit : _GEN_58 ? _slots_15_io_out_uop_flush_on_commit : _slots_14_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_60 ? _slots_17_io_out_uop_ldst_is_rs1 : _GEN_59 ? _slots_16_io_out_uop_ldst_is_rs1 : _GEN_58 ? _slots_15_io_out_uop_ldst_is_rs1 : _slots_14_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_60 ? _slots_17_io_out_uop_ldst : _GEN_59 ? _slots_16_io_out_uop_ldst : _GEN_58 ? _slots_15_io_out_uop_ldst : _slots_14_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_60 ? _slots_17_io_out_uop_lrs1 : _GEN_59 ? _slots_16_io_out_uop_lrs1 : _GEN_58 ? _slots_15_io_out_uop_lrs1 : _slots_14_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_60 ? _slots_17_io_out_uop_lrs2 : _GEN_59 ? _slots_16_io_out_uop_lrs2 : _GEN_58 ? _slots_15_io_out_uop_lrs2 : _slots_14_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_60 ? _slots_17_io_out_uop_lrs3 : _GEN_59 ? _slots_16_io_out_uop_lrs3 : _GEN_58 ? _slots_15_io_out_uop_lrs3 : _slots_14_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_60 ? _slots_17_io_out_uop_ldst_val : _GEN_59 ? _slots_16_io_out_uop_ldst_val : _GEN_58 ? _slots_15_io_out_uop_ldst_val : _slots_14_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_60 ? _slots_17_io_out_uop_dst_rtype : _GEN_59 ? _slots_16_io_out_uop_dst_rtype : _GEN_58 ? _slots_15_io_out_uop_dst_rtype : _slots_14_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_60 ? _slots_17_io_out_uop_lrs1_rtype : _GEN_59 ? _slots_16_io_out_uop_lrs1_rtype : _GEN_58 ? _slots_15_io_out_uop_lrs1_rtype : _slots_14_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_60 ? _slots_17_io_out_uop_lrs2_rtype : _GEN_59 ? _slots_16_io_out_uop_lrs2_rtype : _GEN_58 ? _slots_15_io_out_uop_lrs2_rtype : _slots_14_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_60 ? _slots_17_io_out_uop_frs3_en : _GEN_59 ? _slots_16_io_out_uop_frs3_en : _GEN_58 ? _slots_15_io_out_uop_frs3_en : _slots_14_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_60 ? _slots_17_io_out_uop_fp_val : _GEN_59 ? _slots_16_io_out_uop_fp_val : _GEN_58 ? _slots_15_io_out_uop_fp_val : _slots_14_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_60 ? _slots_17_io_out_uop_fp_single : _GEN_59 ? _slots_16_io_out_uop_fp_single : _GEN_58 ? _slots_15_io_out_uop_fp_single : _slots_14_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_60 ? _slots_17_io_out_uop_xcpt_pf_if : _GEN_59 ? _slots_16_io_out_uop_xcpt_pf_if : _GEN_58 ? _slots_15_io_out_uop_xcpt_pf_if : _slots_14_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_60 ? _slots_17_io_out_uop_xcpt_ae_if : _GEN_59 ? _slots_16_io_out_uop_xcpt_ae_if : _GEN_58 ? _slots_15_io_out_uop_xcpt_ae_if : _slots_14_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_60 ? _slots_17_io_out_uop_xcpt_ma_if : _GEN_59 ? _slots_16_io_out_uop_xcpt_ma_if : _GEN_58 ? _slots_15_io_out_uop_xcpt_ma_if : _slots_14_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_60 ? _slots_17_io_out_uop_bp_debug_if : _GEN_59 ? _slots_16_io_out_uop_bp_debug_if : _GEN_58 ? _slots_15_io_out_uop_bp_debug_if : _slots_14_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_60 ? _slots_17_io_out_uop_bp_xcpt_if : _GEN_59 ? _slots_16_io_out_uop_bp_xcpt_if : _GEN_58 ? _slots_15_io_out_uop_bp_xcpt_if : _slots_14_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_60 ? _slots_17_io_out_uop_debug_fsrc : _GEN_59 ? _slots_16_io_out_uop_debug_fsrc : _GEN_58 ? _slots_15_io_out_uop_debug_fsrc : _slots_14_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_60 ? _slots_17_io_out_uop_debug_tsrc : _GEN_59 ? _slots_16_io_out_uop_debug_tsrc : _GEN_58 ? _slots_15_io_out_uop_debug_tsrc : _slots_14_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_13_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_13_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_13_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_13_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_13_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_13_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_13_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_13_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_13_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_13_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_13_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_13_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_13_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_13_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_13_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_13_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_13_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_13_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_13_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_13_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_13_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_13_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_13_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_13_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_13_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_13_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_13_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_13_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_13_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_13_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_13_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_13_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_13_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_13_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_13_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_13_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_13_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_13_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_13_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_13_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_13_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_13_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_13_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_13_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_13_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_13_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_13_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_13_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_13_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_13_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_13_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_13_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_13_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_13_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_13_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_13_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_13_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_13_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_13_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_13_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_13_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_13_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_13_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_13_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_13_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_13_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_13_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_13_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_13_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_13_io_uop_uopc),
    .io_uop_inst                    (_slots_13_io_uop_inst),
    .io_uop_debug_inst              (_slots_13_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_13_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_13_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_13_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_13_io_uop_fu_code),
    .io_uop_iw_state                (_slots_13_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_13_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_13_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_13_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_13_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_13_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_13_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_13_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_13_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_13_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_13_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_13_io_uop_pc_lob),
    .io_uop_taken                   (_slots_13_io_uop_taken),
    .io_uop_imm_packed              (_slots_13_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_13_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_13_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_13_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_13_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_13_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_13_io_uop_pdst),
    .io_uop_prs1                    (_slots_13_io_uop_prs1),
    .io_uop_prs2                    (_slots_13_io_uop_prs2),
    .io_uop_prs3                    (_slots_13_io_uop_prs3),
    .io_uop_ppred                   (_slots_13_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_13_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_13_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_13_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_13_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_13_io_uop_stale_pdst),
    .io_uop_exception               (_slots_13_io_uop_exception),
    .io_uop_exc_cause               (_slots_13_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_13_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_13_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_13_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_13_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_13_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_13_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_13_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_13_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_13_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_13_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_13_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_13_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_13_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_13_io_uop_ldst),
    .io_uop_lrs1                    (_slots_13_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_13_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_13_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_13_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_13_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_13_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_13_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_13_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_13_io_uop_fp_val),
    .io_uop_fp_single               (_slots_13_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_13_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_13_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_13_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_13_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_13_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_13_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_13_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_14 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_14_io_valid),
    .io_will_be_valid               (_slots_14_io_will_be_valid),
    .io_request                     (_slots_14_io_request),
    .io_grant                       (issue_slots_14_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_13),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_14_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_63 ? _slots_18_io_out_uop_uopc : _GEN_62 ? _slots_17_io_out_uop_uopc : _GEN_61 ? _slots_16_io_out_uop_uopc : _slots_15_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_63 ? _slots_18_io_out_uop_inst : _GEN_62 ? _slots_17_io_out_uop_inst : _GEN_61 ? _slots_16_io_out_uop_inst : _slots_15_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_63 ? _slots_18_io_out_uop_debug_inst : _GEN_62 ? _slots_17_io_out_uop_debug_inst : _GEN_61 ? _slots_16_io_out_uop_debug_inst : _slots_15_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_63 ? _slots_18_io_out_uop_is_rvc : _GEN_62 ? _slots_17_io_out_uop_is_rvc : _GEN_61 ? _slots_16_io_out_uop_is_rvc : _slots_15_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_63 ? _slots_18_io_out_uop_debug_pc : _GEN_62 ? _slots_17_io_out_uop_debug_pc : _GEN_61 ? _slots_16_io_out_uop_debug_pc : _slots_15_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_63 ? _slots_18_io_out_uop_iq_type : _GEN_62 ? _slots_17_io_out_uop_iq_type : _GEN_61 ? _slots_16_io_out_uop_iq_type : _slots_15_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_63 ? _slots_18_io_out_uop_fu_code : _GEN_62 ? _slots_17_io_out_uop_fu_code : _GEN_61 ? _slots_16_io_out_uop_fu_code : _slots_15_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_63 ? _slots_18_io_out_uop_iw_state : _GEN_62 ? _slots_17_io_out_uop_iw_state : _GEN_61 ? _slots_16_io_out_uop_iw_state : _slots_15_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_63 ? _slots_18_io_out_uop_iw_p1_poisoned : _GEN_62 ? _slots_17_io_out_uop_iw_p1_poisoned : _GEN_61 ? _slots_16_io_out_uop_iw_p1_poisoned : _slots_15_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_63 ? _slots_18_io_out_uop_iw_p2_poisoned : _GEN_62 ? _slots_17_io_out_uop_iw_p2_poisoned : _GEN_61 ? _slots_16_io_out_uop_iw_p2_poisoned : _slots_15_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_63 ? _slots_18_io_out_uop_is_br : _GEN_62 ? _slots_17_io_out_uop_is_br : _GEN_61 ? _slots_16_io_out_uop_is_br : _slots_15_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_63 ? _slots_18_io_out_uop_is_jalr : _GEN_62 ? _slots_17_io_out_uop_is_jalr : _GEN_61 ? _slots_16_io_out_uop_is_jalr : _slots_15_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_63 ? _slots_18_io_out_uop_is_jal : _GEN_62 ? _slots_17_io_out_uop_is_jal : _GEN_61 ? _slots_16_io_out_uop_is_jal : _slots_15_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_63 ? _slots_18_io_out_uop_is_sfb : _GEN_62 ? _slots_17_io_out_uop_is_sfb : _GEN_61 ? _slots_16_io_out_uop_is_sfb : _slots_15_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_63 ? _slots_18_io_out_uop_br_mask : _GEN_62 ? _slots_17_io_out_uop_br_mask : _GEN_61 ? _slots_16_io_out_uop_br_mask : _slots_15_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_63 ? _slots_18_io_out_uop_br_tag : _GEN_62 ? _slots_17_io_out_uop_br_tag : _GEN_61 ? _slots_16_io_out_uop_br_tag : _slots_15_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_63 ? _slots_18_io_out_uop_ftq_idx : _GEN_62 ? _slots_17_io_out_uop_ftq_idx : _GEN_61 ? _slots_16_io_out_uop_ftq_idx : _slots_15_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_63 ? _slots_18_io_out_uop_edge_inst : _GEN_62 ? _slots_17_io_out_uop_edge_inst : _GEN_61 ? _slots_16_io_out_uop_edge_inst : _slots_15_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_63 ? _slots_18_io_out_uop_pc_lob : _GEN_62 ? _slots_17_io_out_uop_pc_lob : _GEN_61 ? _slots_16_io_out_uop_pc_lob : _slots_15_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_63 ? _slots_18_io_out_uop_taken : _GEN_62 ? _slots_17_io_out_uop_taken : _GEN_61 ? _slots_16_io_out_uop_taken : _slots_15_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_63 ? _slots_18_io_out_uop_imm_packed : _GEN_62 ? _slots_17_io_out_uop_imm_packed : _GEN_61 ? _slots_16_io_out_uop_imm_packed : _slots_15_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_63 ? _slots_18_io_out_uop_csr_addr : _GEN_62 ? _slots_17_io_out_uop_csr_addr : _GEN_61 ? _slots_16_io_out_uop_csr_addr : _slots_15_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_63 ? _slots_18_io_out_uop_rob_idx : _GEN_62 ? _slots_17_io_out_uop_rob_idx : _GEN_61 ? _slots_16_io_out_uop_rob_idx : _slots_15_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_63 ? _slots_18_io_out_uop_ldq_idx : _GEN_62 ? _slots_17_io_out_uop_ldq_idx : _GEN_61 ? _slots_16_io_out_uop_ldq_idx : _slots_15_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_63 ? _slots_18_io_out_uop_stq_idx : _GEN_62 ? _slots_17_io_out_uop_stq_idx : _GEN_61 ? _slots_16_io_out_uop_stq_idx : _slots_15_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_63 ? _slots_18_io_out_uop_rxq_idx : _GEN_62 ? _slots_17_io_out_uop_rxq_idx : _GEN_61 ? _slots_16_io_out_uop_rxq_idx : _slots_15_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_63 ? _slots_18_io_out_uop_pdst : _GEN_62 ? _slots_17_io_out_uop_pdst : _GEN_61 ? _slots_16_io_out_uop_pdst : _slots_15_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_63 ? _slots_18_io_out_uop_prs1 : _GEN_62 ? _slots_17_io_out_uop_prs1 : _GEN_61 ? _slots_16_io_out_uop_prs1 : _slots_15_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_63 ? _slots_18_io_out_uop_prs2 : _GEN_62 ? _slots_17_io_out_uop_prs2 : _GEN_61 ? _slots_16_io_out_uop_prs2 : _slots_15_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_63 ? _slots_18_io_out_uop_prs3 : _GEN_62 ? _slots_17_io_out_uop_prs3 : _GEN_61 ? _slots_16_io_out_uop_prs3 : _slots_15_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_63 ? _slots_18_io_out_uop_ppred : _GEN_62 ? _slots_17_io_out_uop_ppred : _GEN_61 ? _slots_16_io_out_uop_ppred : _slots_15_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_63 ? _slots_18_io_out_uop_prs1_busy : _GEN_62 ? _slots_17_io_out_uop_prs1_busy : _GEN_61 ? _slots_16_io_out_uop_prs1_busy : _slots_15_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_63 ? _slots_18_io_out_uop_prs2_busy : _GEN_62 ? _slots_17_io_out_uop_prs2_busy : _GEN_61 ? _slots_16_io_out_uop_prs2_busy : _slots_15_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_63 ? _slots_18_io_out_uop_prs3_busy : _GEN_62 ? _slots_17_io_out_uop_prs3_busy : _GEN_61 ? _slots_16_io_out_uop_prs3_busy : _slots_15_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_63 ? _slots_18_io_out_uop_ppred_busy : _GEN_62 ? _slots_17_io_out_uop_ppred_busy : _GEN_61 ? _slots_16_io_out_uop_ppred_busy : _slots_15_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_63 ? _slots_18_io_out_uop_stale_pdst : _GEN_62 ? _slots_17_io_out_uop_stale_pdst : _GEN_61 ? _slots_16_io_out_uop_stale_pdst : _slots_15_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_63 ? _slots_18_io_out_uop_exception : _GEN_62 ? _slots_17_io_out_uop_exception : _GEN_61 ? _slots_16_io_out_uop_exception : _slots_15_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_63 ? _slots_18_io_out_uop_exc_cause : _GEN_62 ? _slots_17_io_out_uop_exc_cause : _GEN_61 ? _slots_16_io_out_uop_exc_cause : _slots_15_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_63 ? _slots_18_io_out_uop_bypassable : _GEN_62 ? _slots_17_io_out_uop_bypassable : _GEN_61 ? _slots_16_io_out_uop_bypassable : _slots_15_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_63 ? _slots_18_io_out_uop_mem_cmd : _GEN_62 ? _slots_17_io_out_uop_mem_cmd : _GEN_61 ? _slots_16_io_out_uop_mem_cmd : _slots_15_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_63 ? _slots_18_io_out_uop_mem_size : _GEN_62 ? _slots_17_io_out_uop_mem_size : _GEN_61 ? _slots_16_io_out_uop_mem_size : _slots_15_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_63 ? _slots_18_io_out_uop_mem_signed : _GEN_62 ? _slots_17_io_out_uop_mem_signed : _GEN_61 ? _slots_16_io_out_uop_mem_signed : _slots_15_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_63 ? _slots_18_io_out_uop_is_fence : _GEN_62 ? _slots_17_io_out_uop_is_fence : _GEN_61 ? _slots_16_io_out_uop_is_fence : _slots_15_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_63 ? _slots_18_io_out_uop_is_fencei : _GEN_62 ? _slots_17_io_out_uop_is_fencei : _GEN_61 ? _slots_16_io_out_uop_is_fencei : _slots_15_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_63 ? _slots_18_io_out_uop_is_amo : _GEN_62 ? _slots_17_io_out_uop_is_amo : _GEN_61 ? _slots_16_io_out_uop_is_amo : _slots_15_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_63 ? _slots_18_io_out_uop_uses_ldq : _GEN_62 ? _slots_17_io_out_uop_uses_ldq : _GEN_61 ? _slots_16_io_out_uop_uses_ldq : _slots_15_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_63 ? _slots_18_io_out_uop_uses_stq : _GEN_62 ? _slots_17_io_out_uop_uses_stq : _GEN_61 ? _slots_16_io_out_uop_uses_stq : _slots_15_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_63 ? _slots_18_io_out_uop_is_sys_pc2epc : _GEN_62 ? _slots_17_io_out_uop_is_sys_pc2epc : _GEN_61 ? _slots_16_io_out_uop_is_sys_pc2epc : _slots_15_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_63 ? _slots_18_io_out_uop_is_unique : _GEN_62 ? _slots_17_io_out_uop_is_unique : _GEN_61 ? _slots_16_io_out_uop_is_unique : _slots_15_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_63 ? _slots_18_io_out_uop_flush_on_commit : _GEN_62 ? _slots_17_io_out_uop_flush_on_commit : _GEN_61 ? _slots_16_io_out_uop_flush_on_commit : _slots_15_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_63 ? _slots_18_io_out_uop_ldst_is_rs1 : _GEN_62 ? _slots_17_io_out_uop_ldst_is_rs1 : _GEN_61 ? _slots_16_io_out_uop_ldst_is_rs1 : _slots_15_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_63 ? _slots_18_io_out_uop_ldst : _GEN_62 ? _slots_17_io_out_uop_ldst : _GEN_61 ? _slots_16_io_out_uop_ldst : _slots_15_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_63 ? _slots_18_io_out_uop_lrs1 : _GEN_62 ? _slots_17_io_out_uop_lrs1 : _GEN_61 ? _slots_16_io_out_uop_lrs1 : _slots_15_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_63 ? _slots_18_io_out_uop_lrs2 : _GEN_62 ? _slots_17_io_out_uop_lrs2 : _GEN_61 ? _slots_16_io_out_uop_lrs2 : _slots_15_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_63 ? _slots_18_io_out_uop_lrs3 : _GEN_62 ? _slots_17_io_out_uop_lrs3 : _GEN_61 ? _slots_16_io_out_uop_lrs3 : _slots_15_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_63 ? _slots_18_io_out_uop_ldst_val : _GEN_62 ? _slots_17_io_out_uop_ldst_val : _GEN_61 ? _slots_16_io_out_uop_ldst_val : _slots_15_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_63 ? _slots_18_io_out_uop_dst_rtype : _GEN_62 ? _slots_17_io_out_uop_dst_rtype : _GEN_61 ? _slots_16_io_out_uop_dst_rtype : _slots_15_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_63 ? _slots_18_io_out_uop_lrs1_rtype : _GEN_62 ? _slots_17_io_out_uop_lrs1_rtype : _GEN_61 ? _slots_16_io_out_uop_lrs1_rtype : _slots_15_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_63 ? _slots_18_io_out_uop_lrs2_rtype : _GEN_62 ? _slots_17_io_out_uop_lrs2_rtype : _GEN_61 ? _slots_16_io_out_uop_lrs2_rtype : _slots_15_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_63 ? _slots_18_io_out_uop_frs3_en : _GEN_62 ? _slots_17_io_out_uop_frs3_en : _GEN_61 ? _slots_16_io_out_uop_frs3_en : _slots_15_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_63 ? _slots_18_io_out_uop_fp_val : _GEN_62 ? _slots_17_io_out_uop_fp_val : _GEN_61 ? _slots_16_io_out_uop_fp_val : _slots_15_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_63 ? _slots_18_io_out_uop_fp_single : _GEN_62 ? _slots_17_io_out_uop_fp_single : _GEN_61 ? _slots_16_io_out_uop_fp_single : _slots_15_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_63 ? _slots_18_io_out_uop_xcpt_pf_if : _GEN_62 ? _slots_17_io_out_uop_xcpt_pf_if : _GEN_61 ? _slots_16_io_out_uop_xcpt_pf_if : _slots_15_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_63 ? _slots_18_io_out_uop_xcpt_ae_if : _GEN_62 ? _slots_17_io_out_uop_xcpt_ae_if : _GEN_61 ? _slots_16_io_out_uop_xcpt_ae_if : _slots_15_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_63 ? _slots_18_io_out_uop_xcpt_ma_if : _GEN_62 ? _slots_17_io_out_uop_xcpt_ma_if : _GEN_61 ? _slots_16_io_out_uop_xcpt_ma_if : _slots_15_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_63 ? _slots_18_io_out_uop_bp_debug_if : _GEN_62 ? _slots_17_io_out_uop_bp_debug_if : _GEN_61 ? _slots_16_io_out_uop_bp_debug_if : _slots_15_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_63 ? _slots_18_io_out_uop_bp_xcpt_if : _GEN_62 ? _slots_17_io_out_uop_bp_xcpt_if : _GEN_61 ? _slots_16_io_out_uop_bp_xcpt_if : _slots_15_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_63 ? _slots_18_io_out_uop_debug_fsrc : _GEN_62 ? _slots_17_io_out_uop_debug_fsrc : _GEN_61 ? _slots_16_io_out_uop_debug_fsrc : _slots_15_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_63 ? _slots_18_io_out_uop_debug_tsrc : _GEN_62 ? _slots_17_io_out_uop_debug_tsrc : _GEN_61 ? _slots_16_io_out_uop_debug_tsrc : _slots_15_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_14_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_14_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_14_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_14_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_14_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_14_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_14_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_14_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_14_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_14_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_14_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_14_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_14_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_14_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_14_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_14_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_14_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_14_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_14_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_14_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_14_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_14_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_14_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_14_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_14_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_14_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_14_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_14_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_14_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_14_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_14_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_14_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_14_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_14_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_14_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_14_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_14_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_14_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_14_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_14_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_14_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_14_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_14_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_14_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_14_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_14_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_14_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_14_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_14_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_14_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_14_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_14_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_14_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_14_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_14_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_14_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_14_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_14_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_14_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_14_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_14_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_14_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_14_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_14_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_14_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_14_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_14_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_14_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_14_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_14_io_uop_uopc),
    .io_uop_inst                    (_slots_14_io_uop_inst),
    .io_uop_debug_inst              (_slots_14_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_14_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_14_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_14_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_14_io_uop_fu_code),
    .io_uop_iw_state                (_slots_14_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_14_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_14_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_14_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_14_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_14_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_14_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_14_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_14_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_14_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_14_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_14_io_uop_pc_lob),
    .io_uop_taken                   (_slots_14_io_uop_taken),
    .io_uop_imm_packed              (_slots_14_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_14_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_14_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_14_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_14_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_14_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_14_io_uop_pdst),
    .io_uop_prs1                    (_slots_14_io_uop_prs1),
    .io_uop_prs2                    (_slots_14_io_uop_prs2),
    .io_uop_prs3                    (_slots_14_io_uop_prs3),
    .io_uop_ppred                   (_slots_14_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_14_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_14_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_14_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_14_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_14_io_uop_stale_pdst),
    .io_uop_exception               (_slots_14_io_uop_exception),
    .io_uop_exc_cause               (_slots_14_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_14_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_14_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_14_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_14_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_14_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_14_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_14_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_14_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_14_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_14_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_14_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_14_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_14_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_14_io_uop_ldst),
    .io_uop_lrs1                    (_slots_14_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_14_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_14_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_14_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_14_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_14_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_14_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_14_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_14_io_uop_fp_val),
    .io_uop_fp_single               (_slots_14_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_14_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_14_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_14_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_14_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_14_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_14_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_14_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_15 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_15_io_valid),
    .io_will_be_valid               (_slots_15_io_will_be_valid),
    .io_request                     (_slots_15_io_request),
    .io_grant                       (issue_slots_15_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_14),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_15_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_66 ? _slots_19_io_out_uop_uopc : _GEN_65 ? _slots_18_io_out_uop_uopc : _GEN_64 ? _slots_17_io_out_uop_uopc : _slots_16_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_66 ? _slots_19_io_out_uop_inst : _GEN_65 ? _slots_18_io_out_uop_inst : _GEN_64 ? _slots_17_io_out_uop_inst : _slots_16_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_66 ? _slots_19_io_out_uop_debug_inst : _GEN_65 ? _slots_18_io_out_uop_debug_inst : _GEN_64 ? _slots_17_io_out_uop_debug_inst : _slots_16_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_66 ? _slots_19_io_out_uop_is_rvc : _GEN_65 ? _slots_18_io_out_uop_is_rvc : _GEN_64 ? _slots_17_io_out_uop_is_rvc : _slots_16_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_66 ? _slots_19_io_out_uop_debug_pc : _GEN_65 ? _slots_18_io_out_uop_debug_pc : _GEN_64 ? _slots_17_io_out_uop_debug_pc : _slots_16_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_66 ? _slots_19_io_out_uop_iq_type : _GEN_65 ? _slots_18_io_out_uop_iq_type : _GEN_64 ? _slots_17_io_out_uop_iq_type : _slots_16_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_66 ? _slots_19_io_out_uop_fu_code : _GEN_65 ? _slots_18_io_out_uop_fu_code : _GEN_64 ? _slots_17_io_out_uop_fu_code : _slots_16_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_66 ? _slots_19_io_out_uop_iw_state : _GEN_65 ? _slots_18_io_out_uop_iw_state : _GEN_64 ? _slots_17_io_out_uop_iw_state : _slots_16_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_66 ? _slots_19_io_out_uop_iw_p1_poisoned : _GEN_65 ? _slots_18_io_out_uop_iw_p1_poisoned : _GEN_64 ? _slots_17_io_out_uop_iw_p1_poisoned : _slots_16_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_66 ? _slots_19_io_out_uop_iw_p2_poisoned : _GEN_65 ? _slots_18_io_out_uop_iw_p2_poisoned : _GEN_64 ? _slots_17_io_out_uop_iw_p2_poisoned : _slots_16_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_66 ? _slots_19_io_out_uop_is_br : _GEN_65 ? _slots_18_io_out_uop_is_br : _GEN_64 ? _slots_17_io_out_uop_is_br : _slots_16_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_66 ? _slots_19_io_out_uop_is_jalr : _GEN_65 ? _slots_18_io_out_uop_is_jalr : _GEN_64 ? _slots_17_io_out_uop_is_jalr : _slots_16_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_66 ? _slots_19_io_out_uop_is_jal : _GEN_65 ? _slots_18_io_out_uop_is_jal : _GEN_64 ? _slots_17_io_out_uop_is_jal : _slots_16_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_66 ? _slots_19_io_out_uop_is_sfb : _GEN_65 ? _slots_18_io_out_uop_is_sfb : _GEN_64 ? _slots_17_io_out_uop_is_sfb : _slots_16_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_66 ? _slots_19_io_out_uop_br_mask : _GEN_65 ? _slots_18_io_out_uop_br_mask : _GEN_64 ? _slots_17_io_out_uop_br_mask : _slots_16_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_66 ? _slots_19_io_out_uop_br_tag : _GEN_65 ? _slots_18_io_out_uop_br_tag : _GEN_64 ? _slots_17_io_out_uop_br_tag : _slots_16_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_66 ? _slots_19_io_out_uop_ftq_idx : _GEN_65 ? _slots_18_io_out_uop_ftq_idx : _GEN_64 ? _slots_17_io_out_uop_ftq_idx : _slots_16_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_66 ? _slots_19_io_out_uop_edge_inst : _GEN_65 ? _slots_18_io_out_uop_edge_inst : _GEN_64 ? _slots_17_io_out_uop_edge_inst : _slots_16_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_66 ? _slots_19_io_out_uop_pc_lob : _GEN_65 ? _slots_18_io_out_uop_pc_lob : _GEN_64 ? _slots_17_io_out_uop_pc_lob : _slots_16_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_66 ? _slots_19_io_out_uop_taken : _GEN_65 ? _slots_18_io_out_uop_taken : _GEN_64 ? _slots_17_io_out_uop_taken : _slots_16_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_66 ? _slots_19_io_out_uop_imm_packed : _GEN_65 ? _slots_18_io_out_uop_imm_packed : _GEN_64 ? _slots_17_io_out_uop_imm_packed : _slots_16_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_66 ? _slots_19_io_out_uop_csr_addr : _GEN_65 ? _slots_18_io_out_uop_csr_addr : _GEN_64 ? _slots_17_io_out_uop_csr_addr : _slots_16_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_66 ? _slots_19_io_out_uop_rob_idx : _GEN_65 ? _slots_18_io_out_uop_rob_idx : _GEN_64 ? _slots_17_io_out_uop_rob_idx : _slots_16_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_66 ? _slots_19_io_out_uop_ldq_idx : _GEN_65 ? _slots_18_io_out_uop_ldq_idx : _GEN_64 ? _slots_17_io_out_uop_ldq_idx : _slots_16_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_66 ? _slots_19_io_out_uop_stq_idx : _GEN_65 ? _slots_18_io_out_uop_stq_idx : _GEN_64 ? _slots_17_io_out_uop_stq_idx : _slots_16_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_66 ? _slots_19_io_out_uop_rxq_idx : _GEN_65 ? _slots_18_io_out_uop_rxq_idx : _GEN_64 ? _slots_17_io_out_uop_rxq_idx : _slots_16_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_66 ? _slots_19_io_out_uop_pdst : _GEN_65 ? _slots_18_io_out_uop_pdst : _GEN_64 ? _slots_17_io_out_uop_pdst : _slots_16_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_66 ? _slots_19_io_out_uop_prs1 : _GEN_65 ? _slots_18_io_out_uop_prs1 : _GEN_64 ? _slots_17_io_out_uop_prs1 : _slots_16_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_66 ? _slots_19_io_out_uop_prs2 : _GEN_65 ? _slots_18_io_out_uop_prs2 : _GEN_64 ? _slots_17_io_out_uop_prs2 : _slots_16_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_66 ? _slots_19_io_out_uop_prs3 : _GEN_65 ? _slots_18_io_out_uop_prs3 : _GEN_64 ? _slots_17_io_out_uop_prs3 : _slots_16_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_66 ? _slots_19_io_out_uop_ppred : _GEN_65 ? _slots_18_io_out_uop_ppred : _GEN_64 ? _slots_17_io_out_uop_ppred : _slots_16_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_66 ? _slots_19_io_out_uop_prs1_busy : _GEN_65 ? _slots_18_io_out_uop_prs1_busy : _GEN_64 ? _slots_17_io_out_uop_prs1_busy : _slots_16_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_66 ? _slots_19_io_out_uop_prs2_busy : _GEN_65 ? _slots_18_io_out_uop_prs2_busy : _GEN_64 ? _slots_17_io_out_uop_prs2_busy : _slots_16_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_66 ? _slots_19_io_out_uop_prs3_busy : _GEN_65 ? _slots_18_io_out_uop_prs3_busy : _GEN_64 ? _slots_17_io_out_uop_prs3_busy : _slots_16_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_66 ? _slots_19_io_out_uop_ppred_busy : _GEN_65 ? _slots_18_io_out_uop_ppred_busy : _GEN_64 ? _slots_17_io_out_uop_ppred_busy : _slots_16_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_66 ? _slots_19_io_out_uop_stale_pdst : _GEN_65 ? _slots_18_io_out_uop_stale_pdst : _GEN_64 ? _slots_17_io_out_uop_stale_pdst : _slots_16_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_66 ? _slots_19_io_out_uop_exception : _GEN_65 ? _slots_18_io_out_uop_exception : _GEN_64 ? _slots_17_io_out_uop_exception : _slots_16_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_66 ? _slots_19_io_out_uop_exc_cause : _GEN_65 ? _slots_18_io_out_uop_exc_cause : _GEN_64 ? _slots_17_io_out_uop_exc_cause : _slots_16_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_66 ? _slots_19_io_out_uop_bypassable : _GEN_65 ? _slots_18_io_out_uop_bypassable : _GEN_64 ? _slots_17_io_out_uop_bypassable : _slots_16_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_66 ? _slots_19_io_out_uop_mem_cmd : _GEN_65 ? _slots_18_io_out_uop_mem_cmd : _GEN_64 ? _slots_17_io_out_uop_mem_cmd : _slots_16_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_66 ? _slots_19_io_out_uop_mem_size : _GEN_65 ? _slots_18_io_out_uop_mem_size : _GEN_64 ? _slots_17_io_out_uop_mem_size : _slots_16_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_66 ? _slots_19_io_out_uop_mem_signed : _GEN_65 ? _slots_18_io_out_uop_mem_signed : _GEN_64 ? _slots_17_io_out_uop_mem_signed : _slots_16_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_66 ? _slots_19_io_out_uop_is_fence : _GEN_65 ? _slots_18_io_out_uop_is_fence : _GEN_64 ? _slots_17_io_out_uop_is_fence : _slots_16_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_66 ? _slots_19_io_out_uop_is_fencei : _GEN_65 ? _slots_18_io_out_uop_is_fencei : _GEN_64 ? _slots_17_io_out_uop_is_fencei : _slots_16_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_66 ? _slots_19_io_out_uop_is_amo : _GEN_65 ? _slots_18_io_out_uop_is_amo : _GEN_64 ? _slots_17_io_out_uop_is_amo : _slots_16_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_66 ? _slots_19_io_out_uop_uses_ldq : _GEN_65 ? _slots_18_io_out_uop_uses_ldq : _GEN_64 ? _slots_17_io_out_uop_uses_ldq : _slots_16_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_66 ? _slots_19_io_out_uop_uses_stq : _GEN_65 ? _slots_18_io_out_uop_uses_stq : _GEN_64 ? _slots_17_io_out_uop_uses_stq : _slots_16_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_66 ? _slots_19_io_out_uop_is_sys_pc2epc : _GEN_65 ? _slots_18_io_out_uop_is_sys_pc2epc : _GEN_64 ? _slots_17_io_out_uop_is_sys_pc2epc : _slots_16_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_66 ? _slots_19_io_out_uop_is_unique : _GEN_65 ? _slots_18_io_out_uop_is_unique : _GEN_64 ? _slots_17_io_out_uop_is_unique : _slots_16_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_66 ? _slots_19_io_out_uop_flush_on_commit : _GEN_65 ? _slots_18_io_out_uop_flush_on_commit : _GEN_64 ? _slots_17_io_out_uop_flush_on_commit : _slots_16_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_66 ? _slots_19_io_out_uop_ldst_is_rs1 : _GEN_65 ? _slots_18_io_out_uop_ldst_is_rs1 : _GEN_64 ? _slots_17_io_out_uop_ldst_is_rs1 : _slots_16_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_66 ? _slots_19_io_out_uop_ldst : _GEN_65 ? _slots_18_io_out_uop_ldst : _GEN_64 ? _slots_17_io_out_uop_ldst : _slots_16_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_66 ? _slots_19_io_out_uop_lrs1 : _GEN_65 ? _slots_18_io_out_uop_lrs1 : _GEN_64 ? _slots_17_io_out_uop_lrs1 : _slots_16_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_66 ? _slots_19_io_out_uop_lrs2 : _GEN_65 ? _slots_18_io_out_uop_lrs2 : _GEN_64 ? _slots_17_io_out_uop_lrs2 : _slots_16_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_66 ? _slots_19_io_out_uop_lrs3 : _GEN_65 ? _slots_18_io_out_uop_lrs3 : _GEN_64 ? _slots_17_io_out_uop_lrs3 : _slots_16_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_66 ? _slots_19_io_out_uop_ldst_val : _GEN_65 ? _slots_18_io_out_uop_ldst_val : _GEN_64 ? _slots_17_io_out_uop_ldst_val : _slots_16_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_66 ? _slots_19_io_out_uop_dst_rtype : _GEN_65 ? _slots_18_io_out_uop_dst_rtype : _GEN_64 ? _slots_17_io_out_uop_dst_rtype : _slots_16_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_66 ? _slots_19_io_out_uop_lrs1_rtype : _GEN_65 ? _slots_18_io_out_uop_lrs1_rtype : _GEN_64 ? _slots_17_io_out_uop_lrs1_rtype : _slots_16_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_66 ? _slots_19_io_out_uop_lrs2_rtype : _GEN_65 ? _slots_18_io_out_uop_lrs2_rtype : _GEN_64 ? _slots_17_io_out_uop_lrs2_rtype : _slots_16_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_66 ? _slots_19_io_out_uop_frs3_en : _GEN_65 ? _slots_18_io_out_uop_frs3_en : _GEN_64 ? _slots_17_io_out_uop_frs3_en : _slots_16_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_66 ? _slots_19_io_out_uop_fp_val : _GEN_65 ? _slots_18_io_out_uop_fp_val : _GEN_64 ? _slots_17_io_out_uop_fp_val : _slots_16_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_66 ? _slots_19_io_out_uop_fp_single : _GEN_65 ? _slots_18_io_out_uop_fp_single : _GEN_64 ? _slots_17_io_out_uop_fp_single : _slots_16_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_66 ? _slots_19_io_out_uop_xcpt_pf_if : _GEN_65 ? _slots_18_io_out_uop_xcpt_pf_if : _GEN_64 ? _slots_17_io_out_uop_xcpt_pf_if : _slots_16_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_66 ? _slots_19_io_out_uop_xcpt_ae_if : _GEN_65 ? _slots_18_io_out_uop_xcpt_ae_if : _GEN_64 ? _slots_17_io_out_uop_xcpt_ae_if : _slots_16_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_66 ? _slots_19_io_out_uop_xcpt_ma_if : _GEN_65 ? _slots_18_io_out_uop_xcpt_ma_if : _GEN_64 ? _slots_17_io_out_uop_xcpt_ma_if : _slots_16_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_66 ? _slots_19_io_out_uop_bp_debug_if : _GEN_65 ? _slots_18_io_out_uop_bp_debug_if : _GEN_64 ? _slots_17_io_out_uop_bp_debug_if : _slots_16_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_66 ? _slots_19_io_out_uop_bp_xcpt_if : _GEN_65 ? _slots_18_io_out_uop_bp_xcpt_if : _GEN_64 ? _slots_17_io_out_uop_bp_xcpt_if : _slots_16_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_66 ? _slots_19_io_out_uop_debug_fsrc : _GEN_65 ? _slots_18_io_out_uop_debug_fsrc : _GEN_64 ? _slots_17_io_out_uop_debug_fsrc : _slots_16_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_66 ? _slots_19_io_out_uop_debug_tsrc : _GEN_65 ? _slots_18_io_out_uop_debug_tsrc : _GEN_64 ? _slots_17_io_out_uop_debug_tsrc : _slots_16_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_15_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_15_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_15_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_15_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_15_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_15_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_15_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_15_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_15_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_15_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_15_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_15_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_15_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_15_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_15_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_15_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_15_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_15_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_15_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_15_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_15_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_15_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_15_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_15_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_15_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_15_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_15_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_15_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_15_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_15_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_15_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_15_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_15_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_15_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_15_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_15_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_15_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_15_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_15_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_15_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_15_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_15_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_15_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_15_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_15_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_15_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_15_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_15_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_15_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_15_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_15_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_15_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_15_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_15_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_15_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_15_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_15_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_15_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_15_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_15_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_15_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_15_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_15_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_15_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_15_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_15_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_15_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_15_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_15_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_15_io_uop_uopc),
    .io_uop_inst                    (_slots_15_io_uop_inst),
    .io_uop_debug_inst              (_slots_15_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_15_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_15_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_15_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_15_io_uop_fu_code),
    .io_uop_iw_state                (_slots_15_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_15_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_15_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_15_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_15_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_15_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_15_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_15_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_15_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_15_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_15_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_15_io_uop_pc_lob),
    .io_uop_taken                   (_slots_15_io_uop_taken),
    .io_uop_imm_packed              (_slots_15_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_15_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_15_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_15_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_15_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_15_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_15_io_uop_pdst),
    .io_uop_prs1                    (_slots_15_io_uop_prs1),
    .io_uop_prs2                    (_slots_15_io_uop_prs2),
    .io_uop_prs3                    (_slots_15_io_uop_prs3),
    .io_uop_ppred                   (_slots_15_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_15_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_15_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_15_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_15_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_15_io_uop_stale_pdst),
    .io_uop_exception               (_slots_15_io_uop_exception),
    .io_uop_exc_cause               (_slots_15_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_15_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_15_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_15_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_15_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_15_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_15_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_15_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_15_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_15_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_15_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_15_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_15_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_15_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_15_io_uop_ldst),
    .io_uop_lrs1                    (_slots_15_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_15_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_15_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_15_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_15_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_15_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_15_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_15_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_15_io_uop_fp_val),
    .io_uop_fp_single               (_slots_15_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_15_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_15_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_15_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_15_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_15_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_15_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_15_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_16 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_16_io_valid),
    .io_will_be_valid               (_slots_16_io_will_be_valid),
    .io_request                     (_slots_16_io_request),
    .io_grant                       (issue_slots_16_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_15),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_16_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_69 ? _slots_20_io_out_uop_uopc : _GEN_68 ? _slots_19_io_out_uop_uopc : _GEN_67 ? _slots_18_io_out_uop_uopc : _slots_17_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_69 ? _slots_20_io_out_uop_inst : _GEN_68 ? _slots_19_io_out_uop_inst : _GEN_67 ? _slots_18_io_out_uop_inst : _slots_17_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_69 ? _slots_20_io_out_uop_debug_inst : _GEN_68 ? _slots_19_io_out_uop_debug_inst : _GEN_67 ? _slots_18_io_out_uop_debug_inst : _slots_17_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_69 ? _slots_20_io_out_uop_is_rvc : _GEN_68 ? _slots_19_io_out_uop_is_rvc : _GEN_67 ? _slots_18_io_out_uop_is_rvc : _slots_17_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_69 ? _slots_20_io_out_uop_debug_pc : _GEN_68 ? _slots_19_io_out_uop_debug_pc : _GEN_67 ? _slots_18_io_out_uop_debug_pc : _slots_17_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_69 ? _slots_20_io_out_uop_iq_type : _GEN_68 ? _slots_19_io_out_uop_iq_type : _GEN_67 ? _slots_18_io_out_uop_iq_type : _slots_17_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_69 ? _slots_20_io_out_uop_fu_code : _GEN_68 ? _slots_19_io_out_uop_fu_code : _GEN_67 ? _slots_18_io_out_uop_fu_code : _slots_17_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_69 ? _slots_20_io_out_uop_iw_state : _GEN_68 ? _slots_19_io_out_uop_iw_state : _GEN_67 ? _slots_18_io_out_uop_iw_state : _slots_17_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_69 ? _slots_20_io_out_uop_iw_p1_poisoned : _GEN_68 ? _slots_19_io_out_uop_iw_p1_poisoned : _GEN_67 ? _slots_18_io_out_uop_iw_p1_poisoned : _slots_17_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_69 ? _slots_20_io_out_uop_iw_p2_poisoned : _GEN_68 ? _slots_19_io_out_uop_iw_p2_poisoned : _GEN_67 ? _slots_18_io_out_uop_iw_p2_poisoned : _slots_17_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_69 ? _slots_20_io_out_uop_is_br : _GEN_68 ? _slots_19_io_out_uop_is_br : _GEN_67 ? _slots_18_io_out_uop_is_br : _slots_17_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_69 ? _slots_20_io_out_uop_is_jalr : _GEN_68 ? _slots_19_io_out_uop_is_jalr : _GEN_67 ? _slots_18_io_out_uop_is_jalr : _slots_17_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_69 ? _slots_20_io_out_uop_is_jal : _GEN_68 ? _slots_19_io_out_uop_is_jal : _GEN_67 ? _slots_18_io_out_uop_is_jal : _slots_17_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_69 ? _slots_20_io_out_uop_is_sfb : _GEN_68 ? _slots_19_io_out_uop_is_sfb : _GEN_67 ? _slots_18_io_out_uop_is_sfb : _slots_17_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_69 ? _slots_20_io_out_uop_br_mask : _GEN_68 ? _slots_19_io_out_uop_br_mask : _GEN_67 ? _slots_18_io_out_uop_br_mask : _slots_17_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_69 ? _slots_20_io_out_uop_br_tag : _GEN_68 ? _slots_19_io_out_uop_br_tag : _GEN_67 ? _slots_18_io_out_uop_br_tag : _slots_17_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_69 ? _slots_20_io_out_uop_ftq_idx : _GEN_68 ? _slots_19_io_out_uop_ftq_idx : _GEN_67 ? _slots_18_io_out_uop_ftq_idx : _slots_17_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_69 ? _slots_20_io_out_uop_edge_inst : _GEN_68 ? _slots_19_io_out_uop_edge_inst : _GEN_67 ? _slots_18_io_out_uop_edge_inst : _slots_17_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_69 ? _slots_20_io_out_uop_pc_lob : _GEN_68 ? _slots_19_io_out_uop_pc_lob : _GEN_67 ? _slots_18_io_out_uop_pc_lob : _slots_17_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_69 ? _slots_20_io_out_uop_taken : _GEN_68 ? _slots_19_io_out_uop_taken : _GEN_67 ? _slots_18_io_out_uop_taken : _slots_17_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_69 ? _slots_20_io_out_uop_imm_packed : _GEN_68 ? _slots_19_io_out_uop_imm_packed : _GEN_67 ? _slots_18_io_out_uop_imm_packed : _slots_17_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_69 ? _slots_20_io_out_uop_csr_addr : _GEN_68 ? _slots_19_io_out_uop_csr_addr : _GEN_67 ? _slots_18_io_out_uop_csr_addr : _slots_17_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_69 ? _slots_20_io_out_uop_rob_idx : _GEN_68 ? _slots_19_io_out_uop_rob_idx : _GEN_67 ? _slots_18_io_out_uop_rob_idx : _slots_17_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_69 ? _slots_20_io_out_uop_ldq_idx : _GEN_68 ? _slots_19_io_out_uop_ldq_idx : _GEN_67 ? _slots_18_io_out_uop_ldq_idx : _slots_17_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_69 ? _slots_20_io_out_uop_stq_idx : _GEN_68 ? _slots_19_io_out_uop_stq_idx : _GEN_67 ? _slots_18_io_out_uop_stq_idx : _slots_17_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_69 ? _slots_20_io_out_uop_rxq_idx : _GEN_68 ? _slots_19_io_out_uop_rxq_idx : _GEN_67 ? _slots_18_io_out_uop_rxq_idx : _slots_17_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_69 ? _slots_20_io_out_uop_pdst : _GEN_68 ? _slots_19_io_out_uop_pdst : _GEN_67 ? _slots_18_io_out_uop_pdst : _slots_17_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_69 ? _slots_20_io_out_uop_prs1 : _GEN_68 ? _slots_19_io_out_uop_prs1 : _GEN_67 ? _slots_18_io_out_uop_prs1 : _slots_17_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_69 ? _slots_20_io_out_uop_prs2 : _GEN_68 ? _slots_19_io_out_uop_prs2 : _GEN_67 ? _slots_18_io_out_uop_prs2 : _slots_17_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_69 ? _slots_20_io_out_uop_prs3 : _GEN_68 ? _slots_19_io_out_uop_prs3 : _GEN_67 ? _slots_18_io_out_uop_prs3 : _slots_17_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_69 ? _slots_20_io_out_uop_ppred : _GEN_68 ? _slots_19_io_out_uop_ppred : _GEN_67 ? _slots_18_io_out_uop_ppred : _slots_17_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_69 ? _slots_20_io_out_uop_prs1_busy : _GEN_68 ? _slots_19_io_out_uop_prs1_busy : _GEN_67 ? _slots_18_io_out_uop_prs1_busy : _slots_17_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_69 ? _slots_20_io_out_uop_prs2_busy : _GEN_68 ? _slots_19_io_out_uop_prs2_busy : _GEN_67 ? _slots_18_io_out_uop_prs2_busy : _slots_17_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_69 ? _slots_20_io_out_uop_prs3_busy : _GEN_68 ? _slots_19_io_out_uop_prs3_busy : _GEN_67 ? _slots_18_io_out_uop_prs3_busy : _slots_17_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_69 ? _slots_20_io_out_uop_ppred_busy : _GEN_68 ? _slots_19_io_out_uop_ppred_busy : _GEN_67 ? _slots_18_io_out_uop_ppred_busy : _slots_17_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_69 ? _slots_20_io_out_uop_stale_pdst : _GEN_68 ? _slots_19_io_out_uop_stale_pdst : _GEN_67 ? _slots_18_io_out_uop_stale_pdst : _slots_17_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_69 ? _slots_20_io_out_uop_exception : _GEN_68 ? _slots_19_io_out_uop_exception : _GEN_67 ? _slots_18_io_out_uop_exception : _slots_17_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_69 ? _slots_20_io_out_uop_exc_cause : _GEN_68 ? _slots_19_io_out_uop_exc_cause : _GEN_67 ? _slots_18_io_out_uop_exc_cause : _slots_17_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_69 ? _slots_20_io_out_uop_bypassable : _GEN_68 ? _slots_19_io_out_uop_bypassable : _GEN_67 ? _slots_18_io_out_uop_bypassable : _slots_17_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_69 ? _slots_20_io_out_uop_mem_cmd : _GEN_68 ? _slots_19_io_out_uop_mem_cmd : _GEN_67 ? _slots_18_io_out_uop_mem_cmd : _slots_17_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_69 ? _slots_20_io_out_uop_mem_size : _GEN_68 ? _slots_19_io_out_uop_mem_size : _GEN_67 ? _slots_18_io_out_uop_mem_size : _slots_17_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_69 ? _slots_20_io_out_uop_mem_signed : _GEN_68 ? _slots_19_io_out_uop_mem_signed : _GEN_67 ? _slots_18_io_out_uop_mem_signed : _slots_17_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_69 ? _slots_20_io_out_uop_is_fence : _GEN_68 ? _slots_19_io_out_uop_is_fence : _GEN_67 ? _slots_18_io_out_uop_is_fence : _slots_17_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_69 ? _slots_20_io_out_uop_is_fencei : _GEN_68 ? _slots_19_io_out_uop_is_fencei : _GEN_67 ? _slots_18_io_out_uop_is_fencei : _slots_17_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_69 ? _slots_20_io_out_uop_is_amo : _GEN_68 ? _slots_19_io_out_uop_is_amo : _GEN_67 ? _slots_18_io_out_uop_is_amo : _slots_17_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_69 ? _slots_20_io_out_uop_uses_ldq : _GEN_68 ? _slots_19_io_out_uop_uses_ldq : _GEN_67 ? _slots_18_io_out_uop_uses_ldq : _slots_17_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_69 ? _slots_20_io_out_uop_uses_stq : _GEN_68 ? _slots_19_io_out_uop_uses_stq : _GEN_67 ? _slots_18_io_out_uop_uses_stq : _slots_17_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_69 ? _slots_20_io_out_uop_is_sys_pc2epc : _GEN_68 ? _slots_19_io_out_uop_is_sys_pc2epc : _GEN_67 ? _slots_18_io_out_uop_is_sys_pc2epc : _slots_17_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_69 ? _slots_20_io_out_uop_is_unique : _GEN_68 ? _slots_19_io_out_uop_is_unique : _GEN_67 ? _slots_18_io_out_uop_is_unique : _slots_17_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_69 ? _slots_20_io_out_uop_flush_on_commit : _GEN_68 ? _slots_19_io_out_uop_flush_on_commit : _GEN_67 ? _slots_18_io_out_uop_flush_on_commit : _slots_17_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_69 ? _slots_20_io_out_uop_ldst_is_rs1 : _GEN_68 ? _slots_19_io_out_uop_ldst_is_rs1 : _GEN_67 ? _slots_18_io_out_uop_ldst_is_rs1 : _slots_17_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_69 ? _slots_20_io_out_uop_ldst : _GEN_68 ? _slots_19_io_out_uop_ldst : _GEN_67 ? _slots_18_io_out_uop_ldst : _slots_17_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_69 ? _slots_20_io_out_uop_lrs1 : _GEN_68 ? _slots_19_io_out_uop_lrs1 : _GEN_67 ? _slots_18_io_out_uop_lrs1 : _slots_17_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_69 ? _slots_20_io_out_uop_lrs2 : _GEN_68 ? _slots_19_io_out_uop_lrs2 : _GEN_67 ? _slots_18_io_out_uop_lrs2 : _slots_17_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_69 ? _slots_20_io_out_uop_lrs3 : _GEN_68 ? _slots_19_io_out_uop_lrs3 : _GEN_67 ? _slots_18_io_out_uop_lrs3 : _slots_17_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_69 ? _slots_20_io_out_uop_ldst_val : _GEN_68 ? _slots_19_io_out_uop_ldst_val : _GEN_67 ? _slots_18_io_out_uop_ldst_val : _slots_17_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_69 ? _slots_20_io_out_uop_dst_rtype : _GEN_68 ? _slots_19_io_out_uop_dst_rtype : _GEN_67 ? _slots_18_io_out_uop_dst_rtype : _slots_17_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_69 ? _slots_20_io_out_uop_lrs1_rtype : _GEN_68 ? _slots_19_io_out_uop_lrs1_rtype : _GEN_67 ? _slots_18_io_out_uop_lrs1_rtype : _slots_17_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_69 ? _slots_20_io_out_uop_lrs2_rtype : _GEN_68 ? _slots_19_io_out_uop_lrs2_rtype : _GEN_67 ? _slots_18_io_out_uop_lrs2_rtype : _slots_17_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_69 ? _slots_20_io_out_uop_frs3_en : _GEN_68 ? _slots_19_io_out_uop_frs3_en : _GEN_67 ? _slots_18_io_out_uop_frs3_en : _slots_17_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_69 ? _slots_20_io_out_uop_fp_val : _GEN_68 ? _slots_19_io_out_uop_fp_val : _GEN_67 ? _slots_18_io_out_uop_fp_val : _slots_17_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_69 ? _slots_20_io_out_uop_fp_single : _GEN_68 ? _slots_19_io_out_uop_fp_single : _GEN_67 ? _slots_18_io_out_uop_fp_single : _slots_17_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_69 ? _slots_20_io_out_uop_xcpt_pf_if : _GEN_68 ? _slots_19_io_out_uop_xcpt_pf_if : _GEN_67 ? _slots_18_io_out_uop_xcpt_pf_if : _slots_17_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_69 ? _slots_20_io_out_uop_xcpt_ae_if : _GEN_68 ? _slots_19_io_out_uop_xcpt_ae_if : _GEN_67 ? _slots_18_io_out_uop_xcpt_ae_if : _slots_17_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_69 ? _slots_20_io_out_uop_xcpt_ma_if : _GEN_68 ? _slots_19_io_out_uop_xcpt_ma_if : _GEN_67 ? _slots_18_io_out_uop_xcpt_ma_if : _slots_17_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_69 ? _slots_20_io_out_uop_bp_debug_if : _GEN_68 ? _slots_19_io_out_uop_bp_debug_if : _GEN_67 ? _slots_18_io_out_uop_bp_debug_if : _slots_17_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_69 ? _slots_20_io_out_uop_bp_xcpt_if : _GEN_68 ? _slots_19_io_out_uop_bp_xcpt_if : _GEN_67 ? _slots_18_io_out_uop_bp_xcpt_if : _slots_17_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_69 ? _slots_20_io_out_uop_debug_fsrc : _GEN_68 ? _slots_19_io_out_uop_debug_fsrc : _GEN_67 ? _slots_18_io_out_uop_debug_fsrc : _slots_17_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_69 ? _slots_20_io_out_uop_debug_tsrc : _GEN_68 ? _slots_19_io_out_uop_debug_tsrc : _GEN_67 ? _slots_18_io_out_uop_debug_tsrc : _slots_17_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_16_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_16_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_16_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_16_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_16_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_16_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_16_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_16_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_16_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_16_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_16_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_16_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_16_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_16_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_16_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_16_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_16_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_16_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_16_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_16_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_16_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_16_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_16_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_16_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_16_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_16_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_16_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_16_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_16_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_16_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_16_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_16_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_16_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_16_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_16_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_16_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_16_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_16_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_16_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_16_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_16_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_16_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_16_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_16_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_16_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_16_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_16_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_16_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_16_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_16_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_16_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_16_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_16_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_16_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_16_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_16_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_16_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_16_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_16_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_16_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_16_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_16_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_16_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_16_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_16_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_16_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_16_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_16_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_16_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_16_io_uop_uopc),
    .io_uop_inst                    (_slots_16_io_uop_inst),
    .io_uop_debug_inst              (_slots_16_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_16_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_16_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_16_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_16_io_uop_fu_code),
    .io_uop_iw_state                (_slots_16_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_16_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_16_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_16_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_16_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_16_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_16_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_16_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_16_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_16_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_16_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_16_io_uop_pc_lob),
    .io_uop_taken                   (_slots_16_io_uop_taken),
    .io_uop_imm_packed              (_slots_16_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_16_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_16_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_16_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_16_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_16_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_16_io_uop_pdst),
    .io_uop_prs1                    (_slots_16_io_uop_prs1),
    .io_uop_prs2                    (_slots_16_io_uop_prs2),
    .io_uop_prs3                    (_slots_16_io_uop_prs3),
    .io_uop_ppred                   (_slots_16_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_16_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_16_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_16_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_16_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_16_io_uop_stale_pdst),
    .io_uop_exception               (_slots_16_io_uop_exception),
    .io_uop_exc_cause               (_slots_16_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_16_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_16_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_16_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_16_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_16_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_16_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_16_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_16_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_16_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_16_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_16_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_16_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_16_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_16_io_uop_ldst),
    .io_uop_lrs1                    (_slots_16_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_16_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_16_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_16_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_16_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_16_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_16_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_16_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_16_io_uop_fp_val),
    .io_uop_fp_single               (_slots_16_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_16_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_16_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_16_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_16_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_16_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_16_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_16_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_17 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_17_io_valid),
    .io_will_be_valid               (_slots_17_io_will_be_valid),
    .io_request                     (_slots_17_io_request),
    .io_grant                       (issue_slots_17_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_16),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_17_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_72 ? _slots_21_io_out_uop_uopc : _GEN_71 ? _slots_20_io_out_uop_uopc : _GEN_70 ? _slots_19_io_out_uop_uopc : _slots_18_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_72 ? _slots_21_io_out_uop_inst : _GEN_71 ? _slots_20_io_out_uop_inst : _GEN_70 ? _slots_19_io_out_uop_inst : _slots_18_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_72 ? _slots_21_io_out_uop_debug_inst : _GEN_71 ? _slots_20_io_out_uop_debug_inst : _GEN_70 ? _slots_19_io_out_uop_debug_inst : _slots_18_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_72 ? _slots_21_io_out_uop_is_rvc : _GEN_71 ? _slots_20_io_out_uop_is_rvc : _GEN_70 ? _slots_19_io_out_uop_is_rvc : _slots_18_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_72 ? _slots_21_io_out_uop_debug_pc : _GEN_71 ? _slots_20_io_out_uop_debug_pc : _GEN_70 ? _slots_19_io_out_uop_debug_pc : _slots_18_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_72 ? _slots_21_io_out_uop_iq_type : _GEN_71 ? _slots_20_io_out_uop_iq_type : _GEN_70 ? _slots_19_io_out_uop_iq_type : _slots_18_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_72 ? _slots_21_io_out_uop_fu_code : _GEN_71 ? _slots_20_io_out_uop_fu_code : _GEN_70 ? _slots_19_io_out_uop_fu_code : _slots_18_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_72 ? _slots_21_io_out_uop_iw_state : _GEN_71 ? _slots_20_io_out_uop_iw_state : _GEN_70 ? _slots_19_io_out_uop_iw_state : _slots_18_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_72 ? _slots_21_io_out_uop_iw_p1_poisoned : _GEN_71 ? _slots_20_io_out_uop_iw_p1_poisoned : _GEN_70 ? _slots_19_io_out_uop_iw_p1_poisoned : _slots_18_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_72 ? _slots_21_io_out_uop_iw_p2_poisoned : _GEN_71 ? _slots_20_io_out_uop_iw_p2_poisoned : _GEN_70 ? _slots_19_io_out_uop_iw_p2_poisoned : _slots_18_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_72 ? _slots_21_io_out_uop_is_br : _GEN_71 ? _slots_20_io_out_uop_is_br : _GEN_70 ? _slots_19_io_out_uop_is_br : _slots_18_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_72 ? _slots_21_io_out_uop_is_jalr : _GEN_71 ? _slots_20_io_out_uop_is_jalr : _GEN_70 ? _slots_19_io_out_uop_is_jalr : _slots_18_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_72 ? _slots_21_io_out_uop_is_jal : _GEN_71 ? _slots_20_io_out_uop_is_jal : _GEN_70 ? _slots_19_io_out_uop_is_jal : _slots_18_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_72 ? _slots_21_io_out_uop_is_sfb : _GEN_71 ? _slots_20_io_out_uop_is_sfb : _GEN_70 ? _slots_19_io_out_uop_is_sfb : _slots_18_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_72 ? _slots_21_io_out_uop_br_mask : _GEN_71 ? _slots_20_io_out_uop_br_mask : _GEN_70 ? _slots_19_io_out_uop_br_mask : _slots_18_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_72 ? _slots_21_io_out_uop_br_tag : _GEN_71 ? _slots_20_io_out_uop_br_tag : _GEN_70 ? _slots_19_io_out_uop_br_tag : _slots_18_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_72 ? _slots_21_io_out_uop_ftq_idx : _GEN_71 ? _slots_20_io_out_uop_ftq_idx : _GEN_70 ? _slots_19_io_out_uop_ftq_idx : _slots_18_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_72 ? _slots_21_io_out_uop_edge_inst : _GEN_71 ? _slots_20_io_out_uop_edge_inst : _GEN_70 ? _slots_19_io_out_uop_edge_inst : _slots_18_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_72 ? _slots_21_io_out_uop_pc_lob : _GEN_71 ? _slots_20_io_out_uop_pc_lob : _GEN_70 ? _slots_19_io_out_uop_pc_lob : _slots_18_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_72 ? _slots_21_io_out_uop_taken : _GEN_71 ? _slots_20_io_out_uop_taken : _GEN_70 ? _slots_19_io_out_uop_taken : _slots_18_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_72 ? _slots_21_io_out_uop_imm_packed : _GEN_71 ? _slots_20_io_out_uop_imm_packed : _GEN_70 ? _slots_19_io_out_uop_imm_packed : _slots_18_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_72 ? _slots_21_io_out_uop_csr_addr : _GEN_71 ? _slots_20_io_out_uop_csr_addr : _GEN_70 ? _slots_19_io_out_uop_csr_addr : _slots_18_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_72 ? _slots_21_io_out_uop_rob_idx : _GEN_71 ? _slots_20_io_out_uop_rob_idx : _GEN_70 ? _slots_19_io_out_uop_rob_idx : _slots_18_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_72 ? _slots_21_io_out_uop_ldq_idx : _GEN_71 ? _slots_20_io_out_uop_ldq_idx : _GEN_70 ? _slots_19_io_out_uop_ldq_idx : _slots_18_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_72 ? _slots_21_io_out_uop_stq_idx : _GEN_71 ? _slots_20_io_out_uop_stq_idx : _GEN_70 ? _slots_19_io_out_uop_stq_idx : _slots_18_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_72 ? _slots_21_io_out_uop_rxq_idx : _GEN_71 ? _slots_20_io_out_uop_rxq_idx : _GEN_70 ? _slots_19_io_out_uop_rxq_idx : _slots_18_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_72 ? _slots_21_io_out_uop_pdst : _GEN_71 ? _slots_20_io_out_uop_pdst : _GEN_70 ? _slots_19_io_out_uop_pdst : _slots_18_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_72 ? _slots_21_io_out_uop_prs1 : _GEN_71 ? _slots_20_io_out_uop_prs1 : _GEN_70 ? _slots_19_io_out_uop_prs1 : _slots_18_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_72 ? _slots_21_io_out_uop_prs2 : _GEN_71 ? _slots_20_io_out_uop_prs2 : _GEN_70 ? _slots_19_io_out_uop_prs2 : _slots_18_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_72 ? _slots_21_io_out_uop_prs3 : _GEN_71 ? _slots_20_io_out_uop_prs3 : _GEN_70 ? _slots_19_io_out_uop_prs3 : _slots_18_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_72 ? _slots_21_io_out_uop_ppred : _GEN_71 ? _slots_20_io_out_uop_ppred : _GEN_70 ? _slots_19_io_out_uop_ppred : _slots_18_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_72 ? _slots_21_io_out_uop_prs1_busy : _GEN_71 ? _slots_20_io_out_uop_prs1_busy : _GEN_70 ? _slots_19_io_out_uop_prs1_busy : _slots_18_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_72 ? _slots_21_io_out_uop_prs2_busy : _GEN_71 ? _slots_20_io_out_uop_prs2_busy : _GEN_70 ? _slots_19_io_out_uop_prs2_busy : _slots_18_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_72 ? _slots_21_io_out_uop_prs3_busy : _GEN_71 ? _slots_20_io_out_uop_prs3_busy : _GEN_70 ? _slots_19_io_out_uop_prs3_busy : _slots_18_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_72 ? _slots_21_io_out_uop_ppred_busy : _GEN_71 ? _slots_20_io_out_uop_ppred_busy : _GEN_70 ? _slots_19_io_out_uop_ppred_busy : _slots_18_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_72 ? _slots_21_io_out_uop_stale_pdst : _GEN_71 ? _slots_20_io_out_uop_stale_pdst : _GEN_70 ? _slots_19_io_out_uop_stale_pdst : _slots_18_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_72 ? _slots_21_io_out_uop_exception : _GEN_71 ? _slots_20_io_out_uop_exception : _GEN_70 ? _slots_19_io_out_uop_exception : _slots_18_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_72 ? _slots_21_io_out_uop_exc_cause : _GEN_71 ? _slots_20_io_out_uop_exc_cause : _GEN_70 ? _slots_19_io_out_uop_exc_cause : _slots_18_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_72 ? _slots_21_io_out_uop_bypassable : _GEN_71 ? _slots_20_io_out_uop_bypassable : _GEN_70 ? _slots_19_io_out_uop_bypassable : _slots_18_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_72 ? _slots_21_io_out_uop_mem_cmd : _GEN_71 ? _slots_20_io_out_uop_mem_cmd : _GEN_70 ? _slots_19_io_out_uop_mem_cmd : _slots_18_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_72 ? _slots_21_io_out_uop_mem_size : _GEN_71 ? _slots_20_io_out_uop_mem_size : _GEN_70 ? _slots_19_io_out_uop_mem_size : _slots_18_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_72 ? _slots_21_io_out_uop_mem_signed : _GEN_71 ? _slots_20_io_out_uop_mem_signed : _GEN_70 ? _slots_19_io_out_uop_mem_signed : _slots_18_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_72 ? _slots_21_io_out_uop_is_fence : _GEN_71 ? _slots_20_io_out_uop_is_fence : _GEN_70 ? _slots_19_io_out_uop_is_fence : _slots_18_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_72 ? _slots_21_io_out_uop_is_fencei : _GEN_71 ? _slots_20_io_out_uop_is_fencei : _GEN_70 ? _slots_19_io_out_uop_is_fencei : _slots_18_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_72 ? _slots_21_io_out_uop_is_amo : _GEN_71 ? _slots_20_io_out_uop_is_amo : _GEN_70 ? _slots_19_io_out_uop_is_amo : _slots_18_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_72 ? _slots_21_io_out_uop_uses_ldq : _GEN_71 ? _slots_20_io_out_uop_uses_ldq : _GEN_70 ? _slots_19_io_out_uop_uses_ldq : _slots_18_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_72 ? _slots_21_io_out_uop_uses_stq : _GEN_71 ? _slots_20_io_out_uop_uses_stq : _GEN_70 ? _slots_19_io_out_uop_uses_stq : _slots_18_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_72 ? _slots_21_io_out_uop_is_sys_pc2epc : _GEN_71 ? _slots_20_io_out_uop_is_sys_pc2epc : _GEN_70 ? _slots_19_io_out_uop_is_sys_pc2epc : _slots_18_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_72 ? _slots_21_io_out_uop_is_unique : _GEN_71 ? _slots_20_io_out_uop_is_unique : _GEN_70 ? _slots_19_io_out_uop_is_unique : _slots_18_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_72 ? _slots_21_io_out_uop_flush_on_commit : _GEN_71 ? _slots_20_io_out_uop_flush_on_commit : _GEN_70 ? _slots_19_io_out_uop_flush_on_commit : _slots_18_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_72 ? _slots_21_io_out_uop_ldst_is_rs1 : _GEN_71 ? _slots_20_io_out_uop_ldst_is_rs1 : _GEN_70 ? _slots_19_io_out_uop_ldst_is_rs1 : _slots_18_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_72 ? _slots_21_io_out_uop_ldst : _GEN_71 ? _slots_20_io_out_uop_ldst : _GEN_70 ? _slots_19_io_out_uop_ldst : _slots_18_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_72 ? _slots_21_io_out_uop_lrs1 : _GEN_71 ? _slots_20_io_out_uop_lrs1 : _GEN_70 ? _slots_19_io_out_uop_lrs1 : _slots_18_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_72 ? _slots_21_io_out_uop_lrs2 : _GEN_71 ? _slots_20_io_out_uop_lrs2 : _GEN_70 ? _slots_19_io_out_uop_lrs2 : _slots_18_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_72 ? _slots_21_io_out_uop_lrs3 : _GEN_71 ? _slots_20_io_out_uop_lrs3 : _GEN_70 ? _slots_19_io_out_uop_lrs3 : _slots_18_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_72 ? _slots_21_io_out_uop_ldst_val : _GEN_71 ? _slots_20_io_out_uop_ldst_val : _GEN_70 ? _slots_19_io_out_uop_ldst_val : _slots_18_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_72 ? _slots_21_io_out_uop_dst_rtype : _GEN_71 ? _slots_20_io_out_uop_dst_rtype : _GEN_70 ? _slots_19_io_out_uop_dst_rtype : _slots_18_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_72 ? _slots_21_io_out_uop_lrs1_rtype : _GEN_71 ? _slots_20_io_out_uop_lrs1_rtype : _GEN_70 ? _slots_19_io_out_uop_lrs1_rtype : _slots_18_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_72 ? _slots_21_io_out_uop_lrs2_rtype : _GEN_71 ? _slots_20_io_out_uop_lrs2_rtype : _GEN_70 ? _slots_19_io_out_uop_lrs2_rtype : _slots_18_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_72 ? _slots_21_io_out_uop_frs3_en : _GEN_71 ? _slots_20_io_out_uop_frs3_en : _GEN_70 ? _slots_19_io_out_uop_frs3_en : _slots_18_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_72 ? _slots_21_io_out_uop_fp_val : _GEN_71 ? _slots_20_io_out_uop_fp_val : _GEN_70 ? _slots_19_io_out_uop_fp_val : _slots_18_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_72 ? _slots_21_io_out_uop_fp_single : _GEN_71 ? _slots_20_io_out_uop_fp_single : _GEN_70 ? _slots_19_io_out_uop_fp_single : _slots_18_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_72 ? _slots_21_io_out_uop_xcpt_pf_if : _GEN_71 ? _slots_20_io_out_uop_xcpt_pf_if : _GEN_70 ? _slots_19_io_out_uop_xcpt_pf_if : _slots_18_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_72 ? _slots_21_io_out_uop_xcpt_ae_if : _GEN_71 ? _slots_20_io_out_uop_xcpt_ae_if : _GEN_70 ? _slots_19_io_out_uop_xcpt_ae_if : _slots_18_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_72 ? _slots_21_io_out_uop_xcpt_ma_if : _GEN_71 ? _slots_20_io_out_uop_xcpt_ma_if : _GEN_70 ? _slots_19_io_out_uop_xcpt_ma_if : _slots_18_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_72 ? _slots_21_io_out_uop_bp_debug_if : _GEN_71 ? _slots_20_io_out_uop_bp_debug_if : _GEN_70 ? _slots_19_io_out_uop_bp_debug_if : _slots_18_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_72 ? _slots_21_io_out_uop_bp_xcpt_if : _GEN_71 ? _slots_20_io_out_uop_bp_xcpt_if : _GEN_70 ? _slots_19_io_out_uop_bp_xcpt_if : _slots_18_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_72 ? _slots_21_io_out_uop_debug_fsrc : _GEN_71 ? _slots_20_io_out_uop_debug_fsrc : _GEN_70 ? _slots_19_io_out_uop_debug_fsrc : _slots_18_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_72 ? _slots_21_io_out_uop_debug_tsrc : _GEN_71 ? _slots_20_io_out_uop_debug_tsrc : _GEN_70 ? _slots_19_io_out_uop_debug_tsrc : _slots_18_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_17_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_17_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_17_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_17_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_17_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_17_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_17_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_17_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_17_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_17_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_17_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_17_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_17_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_17_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_17_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_17_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_17_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_17_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_17_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_17_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_17_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_17_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_17_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_17_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_17_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_17_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_17_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_17_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_17_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_17_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_17_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_17_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_17_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_17_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_17_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_17_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_17_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_17_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_17_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_17_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_17_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_17_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_17_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_17_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_17_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_17_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_17_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_17_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_17_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_17_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_17_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_17_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_17_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_17_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_17_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_17_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_17_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_17_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_17_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_17_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_17_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_17_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_17_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_17_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_17_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_17_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_17_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_17_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_17_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_17_io_uop_uopc),
    .io_uop_inst                    (_slots_17_io_uop_inst),
    .io_uop_debug_inst              (_slots_17_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_17_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_17_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_17_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_17_io_uop_fu_code),
    .io_uop_iw_state                (_slots_17_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_17_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_17_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_17_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_17_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_17_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_17_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_17_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_17_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_17_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_17_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_17_io_uop_pc_lob),
    .io_uop_taken                   (_slots_17_io_uop_taken),
    .io_uop_imm_packed              (_slots_17_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_17_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_17_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_17_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_17_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_17_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_17_io_uop_pdst),
    .io_uop_prs1                    (_slots_17_io_uop_prs1),
    .io_uop_prs2                    (_slots_17_io_uop_prs2),
    .io_uop_prs3                    (_slots_17_io_uop_prs3),
    .io_uop_ppred                   (_slots_17_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_17_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_17_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_17_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_17_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_17_io_uop_stale_pdst),
    .io_uop_exception               (_slots_17_io_uop_exception),
    .io_uop_exc_cause               (_slots_17_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_17_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_17_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_17_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_17_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_17_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_17_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_17_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_17_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_17_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_17_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_17_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_17_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_17_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_17_io_uop_ldst),
    .io_uop_lrs1                    (_slots_17_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_17_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_17_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_17_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_17_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_17_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_17_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_17_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_17_io_uop_fp_val),
    .io_uop_fp_single               (_slots_17_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_17_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_17_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_17_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_17_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_17_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_17_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_17_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_18 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_18_io_valid),
    .io_will_be_valid               (_slots_18_io_will_be_valid),
    .io_request                     (_slots_18_io_request),
    .io_grant                       (issue_slots_18_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_17),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_18_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_75 ? _slots_22_io_out_uop_uopc : _GEN_74 ? _slots_21_io_out_uop_uopc : _GEN_73 ? _slots_20_io_out_uop_uopc : _slots_19_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_75 ? _slots_22_io_out_uop_inst : _GEN_74 ? _slots_21_io_out_uop_inst : _GEN_73 ? _slots_20_io_out_uop_inst : _slots_19_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_75 ? _slots_22_io_out_uop_debug_inst : _GEN_74 ? _slots_21_io_out_uop_debug_inst : _GEN_73 ? _slots_20_io_out_uop_debug_inst : _slots_19_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_75 ? _slots_22_io_out_uop_is_rvc : _GEN_74 ? _slots_21_io_out_uop_is_rvc : _GEN_73 ? _slots_20_io_out_uop_is_rvc : _slots_19_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_75 ? _slots_22_io_out_uop_debug_pc : _GEN_74 ? _slots_21_io_out_uop_debug_pc : _GEN_73 ? _slots_20_io_out_uop_debug_pc : _slots_19_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_75 ? _slots_22_io_out_uop_iq_type : _GEN_74 ? _slots_21_io_out_uop_iq_type : _GEN_73 ? _slots_20_io_out_uop_iq_type : _slots_19_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_75 ? _slots_22_io_out_uop_fu_code : _GEN_74 ? _slots_21_io_out_uop_fu_code : _GEN_73 ? _slots_20_io_out_uop_fu_code : _slots_19_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_75 ? _slots_22_io_out_uop_iw_state : _GEN_74 ? _slots_21_io_out_uop_iw_state : _GEN_73 ? _slots_20_io_out_uop_iw_state : _slots_19_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_75 ? _slots_22_io_out_uop_iw_p1_poisoned : _GEN_74 ? _slots_21_io_out_uop_iw_p1_poisoned : _GEN_73 ? _slots_20_io_out_uop_iw_p1_poisoned : _slots_19_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_75 ? _slots_22_io_out_uop_iw_p2_poisoned : _GEN_74 ? _slots_21_io_out_uop_iw_p2_poisoned : _GEN_73 ? _slots_20_io_out_uop_iw_p2_poisoned : _slots_19_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_75 ? _slots_22_io_out_uop_is_br : _GEN_74 ? _slots_21_io_out_uop_is_br : _GEN_73 ? _slots_20_io_out_uop_is_br : _slots_19_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_75 ? _slots_22_io_out_uop_is_jalr : _GEN_74 ? _slots_21_io_out_uop_is_jalr : _GEN_73 ? _slots_20_io_out_uop_is_jalr : _slots_19_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_75 ? _slots_22_io_out_uop_is_jal : _GEN_74 ? _slots_21_io_out_uop_is_jal : _GEN_73 ? _slots_20_io_out_uop_is_jal : _slots_19_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_75 ? _slots_22_io_out_uop_is_sfb : _GEN_74 ? _slots_21_io_out_uop_is_sfb : _GEN_73 ? _slots_20_io_out_uop_is_sfb : _slots_19_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_75 ? _slots_22_io_out_uop_br_mask : _GEN_74 ? _slots_21_io_out_uop_br_mask : _GEN_73 ? _slots_20_io_out_uop_br_mask : _slots_19_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_75 ? _slots_22_io_out_uop_br_tag : _GEN_74 ? _slots_21_io_out_uop_br_tag : _GEN_73 ? _slots_20_io_out_uop_br_tag : _slots_19_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_75 ? _slots_22_io_out_uop_ftq_idx : _GEN_74 ? _slots_21_io_out_uop_ftq_idx : _GEN_73 ? _slots_20_io_out_uop_ftq_idx : _slots_19_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_75 ? _slots_22_io_out_uop_edge_inst : _GEN_74 ? _slots_21_io_out_uop_edge_inst : _GEN_73 ? _slots_20_io_out_uop_edge_inst : _slots_19_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_75 ? _slots_22_io_out_uop_pc_lob : _GEN_74 ? _slots_21_io_out_uop_pc_lob : _GEN_73 ? _slots_20_io_out_uop_pc_lob : _slots_19_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_75 ? _slots_22_io_out_uop_taken : _GEN_74 ? _slots_21_io_out_uop_taken : _GEN_73 ? _slots_20_io_out_uop_taken : _slots_19_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_75 ? _slots_22_io_out_uop_imm_packed : _GEN_74 ? _slots_21_io_out_uop_imm_packed : _GEN_73 ? _slots_20_io_out_uop_imm_packed : _slots_19_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_75 ? _slots_22_io_out_uop_csr_addr : _GEN_74 ? _slots_21_io_out_uop_csr_addr : _GEN_73 ? _slots_20_io_out_uop_csr_addr : _slots_19_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_75 ? _slots_22_io_out_uop_rob_idx : _GEN_74 ? _slots_21_io_out_uop_rob_idx : _GEN_73 ? _slots_20_io_out_uop_rob_idx : _slots_19_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_75 ? _slots_22_io_out_uop_ldq_idx : _GEN_74 ? _slots_21_io_out_uop_ldq_idx : _GEN_73 ? _slots_20_io_out_uop_ldq_idx : _slots_19_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_75 ? _slots_22_io_out_uop_stq_idx : _GEN_74 ? _slots_21_io_out_uop_stq_idx : _GEN_73 ? _slots_20_io_out_uop_stq_idx : _slots_19_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_75 ? _slots_22_io_out_uop_rxq_idx : _GEN_74 ? _slots_21_io_out_uop_rxq_idx : _GEN_73 ? _slots_20_io_out_uop_rxq_idx : _slots_19_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_75 ? _slots_22_io_out_uop_pdst : _GEN_74 ? _slots_21_io_out_uop_pdst : _GEN_73 ? _slots_20_io_out_uop_pdst : _slots_19_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_75 ? _slots_22_io_out_uop_prs1 : _GEN_74 ? _slots_21_io_out_uop_prs1 : _GEN_73 ? _slots_20_io_out_uop_prs1 : _slots_19_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_75 ? _slots_22_io_out_uop_prs2 : _GEN_74 ? _slots_21_io_out_uop_prs2 : _GEN_73 ? _slots_20_io_out_uop_prs2 : _slots_19_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_75 ? _slots_22_io_out_uop_prs3 : _GEN_74 ? _slots_21_io_out_uop_prs3 : _GEN_73 ? _slots_20_io_out_uop_prs3 : _slots_19_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_75 ? _slots_22_io_out_uop_ppred : _GEN_74 ? _slots_21_io_out_uop_ppred : _GEN_73 ? _slots_20_io_out_uop_ppred : _slots_19_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_75 ? _slots_22_io_out_uop_prs1_busy : _GEN_74 ? _slots_21_io_out_uop_prs1_busy : _GEN_73 ? _slots_20_io_out_uop_prs1_busy : _slots_19_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_75 ? _slots_22_io_out_uop_prs2_busy : _GEN_74 ? _slots_21_io_out_uop_prs2_busy : _GEN_73 ? _slots_20_io_out_uop_prs2_busy : _slots_19_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_75 ? _slots_22_io_out_uop_prs3_busy : _GEN_74 ? _slots_21_io_out_uop_prs3_busy : _GEN_73 ? _slots_20_io_out_uop_prs3_busy : _slots_19_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_75 ? _slots_22_io_out_uop_ppred_busy : _GEN_74 ? _slots_21_io_out_uop_ppred_busy : _GEN_73 ? _slots_20_io_out_uop_ppred_busy : _slots_19_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_75 ? _slots_22_io_out_uop_stale_pdst : _GEN_74 ? _slots_21_io_out_uop_stale_pdst : _GEN_73 ? _slots_20_io_out_uop_stale_pdst : _slots_19_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_75 ? _slots_22_io_out_uop_exception : _GEN_74 ? _slots_21_io_out_uop_exception : _GEN_73 ? _slots_20_io_out_uop_exception : _slots_19_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_75 ? _slots_22_io_out_uop_exc_cause : _GEN_74 ? _slots_21_io_out_uop_exc_cause : _GEN_73 ? _slots_20_io_out_uop_exc_cause : _slots_19_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_75 ? _slots_22_io_out_uop_bypassable : _GEN_74 ? _slots_21_io_out_uop_bypassable : _GEN_73 ? _slots_20_io_out_uop_bypassable : _slots_19_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_75 ? _slots_22_io_out_uop_mem_cmd : _GEN_74 ? _slots_21_io_out_uop_mem_cmd : _GEN_73 ? _slots_20_io_out_uop_mem_cmd : _slots_19_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_75 ? _slots_22_io_out_uop_mem_size : _GEN_74 ? _slots_21_io_out_uop_mem_size : _GEN_73 ? _slots_20_io_out_uop_mem_size : _slots_19_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_75 ? _slots_22_io_out_uop_mem_signed : _GEN_74 ? _slots_21_io_out_uop_mem_signed : _GEN_73 ? _slots_20_io_out_uop_mem_signed : _slots_19_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_75 ? _slots_22_io_out_uop_is_fence : _GEN_74 ? _slots_21_io_out_uop_is_fence : _GEN_73 ? _slots_20_io_out_uop_is_fence : _slots_19_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_75 ? _slots_22_io_out_uop_is_fencei : _GEN_74 ? _slots_21_io_out_uop_is_fencei : _GEN_73 ? _slots_20_io_out_uop_is_fencei : _slots_19_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_75 ? _slots_22_io_out_uop_is_amo : _GEN_74 ? _slots_21_io_out_uop_is_amo : _GEN_73 ? _slots_20_io_out_uop_is_amo : _slots_19_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_75 ? _slots_22_io_out_uop_uses_ldq : _GEN_74 ? _slots_21_io_out_uop_uses_ldq : _GEN_73 ? _slots_20_io_out_uop_uses_ldq : _slots_19_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_75 ? _slots_22_io_out_uop_uses_stq : _GEN_74 ? _slots_21_io_out_uop_uses_stq : _GEN_73 ? _slots_20_io_out_uop_uses_stq : _slots_19_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_75 ? _slots_22_io_out_uop_is_sys_pc2epc : _GEN_74 ? _slots_21_io_out_uop_is_sys_pc2epc : _GEN_73 ? _slots_20_io_out_uop_is_sys_pc2epc : _slots_19_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_75 ? _slots_22_io_out_uop_is_unique : _GEN_74 ? _slots_21_io_out_uop_is_unique : _GEN_73 ? _slots_20_io_out_uop_is_unique : _slots_19_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_75 ? _slots_22_io_out_uop_flush_on_commit : _GEN_74 ? _slots_21_io_out_uop_flush_on_commit : _GEN_73 ? _slots_20_io_out_uop_flush_on_commit : _slots_19_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_75 ? _slots_22_io_out_uop_ldst_is_rs1 : _GEN_74 ? _slots_21_io_out_uop_ldst_is_rs1 : _GEN_73 ? _slots_20_io_out_uop_ldst_is_rs1 : _slots_19_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_75 ? _slots_22_io_out_uop_ldst : _GEN_74 ? _slots_21_io_out_uop_ldst : _GEN_73 ? _slots_20_io_out_uop_ldst : _slots_19_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_75 ? _slots_22_io_out_uop_lrs1 : _GEN_74 ? _slots_21_io_out_uop_lrs1 : _GEN_73 ? _slots_20_io_out_uop_lrs1 : _slots_19_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_75 ? _slots_22_io_out_uop_lrs2 : _GEN_74 ? _slots_21_io_out_uop_lrs2 : _GEN_73 ? _slots_20_io_out_uop_lrs2 : _slots_19_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_75 ? _slots_22_io_out_uop_lrs3 : _GEN_74 ? _slots_21_io_out_uop_lrs3 : _GEN_73 ? _slots_20_io_out_uop_lrs3 : _slots_19_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_75 ? _slots_22_io_out_uop_ldst_val : _GEN_74 ? _slots_21_io_out_uop_ldst_val : _GEN_73 ? _slots_20_io_out_uop_ldst_val : _slots_19_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_75 ? _slots_22_io_out_uop_dst_rtype : _GEN_74 ? _slots_21_io_out_uop_dst_rtype : _GEN_73 ? _slots_20_io_out_uop_dst_rtype : _slots_19_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_75 ? _slots_22_io_out_uop_lrs1_rtype : _GEN_74 ? _slots_21_io_out_uop_lrs1_rtype : _GEN_73 ? _slots_20_io_out_uop_lrs1_rtype : _slots_19_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_75 ? _slots_22_io_out_uop_lrs2_rtype : _GEN_74 ? _slots_21_io_out_uop_lrs2_rtype : _GEN_73 ? _slots_20_io_out_uop_lrs2_rtype : _slots_19_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_75 ? _slots_22_io_out_uop_frs3_en : _GEN_74 ? _slots_21_io_out_uop_frs3_en : _GEN_73 ? _slots_20_io_out_uop_frs3_en : _slots_19_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_75 ? _slots_22_io_out_uop_fp_val : _GEN_74 ? _slots_21_io_out_uop_fp_val : _GEN_73 ? _slots_20_io_out_uop_fp_val : _slots_19_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_75 ? _slots_22_io_out_uop_fp_single : _GEN_74 ? _slots_21_io_out_uop_fp_single : _GEN_73 ? _slots_20_io_out_uop_fp_single : _slots_19_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_75 ? _slots_22_io_out_uop_xcpt_pf_if : _GEN_74 ? _slots_21_io_out_uop_xcpt_pf_if : _GEN_73 ? _slots_20_io_out_uop_xcpt_pf_if : _slots_19_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_75 ? _slots_22_io_out_uop_xcpt_ae_if : _GEN_74 ? _slots_21_io_out_uop_xcpt_ae_if : _GEN_73 ? _slots_20_io_out_uop_xcpt_ae_if : _slots_19_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_75 ? _slots_22_io_out_uop_xcpt_ma_if : _GEN_74 ? _slots_21_io_out_uop_xcpt_ma_if : _GEN_73 ? _slots_20_io_out_uop_xcpt_ma_if : _slots_19_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_75 ? _slots_22_io_out_uop_bp_debug_if : _GEN_74 ? _slots_21_io_out_uop_bp_debug_if : _GEN_73 ? _slots_20_io_out_uop_bp_debug_if : _slots_19_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_75 ? _slots_22_io_out_uop_bp_xcpt_if : _GEN_74 ? _slots_21_io_out_uop_bp_xcpt_if : _GEN_73 ? _slots_20_io_out_uop_bp_xcpt_if : _slots_19_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_75 ? _slots_22_io_out_uop_debug_fsrc : _GEN_74 ? _slots_21_io_out_uop_debug_fsrc : _GEN_73 ? _slots_20_io_out_uop_debug_fsrc : _slots_19_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_75 ? _slots_22_io_out_uop_debug_tsrc : _GEN_74 ? _slots_21_io_out_uop_debug_tsrc : _GEN_73 ? _slots_20_io_out_uop_debug_tsrc : _slots_19_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_18_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_18_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_18_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_18_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_18_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_18_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_18_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_18_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_18_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_18_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_18_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_18_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_18_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_18_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_18_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_18_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_18_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_18_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_18_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_18_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_18_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_18_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_18_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_18_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_18_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_18_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_18_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_18_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_18_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_18_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_18_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_18_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_18_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_18_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_18_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_18_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_18_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_18_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_18_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_18_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_18_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_18_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_18_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_18_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_18_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_18_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_18_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_18_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_18_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_18_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_18_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_18_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_18_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_18_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_18_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_18_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_18_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_18_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_18_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_18_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_18_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_18_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_18_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_18_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_18_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_18_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_18_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_18_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_18_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_18_io_uop_uopc),
    .io_uop_inst                    (_slots_18_io_uop_inst),
    .io_uop_debug_inst              (_slots_18_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_18_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_18_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_18_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_18_io_uop_fu_code),
    .io_uop_iw_state                (_slots_18_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_18_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_18_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_18_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_18_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_18_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_18_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_18_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_18_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_18_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_18_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_18_io_uop_pc_lob),
    .io_uop_taken                   (_slots_18_io_uop_taken),
    .io_uop_imm_packed              (_slots_18_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_18_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_18_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_18_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_18_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_18_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_18_io_uop_pdst),
    .io_uop_prs1                    (_slots_18_io_uop_prs1),
    .io_uop_prs2                    (_slots_18_io_uop_prs2),
    .io_uop_prs3                    (_slots_18_io_uop_prs3),
    .io_uop_ppred                   (_slots_18_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_18_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_18_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_18_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_18_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_18_io_uop_stale_pdst),
    .io_uop_exception               (_slots_18_io_uop_exception),
    .io_uop_exc_cause               (_slots_18_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_18_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_18_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_18_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_18_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_18_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_18_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_18_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_18_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_18_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_18_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_18_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_18_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_18_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_18_io_uop_ldst),
    .io_uop_lrs1                    (_slots_18_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_18_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_18_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_18_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_18_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_18_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_18_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_18_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_18_io_uop_fp_val),
    .io_uop_fp_single               (_slots_18_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_18_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_18_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_18_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_18_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_18_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_18_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_18_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_19 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_19_io_valid),
    .io_will_be_valid               (_slots_19_io_will_be_valid),
    .io_request                     (_slots_19_io_request),
    .io_grant                       (issue_slots_19_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_18),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_19_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_78 ? _slots_23_io_out_uop_uopc : _GEN_77 ? _slots_22_io_out_uop_uopc : _GEN_76 ? _slots_21_io_out_uop_uopc : _slots_20_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_78 ? _slots_23_io_out_uop_inst : _GEN_77 ? _slots_22_io_out_uop_inst : _GEN_76 ? _slots_21_io_out_uop_inst : _slots_20_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_78 ? _slots_23_io_out_uop_debug_inst : _GEN_77 ? _slots_22_io_out_uop_debug_inst : _GEN_76 ? _slots_21_io_out_uop_debug_inst : _slots_20_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_78 ? _slots_23_io_out_uop_is_rvc : _GEN_77 ? _slots_22_io_out_uop_is_rvc : _GEN_76 ? _slots_21_io_out_uop_is_rvc : _slots_20_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_78 ? _slots_23_io_out_uop_debug_pc : _GEN_77 ? _slots_22_io_out_uop_debug_pc : _GEN_76 ? _slots_21_io_out_uop_debug_pc : _slots_20_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_78 ? _slots_23_io_out_uop_iq_type : _GEN_77 ? _slots_22_io_out_uop_iq_type : _GEN_76 ? _slots_21_io_out_uop_iq_type : _slots_20_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_78 ? _slots_23_io_out_uop_fu_code : _GEN_77 ? _slots_22_io_out_uop_fu_code : _GEN_76 ? _slots_21_io_out_uop_fu_code : _slots_20_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_78 ? _slots_23_io_out_uop_iw_state : _GEN_77 ? _slots_22_io_out_uop_iw_state : _GEN_76 ? _slots_21_io_out_uop_iw_state : _slots_20_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_78 ? _slots_23_io_out_uop_iw_p1_poisoned : _GEN_77 ? _slots_22_io_out_uop_iw_p1_poisoned : _GEN_76 ? _slots_21_io_out_uop_iw_p1_poisoned : _slots_20_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_78 ? _slots_23_io_out_uop_iw_p2_poisoned : _GEN_77 ? _slots_22_io_out_uop_iw_p2_poisoned : _GEN_76 ? _slots_21_io_out_uop_iw_p2_poisoned : _slots_20_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_78 ? _slots_23_io_out_uop_is_br : _GEN_77 ? _slots_22_io_out_uop_is_br : _GEN_76 ? _slots_21_io_out_uop_is_br : _slots_20_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_78 ? _slots_23_io_out_uop_is_jalr : _GEN_77 ? _slots_22_io_out_uop_is_jalr : _GEN_76 ? _slots_21_io_out_uop_is_jalr : _slots_20_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_78 ? _slots_23_io_out_uop_is_jal : _GEN_77 ? _slots_22_io_out_uop_is_jal : _GEN_76 ? _slots_21_io_out_uop_is_jal : _slots_20_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_78 ? _slots_23_io_out_uop_is_sfb : _GEN_77 ? _slots_22_io_out_uop_is_sfb : _GEN_76 ? _slots_21_io_out_uop_is_sfb : _slots_20_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_78 ? _slots_23_io_out_uop_br_mask : _GEN_77 ? _slots_22_io_out_uop_br_mask : _GEN_76 ? _slots_21_io_out_uop_br_mask : _slots_20_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_78 ? _slots_23_io_out_uop_br_tag : _GEN_77 ? _slots_22_io_out_uop_br_tag : _GEN_76 ? _slots_21_io_out_uop_br_tag : _slots_20_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_78 ? _slots_23_io_out_uop_ftq_idx : _GEN_77 ? _slots_22_io_out_uop_ftq_idx : _GEN_76 ? _slots_21_io_out_uop_ftq_idx : _slots_20_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_78 ? _slots_23_io_out_uop_edge_inst : _GEN_77 ? _slots_22_io_out_uop_edge_inst : _GEN_76 ? _slots_21_io_out_uop_edge_inst : _slots_20_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_78 ? _slots_23_io_out_uop_pc_lob : _GEN_77 ? _slots_22_io_out_uop_pc_lob : _GEN_76 ? _slots_21_io_out_uop_pc_lob : _slots_20_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_78 ? _slots_23_io_out_uop_taken : _GEN_77 ? _slots_22_io_out_uop_taken : _GEN_76 ? _slots_21_io_out_uop_taken : _slots_20_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_78 ? _slots_23_io_out_uop_imm_packed : _GEN_77 ? _slots_22_io_out_uop_imm_packed : _GEN_76 ? _slots_21_io_out_uop_imm_packed : _slots_20_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_78 ? _slots_23_io_out_uop_csr_addr : _GEN_77 ? _slots_22_io_out_uop_csr_addr : _GEN_76 ? _slots_21_io_out_uop_csr_addr : _slots_20_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_78 ? _slots_23_io_out_uop_rob_idx : _GEN_77 ? _slots_22_io_out_uop_rob_idx : _GEN_76 ? _slots_21_io_out_uop_rob_idx : _slots_20_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_78 ? _slots_23_io_out_uop_ldq_idx : _GEN_77 ? _slots_22_io_out_uop_ldq_idx : _GEN_76 ? _slots_21_io_out_uop_ldq_idx : _slots_20_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_78 ? _slots_23_io_out_uop_stq_idx : _GEN_77 ? _slots_22_io_out_uop_stq_idx : _GEN_76 ? _slots_21_io_out_uop_stq_idx : _slots_20_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_78 ? _slots_23_io_out_uop_rxq_idx : _GEN_77 ? _slots_22_io_out_uop_rxq_idx : _GEN_76 ? _slots_21_io_out_uop_rxq_idx : _slots_20_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_78 ? _slots_23_io_out_uop_pdst : _GEN_77 ? _slots_22_io_out_uop_pdst : _GEN_76 ? _slots_21_io_out_uop_pdst : _slots_20_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_78 ? _slots_23_io_out_uop_prs1 : _GEN_77 ? _slots_22_io_out_uop_prs1 : _GEN_76 ? _slots_21_io_out_uop_prs1 : _slots_20_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_78 ? _slots_23_io_out_uop_prs2 : _GEN_77 ? _slots_22_io_out_uop_prs2 : _GEN_76 ? _slots_21_io_out_uop_prs2 : _slots_20_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_78 ? _slots_23_io_out_uop_prs3 : _GEN_77 ? _slots_22_io_out_uop_prs3 : _GEN_76 ? _slots_21_io_out_uop_prs3 : _slots_20_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_78 ? _slots_23_io_out_uop_ppred : _GEN_77 ? _slots_22_io_out_uop_ppred : _GEN_76 ? _slots_21_io_out_uop_ppred : _slots_20_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_78 ? _slots_23_io_out_uop_prs1_busy : _GEN_77 ? _slots_22_io_out_uop_prs1_busy : _GEN_76 ? _slots_21_io_out_uop_prs1_busy : _slots_20_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_78 ? _slots_23_io_out_uop_prs2_busy : _GEN_77 ? _slots_22_io_out_uop_prs2_busy : _GEN_76 ? _slots_21_io_out_uop_prs2_busy : _slots_20_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_78 ? _slots_23_io_out_uop_prs3_busy : _GEN_77 ? _slots_22_io_out_uop_prs3_busy : _GEN_76 ? _slots_21_io_out_uop_prs3_busy : _slots_20_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_78 ? _slots_23_io_out_uop_ppred_busy : _GEN_77 ? _slots_22_io_out_uop_ppred_busy : _GEN_76 ? _slots_21_io_out_uop_ppred_busy : _slots_20_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_78 ? _slots_23_io_out_uop_stale_pdst : _GEN_77 ? _slots_22_io_out_uop_stale_pdst : _GEN_76 ? _slots_21_io_out_uop_stale_pdst : _slots_20_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_78 ? _slots_23_io_out_uop_exception : _GEN_77 ? _slots_22_io_out_uop_exception : _GEN_76 ? _slots_21_io_out_uop_exception : _slots_20_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_78 ? _slots_23_io_out_uop_exc_cause : _GEN_77 ? _slots_22_io_out_uop_exc_cause : _GEN_76 ? _slots_21_io_out_uop_exc_cause : _slots_20_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_78 ? _slots_23_io_out_uop_bypassable : _GEN_77 ? _slots_22_io_out_uop_bypassable : _GEN_76 ? _slots_21_io_out_uop_bypassable : _slots_20_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_78 ? _slots_23_io_out_uop_mem_cmd : _GEN_77 ? _slots_22_io_out_uop_mem_cmd : _GEN_76 ? _slots_21_io_out_uop_mem_cmd : _slots_20_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_78 ? _slots_23_io_out_uop_mem_size : _GEN_77 ? _slots_22_io_out_uop_mem_size : _GEN_76 ? _slots_21_io_out_uop_mem_size : _slots_20_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_78 ? _slots_23_io_out_uop_mem_signed : _GEN_77 ? _slots_22_io_out_uop_mem_signed : _GEN_76 ? _slots_21_io_out_uop_mem_signed : _slots_20_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_78 ? _slots_23_io_out_uop_is_fence : _GEN_77 ? _slots_22_io_out_uop_is_fence : _GEN_76 ? _slots_21_io_out_uop_is_fence : _slots_20_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_78 ? _slots_23_io_out_uop_is_fencei : _GEN_77 ? _slots_22_io_out_uop_is_fencei : _GEN_76 ? _slots_21_io_out_uop_is_fencei : _slots_20_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_78 ? _slots_23_io_out_uop_is_amo : _GEN_77 ? _slots_22_io_out_uop_is_amo : _GEN_76 ? _slots_21_io_out_uop_is_amo : _slots_20_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_78 ? _slots_23_io_out_uop_uses_ldq : _GEN_77 ? _slots_22_io_out_uop_uses_ldq : _GEN_76 ? _slots_21_io_out_uop_uses_ldq : _slots_20_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_78 ? _slots_23_io_out_uop_uses_stq : _GEN_77 ? _slots_22_io_out_uop_uses_stq : _GEN_76 ? _slots_21_io_out_uop_uses_stq : _slots_20_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_78 ? _slots_23_io_out_uop_is_sys_pc2epc : _GEN_77 ? _slots_22_io_out_uop_is_sys_pc2epc : _GEN_76 ? _slots_21_io_out_uop_is_sys_pc2epc : _slots_20_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_78 ? _slots_23_io_out_uop_is_unique : _GEN_77 ? _slots_22_io_out_uop_is_unique : _GEN_76 ? _slots_21_io_out_uop_is_unique : _slots_20_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_78 ? _slots_23_io_out_uop_flush_on_commit : _GEN_77 ? _slots_22_io_out_uop_flush_on_commit : _GEN_76 ? _slots_21_io_out_uop_flush_on_commit : _slots_20_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_78 ? _slots_23_io_out_uop_ldst_is_rs1 : _GEN_77 ? _slots_22_io_out_uop_ldst_is_rs1 : _GEN_76 ? _slots_21_io_out_uop_ldst_is_rs1 : _slots_20_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_78 ? _slots_23_io_out_uop_ldst : _GEN_77 ? _slots_22_io_out_uop_ldst : _GEN_76 ? _slots_21_io_out_uop_ldst : _slots_20_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_78 ? _slots_23_io_out_uop_lrs1 : _GEN_77 ? _slots_22_io_out_uop_lrs1 : _GEN_76 ? _slots_21_io_out_uop_lrs1 : _slots_20_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_78 ? _slots_23_io_out_uop_lrs2 : _GEN_77 ? _slots_22_io_out_uop_lrs2 : _GEN_76 ? _slots_21_io_out_uop_lrs2 : _slots_20_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_78 ? _slots_23_io_out_uop_lrs3 : _GEN_77 ? _slots_22_io_out_uop_lrs3 : _GEN_76 ? _slots_21_io_out_uop_lrs3 : _slots_20_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_78 ? _slots_23_io_out_uop_ldst_val : _GEN_77 ? _slots_22_io_out_uop_ldst_val : _GEN_76 ? _slots_21_io_out_uop_ldst_val : _slots_20_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_78 ? _slots_23_io_out_uop_dst_rtype : _GEN_77 ? _slots_22_io_out_uop_dst_rtype : _GEN_76 ? _slots_21_io_out_uop_dst_rtype : _slots_20_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_78 ? _slots_23_io_out_uop_lrs1_rtype : _GEN_77 ? _slots_22_io_out_uop_lrs1_rtype : _GEN_76 ? _slots_21_io_out_uop_lrs1_rtype : _slots_20_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_78 ? _slots_23_io_out_uop_lrs2_rtype : _GEN_77 ? _slots_22_io_out_uop_lrs2_rtype : _GEN_76 ? _slots_21_io_out_uop_lrs2_rtype : _slots_20_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_78 ? _slots_23_io_out_uop_frs3_en : _GEN_77 ? _slots_22_io_out_uop_frs3_en : _GEN_76 ? _slots_21_io_out_uop_frs3_en : _slots_20_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_78 ? _slots_23_io_out_uop_fp_val : _GEN_77 ? _slots_22_io_out_uop_fp_val : _GEN_76 ? _slots_21_io_out_uop_fp_val : _slots_20_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_78 ? _slots_23_io_out_uop_fp_single : _GEN_77 ? _slots_22_io_out_uop_fp_single : _GEN_76 ? _slots_21_io_out_uop_fp_single : _slots_20_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_78 ? _slots_23_io_out_uop_xcpt_pf_if : _GEN_77 ? _slots_22_io_out_uop_xcpt_pf_if : _GEN_76 ? _slots_21_io_out_uop_xcpt_pf_if : _slots_20_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_78 ? _slots_23_io_out_uop_xcpt_ae_if : _GEN_77 ? _slots_22_io_out_uop_xcpt_ae_if : _GEN_76 ? _slots_21_io_out_uop_xcpt_ae_if : _slots_20_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_78 ? _slots_23_io_out_uop_xcpt_ma_if : _GEN_77 ? _slots_22_io_out_uop_xcpt_ma_if : _GEN_76 ? _slots_21_io_out_uop_xcpt_ma_if : _slots_20_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_78 ? _slots_23_io_out_uop_bp_debug_if : _GEN_77 ? _slots_22_io_out_uop_bp_debug_if : _GEN_76 ? _slots_21_io_out_uop_bp_debug_if : _slots_20_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_78 ? _slots_23_io_out_uop_bp_xcpt_if : _GEN_77 ? _slots_22_io_out_uop_bp_xcpt_if : _GEN_76 ? _slots_21_io_out_uop_bp_xcpt_if : _slots_20_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_78 ? _slots_23_io_out_uop_debug_fsrc : _GEN_77 ? _slots_22_io_out_uop_debug_fsrc : _GEN_76 ? _slots_21_io_out_uop_debug_fsrc : _slots_20_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_78 ? _slots_23_io_out_uop_debug_tsrc : _GEN_77 ? _slots_22_io_out_uop_debug_tsrc : _GEN_76 ? _slots_21_io_out_uop_debug_tsrc : _slots_20_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_19_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_19_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_19_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_19_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_19_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_19_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_19_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_19_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_19_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_19_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_19_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_19_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_19_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_19_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_19_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_19_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_19_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_19_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_19_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_19_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_19_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_19_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_19_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_19_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_19_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_19_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_19_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_19_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_19_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_19_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_19_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_19_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_19_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_19_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_19_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_19_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_19_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_19_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_19_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_19_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_19_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_19_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_19_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_19_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_19_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_19_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_19_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_19_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_19_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_19_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_19_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_19_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_19_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_19_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_19_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_19_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_19_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_19_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_19_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_19_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_19_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_19_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_19_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_19_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_19_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_19_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_19_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_19_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_19_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_19_io_uop_uopc),
    .io_uop_inst                    (_slots_19_io_uop_inst),
    .io_uop_debug_inst              (_slots_19_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_19_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_19_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_19_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_19_io_uop_fu_code),
    .io_uop_iw_state                (_slots_19_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_19_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_19_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_19_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_19_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_19_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_19_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_19_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_19_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_19_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_19_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_19_io_uop_pc_lob),
    .io_uop_taken                   (_slots_19_io_uop_taken),
    .io_uop_imm_packed              (_slots_19_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_19_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_19_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_19_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_19_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_19_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_19_io_uop_pdst),
    .io_uop_prs1                    (_slots_19_io_uop_prs1),
    .io_uop_prs2                    (_slots_19_io_uop_prs2),
    .io_uop_prs3                    (_slots_19_io_uop_prs3),
    .io_uop_ppred                   (_slots_19_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_19_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_19_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_19_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_19_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_19_io_uop_stale_pdst),
    .io_uop_exception               (_slots_19_io_uop_exception),
    .io_uop_exc_cause               (_slots_19_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_19_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_19_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_19_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_19_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_19_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_19_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_19_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_19_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_19_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_19_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_19_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_19_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_19_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_19_io_uop_ldst),
    .io_uop_lrs1                    (_slots_19_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_19_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_19_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_19_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_19_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_19_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_19_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_19_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_19_io_uop_fp_val),
    .io_uop_fp_single               (_slots_19_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_19_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_19_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_19_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_19_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_19_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_19_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_19_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_20 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_20_io_valid),
    .io_will_be_valid               (_slots_20_io_will_be_valid),
    .io_request                     (_slots_20_io_request),
    .io_grant                       (issue_slots_20_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_19),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_20_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_81 ? _slots_24_io_out_uop_uopc : _GEN_80 ? _slots_23_io_out_uop_uopc : _GEN_79 ? _slots_22_io_out_uop_uopc : _slots_21_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_81 ? _slots_24_io_out_uop_inst : _GEN_80 ? _slots_23_io_out_uop_inst : _GEN_79 ? _slots_22_io_out_uop_inst : _slots_21_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_81 ? _slots_24_io_out_uop_debug_inst : _GEN_80 ? _slots_23_io_out_uop_debug_inst : _GEN_79 ? _slots_22_io_out_uop_debug_inst : _slots_21_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_81 ? _slots_24_io_out_uop_is_rvc : _GEN_80 ? _slots_23_io_out_uop_is_rvc : _GEN_79 ? _slots_22_io_out_uop_is_rvc : _slots_21_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_81 ? _slots_24_io_out_uop_debug_pc : _GEN_80 ? _slots_23_io_out_uop_debug_pc : _GEN_79 ? _slots_22_io_out_uop_debug_pc : _slots_21_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_81 ? _slots_24_io_out_uop_iq_type : _GEN_80 ? _slots_23_io_out_uop_iq_type : _GEN_79 ? _slots_22_io_out_uop_iq_type : _slots_21_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_81 ? _slots_24_io_out_uop_fu_code : _GEN_80 ? _slots_23_io_out_uop_fu_code : _GEN_79 ? _slots_22_io_out_uop_fu_code : _slots_21_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_81 ? _slots_24_io_out_uop_iw_state : _GEN_80 ? _slots_23_io_out_uop_iw_state : _GEN_79 ? _slots_22_io_out_uop_iw_state : _slots_21_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_81 ? _slots_24_io_out_uop_iw_p1_poisoned : _GEN_80 ? _slots_23_io_out_uop_iw_p1_poisoned : _GEN_79 ? _slots_22_io_out_uop_iw_p1_poisoned : _slots_21_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_81 ? _slots_24_io_out_uop_iw_p2_poisoned : _GEN_80 ? _slots_23_io_out_uop_iw_p2_poisoned : _GEN_79 ? _slots_22_io_out_uop_iw_p2_poisoned : _slots_21_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_81 ? _slots_24_io_out_uop_is_br : _GEN_80 ? _slots_23_io_out_uop_is_br : _GEN_79 ? _slots_22_io_out_uop_is_br : _slots_21_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_81 ? _slots_24_io_out_uop_is_jalr : _GEN_80 ? _slots_23_io_out_uop_is_jalr : _GEN_79 ? _slots_22_io_out_uop_is_jalr : _slots_21_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_81 ? _slots_24_io_out_uop_is_jal : _GEN_80 ? _slots_23_io_out_uop_is_jal : _GEN_79 ? _slots_22_io_out_uop_is_jal : _slots_21_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_81 ? _slots_24_io_out_uop_is_sfb : _GEN_80 ? _slots_23_io_out_uop_is_sfb : _GEN_79 ? _slots_22_io_out_uop_is_sfb : _slots_21_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_81 ? _slots_24_io_out_uop_br_mask : _GEN_80 ? _slots_23_io_out_uop_br_mask : _GEN_79 ? _slots_22_io_out_uop_br_mask : _slots_21_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_81 ? _slots_24_io_out_uop_br_tag : _GEN_80 ? _slots_23_io_out_uop_br_tag : _GEN_79 ? _slots_22_io_out_uop_br_tag : _slots_21_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_81 ? _slots_24_io_out_uop_ftq_idx : _GEN_80 ? _slots_23_io_out_uop_ftq_idx : _GEN_79 ? _slots_22_io_out_uop_ftq_idx : _slots_21_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_81 ? _slots_24_io_out_uop_edge_inst : _GEN_80 ? _slots_23_io_out_uop_edge_inst : _GEN_79 ? _slots_22_io_out_uop_edge_inst : _slots_21_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_81 ? _slots_24_io_out_uop_pc_lob : _GEN_80 ? _slots_23_io_out_uop_pc_lob : _GEN_79 ? _slots_22_io_out_uop_pc_lob : _slots_21_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_81 ? _slots_24_io_out_uop_taken : _GEN_80 ? _slots_23_io_out_uop_taken : _GEN_79 ? _slots_22_io_out_uop_taken : _slots_21_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_81 ? _slots_24_io_out_uop_imm_packed : _GEN_80 ? _slots_23_io_out_uop_imm_packed : _GEN_79 ? _slots_22_io_out_uop_imm_packed : _slots_21_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_81 ? _slots_24_io_out_uop_csr_addr : _GEN_80 ? _slots_23_io_out_uop_csr_addr : _GEN_79 ? _slots_22_io_out_uop_csr_addr : _slots_21_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_81 ? _slots_24_io_out_uop_rob_idx : _GEN_80 ? _slots_23_io_out_uop_rob_idx : _GEN_79 ? _slots_22_io_out_uop_rob_idx : _slots_21_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_81 ? _slots_24_io_out_uop_ldq_idx : _GEN_80 ? _slots_23_io_out_uop_ldq_idx : _GEN_79 ? _slots_22_io_out_uop_ldq_idx : _slots_21_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_81 ? _slots_24_io_out_uop_stq_idx : _GEN_80 ? _slots_23_io_out_uop_stq_idx : _GEN_79 ? _slots_22_io_out_uop_stq_idx : _slots_21_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_81 ? _slots_24_io_out_uop_rxq_idx : _GEN_80 ? _slots_23_io_out_uop_rxq_idx : _GEN_79 ? _slots_22_io_out_uop_rxq_idx : _slots_21_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_81 ? _slots_24_io_out_uop_pdst : _GEN_80 ? _slots_23_io_out_uop_pdst : _GEN_79 ? _slots_22_io_out_uop_pdst : _slots_21_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_81 ? _slots_24_io_out_uop_prs1 : _GEN_80 ? _slots_23_io_out_uop_prs1 : _GEN_79 ? _slots_22_io_out_uop_prs1 : _slots_21_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_81 ? _slots_24_io_out_uop_prs2 : _GEN_80 ? _slots_23_io_out_uop_prs2 : _GEN_79 ? _slots_22_io_out_uop_prs2 : _slots_21_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_81 ? _slots_24_io_out_uop_prs3 : _GEN_80 ? _slots_23_io_out_uop_prs3 : _GEN_79 ? _slots_22_io_out_uop_prs3 : _slots_21_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_81 ? _slots_24_io_out_uop_ppred : _GEN_80 ? _slots_23_io_out_uop_ppred : _GEN_79 ? _slots_22_io_out_uop_ppred : _slots_21_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_81 ? _slots_24_io_out_uop_prs1_busy : _GEN_80 ? _slots_23_io_out_uop_prs1_busy : _GEN_79 ? _slots_22_io_out_uop_prs1_busy : _slots_21_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_81 ? _slots_24_io_out_uop_prs2_busy : _GEN_80 ? _slots_23_io_out_uop_prs2_busy : _GEN_79 ? _slots_22_io_out_uop_prs2_busy : _slots_21_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_81 ? _slots_24_io_out_uop_prs3_busy : _GEN_80 ? _slots_23_io_out_uop_prs3_busy : _GEN_79 ? _slots_22_io_out_uop_prs3_busy : _slots_21_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_81 ? _slots_24_io_out_uop_ppred_busy : _GEN_80 ? _slots_23_io_out_uop_ppred_busy : _GEN_79 ? _slots_22_io_out_uop_ppred_busy : _slots_21_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_81 ? _slots_24_io_out_uop_stale_pdst : _GEN_80 ? _slots_23_io_out_uop_stale_pdst : _GEN_79 ? _slots_22_io_out_uop_stale_pdst : _slots_21_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_81 ? _slots_24_io_out_uop_exception : _GEN_80 ? _slots_23_io_out_uop_exception : _GEN_79 ? _slots_22_io_out_uop_exception : _slots_21_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_81 ? _slots_24_io_out_uop_exc_cause : _GEN_80 ? _slots_23_io_out_uop_exc_cause : _GEN_79 ? _slots_22_io_out_uop_exc_cause : _slots_21_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_81 ? _slots_24_io_out_uop_bypassable : _GEN_80 ? _slots_23_io_out_uop_bypassable : _GEN_79 ? _slots_22_io_out_uop_bypassable : _slots_21_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_81 ? _slots_24_io_out_uop_mem_cmd : _GEN_80 ? _slots_23_io_out_uop_mem_cmd : _GEN_79 ? _slots_22_io_out_uop_mem_cmd : _slots_21_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_81 ? _slots_24_io_out_uop_mem_size : _GEN_80 ? _slots_23_io_out_uop_mem_size : _GEN_79 ? _slots_22_io_out_uop_mem_size : _slots_21_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_81 ? _slots_24_io_out_uop_mem_signed : _GEN_80 ? _slots_23_io_out_uop_mem_signed : _GEN_79 ? _slots_22_io_out_uop_mem_signed : _slots_21_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_81 ? _slots_24_io_out_uop_is_fence : _GEN_80 ? _slots_23_io_out_uop_is_fence : _GEN_79 ? _slots_22_io_out_uop_is_fence : _slots_21_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_81 ? _slots_24_io_out_uop_is_fencei : _GEN_80 ? _slots_23_io_out_uop_is_fencei : _GEN_79 ? _slots_22_io_out_uop_is_fencei : _slots_21_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_81 ? _slots_24_io_out_uop_is_amo : _GEN_80 ? _slots_23_io_out_uop_is_amo : _GEN_79 ? _slots_22_io_out_uop_is_amo : _slots_21_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_81 ? _slots_24_io_out_uop_uses_ldq : _GEN_80 ? _slots_23_io_out_uop_uses_ldq : _GEN_79 ? _slots_22_io_out_uop_uses_ldq : _slots_21_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_81 ? _slots_24_io_out_uop_uses_stq : _GEN_80 ? _slots_23_io_out_uop_uses_stq : _GEN_79 ? _slots_22_io_out_uop_uses_stq : _slots_21_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_81 ? _slots_24_io_out_uop_is_sys_pc2epc : _GEN_80 ? _slots_23_io_out_uop_is_sys_pc2epc : _GEN_79 ? _slots_22_io_out_uop_is_sys_pc2epc : _slots_21_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_81 ? _slots_24_io_out_uop_is_unique : _GEN_80 ? _slots_23_io_out_uop_is_unique : _GEN_79 ? _slots_22_io_out_uop_is_unique : _slots_21_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_81 ? _slots_24_io_out_uop_flush_on_commit : _GEN_80 ? _slots_23_io_out_uop_flush_on_commit : _GEN_79 ? _slots_22_io_out_uop_flush_on_commit : _slots_21_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_81 ? _slots_24_io_out_uop_ldst_is_rs1 : _GEN_80 ? _slots_23_io_out_uop_ldst_is_rs1 : _GEN_79 ? _slots_22_io_out_uop_ldst_is_rs1 : _slots_21_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_81 ? _slots_24_io_out_uop_ldst : _GEN_80 ? _slots_23_io_out_uop_ldst : _GEN_79 ? _slots_22_io_out_uop_ldst : _slots_21_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_81 ? _slots_24_io_out_uop_lrs1 : _GEN_80 ? _slots_23_io_out_uop_lrs1 : _GEN_79 ? _slots_22_io_out_uop_lrs1 : _slots_21_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_81 ? _slots_24_io_out_uop_lrs2 : _GEN_80 ? _slots_23_io_out_uop_lrs2 : _GEN_79 ? _slots_22_io_out_uop_lrs2 : _slots_21_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_81 ? _slots_24_io_out_uop_lrs3 : _GEN_80 ? _slots_23_io_out_uop_lrs3 : _GEN_79 ? _slots_22_io_out_uop_lrs3 : _slots_21_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_81 ? _slots_24_io_out_uop_ldst_val : _GEN_80 ? _slots_23_io_out_uop_ldst_val : _GEN_79 ? _slots_22_io_out_uop_ldst_val : _slots_21_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_81 ? _slots_24_io_out_uop_dst_rtype : _GEN_80 ? _slots_23_io_out_uop_dst_rtype : _GEN_79 ? _slots_22_io_out_uop_dst_rtype : _slots_21_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_81 ? _slots_24_io_out_uop_lrs1_rtype : _GEN_80 ? _slots_23_io_out_uop_lrs1_rtype : _GEN_79 ? _slots_22_io_out_uop_lrs1_rtype : _slots_21_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_81 ? _slots_24_io_out_uop_lrs2_rtype : _GEN_80 ? _slots_23_io_out_uop_lrs2_rtype : _GEN_79 ? _slots_22_io_out_uop_lrs2_rtype : _slots_21_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_81 ? _slots_24_io_out_uop_frs3_en : _GEN_80 ? _slots_23_io_out_uop_frs3_en : _GEN_79 ? _slots_22_io_out_uop_frs3_en : _slots_21_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_81 ? _slots_24_io_out_uop_fp_val : _GEN_80 ? _slots_23_io_out_uop_fp_val : _GEN_79 ? _slots_22_io_out_uop_fp_val : _slots_21_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_81 ? _slots_24_io_out_uop_fp_single : _GEN_80 ? _slots_23_io_out_uop_fp_single : _GEN_79 ? _slots_22_io_out_uop_fp_single : _slots_21_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_81 ? _slots_24_io_out_uop_xcpt_pf_if : _GEN_80 ? _slots_23_io_out_uop_xcpt_pf_if : _GEN_79 ? _slots_22_io_out_uop_xcpt_pf_if : _slots_21_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_81 ? _slots_24_io_out_uop_xcpt_ae_if : _GEN_80 ? _slots_23_io_out_uop_xcpt_ae_if : _GEN_79 ? _slots_22_io_out_uop_xcpt_ae_if : _slots_21_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_81 ? _slots_24_io_out_uop_xcpt_ma_if : _GEN_80 ? _slots_23_io_out_uop_xcpt_ma_if : _GEN_79 ? _slots_22_io_out_uop_xcpt_ma_if : _slots_21_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_81 ? _slots_24_io_out_uop_bp_debug_if : _GEN_80 ? _slots_23_io_out_uop_bp_debug_if : _GEN_79 ? _slots_22_io_out_uop_bp_debug_if : _slots_21_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_81 ? _slots_24_io_out_uop_bp_xcpt_if : _GEN_80 ? _slots_23_io_out_uop_bp_xcpt_if : _GEN_79 ? _slots_22_io_out_uop_bp_xcpt_if : _slots_21_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_81 ? _slots_24_io_out_uop_debug_fsrc : _GEN_80 ? _slots_23_io_out_uop_debug_fsrc : _GEN_79 ? _slots_22_io_out_uop_debug_fsrc : _slots_21_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_81 ? _slots_24_io_out_uop_debug_tsrc : _GEN_80 ? _slots_23_io_out_uop_debug_tsrc : _GEN_79 ? _slots_22_io_out_uop_debug_tsrc : _slots_21_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_20_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_20_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_20_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_20_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_20_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_20_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_20_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_20_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_20_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_20_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_20_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_20_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_20_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_20_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_20_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_20_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_20_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_20_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_20_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_20_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_20_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_20_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_20_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_20_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_20_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_20_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_20_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_20_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_20_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_20_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_20_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_20_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_20_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_20_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_20_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_20_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_20_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_20_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_20_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_20_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_20_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_20_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_20_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_20_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_20_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_20_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_20_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_20_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_20_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_20_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_20_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_20_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_20_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_20_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_20_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_20_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_20_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_20_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_20_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_20_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_20_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_20_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_20_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_20_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_20_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_20_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_20_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_20_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_20_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_20_io_uop_uopc),
    .io_uop_inst                    (_slots_20_io_uop_inst),
    .io_uop_debug_inst              (_slots_20_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_20_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_20_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_20_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_20_io_uop_fu_code),
    .io_uop_iw_state                (_slots_20_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_20_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_20_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_20_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_20_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_20_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_20_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_20_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_20_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_20_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_20_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_20_io_uop_pc_lob),
    .io_uop_taken                   (_slots_20_io_uop_taken),
    .io_uop_imm_packed              (_slots_20_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_20_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_20_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_20_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_20_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_20_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_20_io_uop_pdst),
    .io_uop_prs1                    (_slots_20_io_uop_prs1),
    .io_uop_prs2                    (_slots_20_io_uop_prs2),
    .io_uop_prs3                    (_slots_20_io_uop_prs3),
    .io_uop_ppred                   (_slots_20_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_20_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_20_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_20_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_20_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_20_io_uop_stale_pdst),
    .io_uop_exception               (_slots_20_io_uop_exception),
    .io_uop_exc_cause               (_slots_20_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_20_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_20_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_20_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_20_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_20_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_20_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_20_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_20_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_20_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_20_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_20_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_20_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_20_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_20_io_uop_ldst),
    .io_uop_lrs1                    (_slots_20_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_20_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_20_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_20_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_20_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_20_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_20_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_20_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_20_io_uop_fp_val),
    .io_uop_fp_single               (_slots_20_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_20_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_20_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_20_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_20_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_20_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_20_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_20_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_21 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_21_io_valid),
    .io_will_be_valid               (_slots_21_io_will_be_valid),
    .io_request                     (_slots_21_io_request),
    .io_grant                       (issue_slots_21_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_20),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_21_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_84 ? _slots_25_io_out_uop_uopc : _GEN_83 ? _slots_24_io_out_uop_uopc : _GEN_82 ? _slots_23_io_out_uop_uopc : _slots_22_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_84 ? _slots_25_io_out_uop_inst : _GEN_83 ? _slots_24_io_out_uop_inst : _GEN_82 ? _slots_23_io_out_uop_inst : _slots_22_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_84 ? _slots_25_io_out_uop_debug_inst : _GEN_83 ? _slots_24_io_out_uop_debug_inst : _GEN_82 ? _slots_23_io_out_uop_debug_inst : _slots_22_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_84 ? _slots_25_io_out_uop_is_rvc : _GEN_83 ? _slots_24_io_out_uop_is_rvc : _GEN_82 ? _slots_23_io_out_uop_is_rvc : _slots_22_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_84 ? _slots_25_io_out_uop_debug_pc : _GEN_83 ? _slots_24_io_out_uop_debug_pc : _GEN_82 ? _slots_23_io_out_uop_debug_pc : _slots_22_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_84 ? _slots_25_io_out_uop_iq_type : _GEN_83 ? _slots_24_io_out_uop_iq_type : _GEN_82 ? _slots_23_io_out_uop_iq_type : _slots_22_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_84 ? _slots_25_io_out_uop_fu_code : _GEN_83 ? _slots_24_io_out_uop_fu_code : _GEN_82 ? _slots_23_io_out_uop_fu_code : _slots_22_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_84 ? _slots_25_io_out_uop_iw_state : _GEN_83 ? _slots_24_io_out_uop_iw_state : _GEN_82 ? _slots_23_io_out_uop_iw_state : _slots_22_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_84 ? _slots_25_io_out_uop_iw_p1_poisoned : _GEN_83 ? _slots_24_io_out_uop_iw_p1_poisoned : _GEN_82 ? _slots_23_io_out_uop_iw_p1_poisoned : _slots_22_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_84 ? _slots_25_io_out_uop_iw_p2_poisoned : _GEN_83 ? _slots_24_io_out_uop_iw_p2_poisoned : _GEN_82 ? _slots_23_io_out_uop_iw_p2_poisoned : _slots_22_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_84 ? _slots_25_io_out_uop_is_br : _GEN_83 ? _slots_24_io_out_uop_is_br : _GEN_82 ? _slots_23_io_out_uop_is_br : _slots_22_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_84 ? _slots_25_io_out_uop_is_jalr : _GEN_83 ? _slots_24_io_out_uop_is_jalr : _GEN_82 ? _slots_23_io_out_uop_is_jalr : _slots_22_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_84 ? _slots_25_io_out_uop_is_jal : _GEN_83 ? _slots_24_io_out_uop_is_jal : _GEN_82 ? _slots_23_io_out_uop_is_jal : _slots_22_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_84 ? _slots_25_io_out_uop_is_sfb : _GEN_83 ? _slots_24_io_out_uop_is_sfb : _GEN_82 ? _slots_23_io_out_uop_is_sfb : _slots_22_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_84 ? _slots_25_io_out_uop_br_mask : _GEN_83 ? _slots_24_io_out_uop_br_mask : _GEN_82 ? _slots_23_io_out_uop_br_mask : _slots_22_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_84 ? _slots_25_io_out_uop_br_tag : _GEN_83 ? _slots_24_io_out_uop_br_tag : _GEN_82 ? _slots_23_io_out_uop_br_tag : _slots_22_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_84 ? _slots_25_io_out_uop_ftq_idx : _GEN_83 ? _slots_24_io_out_uop_ftq_idx : _GEN_82 ? _slots_23_io_out_uop_ftq_idx : _slots_22_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_84 ? _slots_25_io_out_uop_edge_inst : _GEN_83 ? _slots_24_io_out_uop_edge_inst : _GEN_82 ? _slots_23_io_out_uop_edge_inst : _slots_22_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_84 ? _slots_25_io_out_uop_pc_lob : _GEN_83 ? _slots_24_io_out_uop_pc_lob : _GEN_82 ? _slots_23_io_out_uop_pc_lob : _slots_22_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_84 ? _slots_25_io_out_uop_taken : _GEN_83 ? _slots_24_io_out_uop_taken : _GEN_82 ? _slots_23_io_out_uop_taken : _slots_22_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_84 ? _slots_25_io_out_uop_imm_packed : _GEN_83 ? _slots_24_io_out_uop_imm_packed : _GEN_82 ? _slots_23_io_out_uop_imm_packed : _slots_22_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_84 ? _slots_25_io_out_uop_csr_addr : _GEN_83 ? _slots_24_io_out_uop_csr_addr : _GEN_82 ? _slots_23_io_out_uop_csr_addr : _slots_22_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_84 ? _slots_25_io_out_uop_rob_idx : _GEN_83 ? _slots_24_io_out_uop_rob_idx : _GEN_82 ? _slots_23_io_out_uop_rob_idx : _slots_22_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_84 ? _slots_25_io_out_uop_ldq_idx : _GEN_83 ? _slots_24_io_out_uop_ldq_idx : _GEN_82 ? _slots_23_io_out_uop_ldq_idx : _slots_22_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_84 ? _slots_25_io_out_uop_stq_idx : _GEN_83 ? _slots_24_io_out_uop_stq_idx : _GEN_82 ? _slots_23_io_out_uop_stq_idx : _slots_22_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_84 ? _slots_25_io_out_uop_rxq_idx : _GEN_83 ? _slots_24_io_out_uop_rxq_idx : _GEN_82 ? _slots_23_io_out_uop_rxq_idx : _slots_22_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_84 ? _slots_25_io_out_uop_pdst : _GEN_83 ? _slots_24_io_out_uop_pdst : _GEN_82 ? _slots_23_io_out_uop_pdst : _slots_22_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_84 ? _slots_25_io_out_uop_prs1 : _GEN_83 ? _slots_24_io_out_uop_prs1 : _GEN_82 ? _slots_23_io_out_uop_prs1 : _slots_22_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_84 ? _slots_25_io_out_uop_prs2 : _GEN_83 ? _slots_24_io_out_uop_prs2 : _GEN_82 ? _slots_23_io_out_uop_prs2 : _slots_22_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_84 ? _slots_25_io_out_uop_prs3 : _GEN_83 ? _slots_24_io_out_uop_prs3 : _GEN_82 ? _slots_23_io_out_uop_prs3 : _slots_22_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_84 ? _slots_25_io_out_uop_ppred : _GEN_83 ? _slots_24_io_out_uop_ppred : _GEN_82 ? _slots_23_io_out_uop_ppred : _slots_22_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_84 ? _slots_25_io_out_uop_prs1_busy : _GEN_83 ? _slots_24_io_out_uop_prs1_busy : _GEN_82 ? _slots_23_io_out_uop_prs1_busy : _slots_22_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_84 ? _slots_25_io_out_uop_prs2_busy : _GEN_83 ? _slots_24_io_out_uop_prs2_busy : _GEN_82 ? _slots_23_io_out_uop_prs2_busy : _slots_22_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_84 ? _slots_25_io_out_uop_prs3_busy : _GEN_83 ? _slots_24_io_out_uop_prs3_busy : _GEN_82 ? _slots_23_io_out_uop_prs3_busy : _slots_22_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_84 ? _slots_25_io_out_uop_ppred_busy : _GEN_83 ? _slots_24_io_out_uop_ppred_busy : _GEN_82 ? _slots_23_io_out_uop_ppred_busy : _slots_22_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_84 ? _slots_25_io_out_uop_stale_pdst : _GEN_83 ? _slots_24_io_out_uop_stale_pdst : _GEN_82 ? _slots_23_io_out_uop_stale_pdst : _slots_22_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_84 ? _slots_25_io_out_uop_exception : _GEN_83 ? _slots_24_io_out_uop_exception : _GEN_82 ? _slots_23_io_out_uop_exception : _slots_22_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_84 ? _slots_25_io_out_uop_exc_cause : _GEN_83 ? _slots_24_io_out_uop_exc_cause : _GEN_82 ? _slots_23_io_out_uop_exc_cause : _slots_22_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_84 ? _slots_25_io_out_uop_bypassable : _GEN_83 ? _slots_24_io_out_uop_bypassable : _GEN_82 ? _slots_23_io_out_uop_bypassable : _slots_22_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_84 ? _slots_25_io_out_uop_mem_cmd : _GEN_83 ? _slots_24_io_out_uop_mem_cmd : _GEN_82 ? _slots_23_io_out_uop_mem_cmd : _slots_22_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_84 ? _slots_25_io_out_uop_mem_size : _GEN_83 ? _slots_24_io_out_uop_mem_size : _GEN_82 ? _slots_23_io_out_uop_mem_size : _slots_22_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_84 ? _slots_25_io_out_uop_mem_signed : _GEN_83 ? _slots_24_io_out_uop_mem_signed : _GEN_82 ? _slots_23_io_out_uop_mem_signed : _slots_22_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_84 ? _slots_25_io_out_uop_is_fence : _GEN_83 ? _slots_24_io_out_uop_is_fence : _GEN_82 ? _slots_23_io_out_uop_is_fence : _slots_22_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_84 ? _slots_25_io_out_uop_is_fencei : _GEN_83 ? _slots_24_io_out_uop_is_fencei : _GEN_82 ? _slots_23_io_out_uop_is_fencei : _slots_22_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_84 ? _slots_25_io_out_uop_is_amo : _GEN_83 ? _slots_24_io_out_uop_is_amo : _GEN_82 ? _slots_23_io_out_uop_is_amo : _slots_22_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_84 ? _slots_25_io_out_uop_uses_ldq : _GEN_83 ? _slots_24_io_out_uop_uses_ldq : _GEN_82 ? _slots_23_io_out_uop_uses_ldq : _slots_22_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_84 ? _slots_25_io_out_uop_uses_stq : _GEN_83 ? _slots_24_io_out_uop_uses_stq : _GEN_82 ? _slots_23_io_out_uop_uses_stq : _slots_22_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_84 ? _slots_25_io_out_uop_is_sys_pc2epc : _GEN_83 ? _slots_24_io_out_uop_is_sys_pc2epc : _GEN_82 ? _slots_23_io_out_uop_is_sys_pc2epc : _slots_22_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_84 ? _slots_25_io_out_uop_is_unique : _GEN_83 ? _slots_24_io_out_uop_is_unique : _GEN_82 ? _slots_23_io_out_uop_is_unique : _slots_22_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_84 ? _slots_25_io_out_uop_flush_on_commit : _GEN_83 ? _slots_24_io_out_uop_flush_on_commit : _GEN_82 ? _slots_23_io_out_uop_flush_on_commit : _slots_22_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_84 ? _slots_25_io_out_uop_ldst_is_rs1 : _GEN_83 ? _slots_24_io_out_uop_ldst_is_rs1 : _GEN_82 ? _slots_23_io_out_uop_ldst_is_rs1 : _slots_22_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_84 ? _slots_25_io_out_uop_ldst : _GEN_83 ? _slots_24_io_out_uop_ldst : _GEN_82 ? _slots_23_io_out_uop_ldst : _slots_22_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_84 ? _slots_25_io_out_uop_lrs1 : _GEN_83 ? _slots_24_io_out_uop_lrs1 : _GEN_82 ? _slots_23_io_out_uop_lrs1 : _slots_22_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_84 ? _slots_25_io_out_uop_lrs2 : _GEN_83 ? _slots_24_io_out_uop_lrs2 : _GEN_82 ? _slots_23_io_out_uop_lrs2 : _slots_22_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_84 ? _slots_25_io_out_uop_lrs3 : _GEN_83 ? _slots_24_io_out_uop_lrs3 : _GEN_82 ? _slots_23_io_out_uop_lrs3 : _slots_22_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_84 ? _slots_25_io_out_uop_ldst_val : _GEN_83 ? _slots_24_io_out_uop_ldst_val : _GEN_82 ? _slots_23_io_out_uop_ldst_val : _slots_22_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_84 ? _slots_25_io_out_uop_dst_rtype : _GEN_83 ? _slots_24_io_out_uop_dst_rtype : _GEN_82 ? _slots_23_io_out_uop_dst_rtype : _slots_22_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_84 ? _slots_25_io_out_uop_lrs1_rtype : _GEN_83 ? _slots_24_io_out_uop_lrs1_rtype : _GEN_82 ? _slots_23_io_out_uop_lrs1_rtype : _slots_22_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_84 ? _slots_25_io_out_uop_lrs2_rtype : _GEN_83 ? _slots_24_io_out_uop_lrs2_rtype : _GEN_82 ? _slots_23_io_out_uop_lrs2_rtype : _slots_22_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_84 ? _slots_25_io_out_uop_frs3_en : _GEN_83 ? _slots_24_io_out_uop_frs3_en : _GEN_82 ? _slots_23_io_out_uop_frs3_en : _slots_22_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_84 ? _slots_25_io_out_uop_fp_val : _GEN_83 ? _slots_24_io_out_uop_fp_val : _GEN_82 ? _slots_23_io_out_uop_fp_val : _slots_22_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_84 ? _slots_25_io_out_uop_fp_single : _GEN_83 ? _slots_24_io_out_uop_fp_single : _GEN_82 ? _slots_23_io_out_uop_fp_single : _slots_22_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_84 ? _slots_25_io_out_uop_xcpt_pf_if : _GEN_83 ? _slots_24_io_out_uop_xcpt_pf_if : _GEN_82 ? _slots_23_io_out_uop_xcpt_pf_if : _slots_22_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_84 ? _slots_25_io_out_uop_xcpt_ae_if : _GEN_83 ? _slots_24_io_out_uop_xcpt_ae_if : _GEN_82 ? _slots_23_io_out_uop_xcpt_ae_if : _slots_22_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_84 ? _slots_25_io_out_uop_xcpt_ma_if : _GEN_83 ? _slots_24_io_out_uop_xcpt_ma_if : _GEN_82 ? _slots_23_io_out_uop_xcpt_ma_if : _slots_22_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_84 ? _slots_25_io_out_uop_bp_debug_if : _GEN_83 ? _slots_24_io_out_uop_bp_debug_if : _GEN_82 ? _slots_23_io_out_uop_bp_debug_if : _slots_22_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_84 ? _slots_25_io_out_uop_bp_xcpt_if : _GEN_83 ? _slots_24_io_out_uop_bp_xcpt_if : _GEN_82 ? _slots_23_io_out_uop_bp_xcpt_if : _slots_22_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_84 ? _slots_25_io_out_uop_debug_fsrc : _GEN_83 ? _slots_24_io_out_uop_debug_fsrc : _GEN_82 ? _slots_23_io_out_uop_debug_fsrc : _slots_22_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_84 ? _slots_25_io_out_uop_debug_tsrc : _GEN_83 ? _slots_24_io_out_uop_debug_tsrc : _GEN_82 ? _slots_23_io_out_uop_debug_tsrc : _slots_22_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_21_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_21_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_21_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_21_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_21_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_21_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_21_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_21_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_21_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_21_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_21_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_21_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_21_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_21_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_21_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_21_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_21_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_21_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_21_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_21_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_21_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_21_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_21_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_21_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_21_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_21_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_21_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_21_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_21_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_21_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_21_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_21_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_21_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_21_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_21_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_21_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_21_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_21_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_21_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_21_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_21_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_21_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_21_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_21_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_21_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_21_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_21_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_21_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_21_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_21_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_21_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_21_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_21_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_21_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_21_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_21_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_21_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_21_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_21_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_21_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_21_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_21_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_21_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_21_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_21_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_21_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_21_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_21_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_21_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_21_io_uop_uopc),
    .io_uop_inst                    (_slots_21_io_uop_inst),
    .io_uop_debug_inst              (_slots_21_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_21_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_21_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_21_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_21_io_uop_fu_code),
    .io_uop_iw_state                (_slots_21_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_21_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_21_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_21_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_21_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_21_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_21_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_21_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_21_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_21_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_21_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_21_io_uop_pc_lob),
    .io_uop_taken                   (_slots_21_io_uop_taken),
    .io_uop_imm_packed              (_slots_21_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_21_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_21_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_21_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_21_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_21_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_21_io_uop_pdst),
    .io_uop_prs1                    (_slots_21_io_uop_prs1),
    .io_uop_prs2                    (_slots_21_io_uop_prs2),
    .io_uop_prs3                    (_slots_21_io_uop_prs3),
    .io_uop_ppred                   (_slots_21_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_21_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_21_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_21_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_21_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_21_io_uop_stale_pdst),
    .io_uop_exception               (_slots_21_io_uop_exception),
    .io_uop_exc_cause               (_slots_21_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_21_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_21_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_21_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_21_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_21_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_21_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_21_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_21_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_21_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_21_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_21_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_21_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_21_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_21_io_uop_ldst),
    .io_uop_lrs1                    (_slots_21_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_21_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_21_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_21_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_21_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_21_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_21_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_21_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_21_io_uop_fp_val),
    .io_uop_fp_single               (_slots_21_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_21_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_21_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_21_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_21_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_21_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_21_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_21_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_22 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_22_io_valid),
    .io_will_be_valid               (_slots_22_io_will_be_valid),
    .io_request                     (_slots_22_io_request),
    .io_grant                       (issue_slots_22_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_21),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_22_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_87 ? _slots_26_io_out_uop_uopc : _GEN_86 ? _slots_25_io_out_uop_uopc : _GEN_85 ? _slots_24_io_out_uop_uopc : _slots_23_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_87 ? _slots_26_io_out_uop_inst : _GEN_86 ? _slots_25_io_out_uop_inst : _GEN_85 ? _slots_24_io_out_uop_inst : _slots_23_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_87 ? _slots_26_io_out_uop_debug_inst : _GEN_86 ? _slots_25_io_out_uop_debug_inst : _GEN_85 ? _slots_24_io_out_uop_debug_inst : _slots_23_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_87 ? _slots_26_io_out_uop_is_rvc : _GEN_86 ? _slots_25_io_out_uop_is_rvc : _GEN_85 ? _slots_24_io_out_uop_is_rvc : _slots_23_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_87 ? _slots_26_io_out_uop_debug_pc : _GEN_86 ? _slots_25_io_out_uop_debug_pc : _GEN_85 ? _slots_24_io_out_uop_debug_pc : _slots_23_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_87 ? _slots_26_io_out_uop_iq_type : _GEN_86 ? _slots_25_io_out_uop_iq_type : _GEN_85 ? _slots_24_io_out_uop_iq_type : _slots_23_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_87 ? _slots_26_io_out_uop_fu_code : _GEN_86 ? _slots_25_io_out_uop_fu_code : _GEN_85 ? _slots_24_io_out_uop_fu_code : _slots_23_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_87 ? _slots_26_io_out_uop_iw_state : _GEN_86 ? _slots_25_io_out_uop_iw_state : _GEN_85 ? _slots_24_io_out_uop_iw_state : _slots_23_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_87 ? _slots_26_io_out_uop_iw_p1_poisoned : _GEN_86 ? _slots_25_io_out_uop_iw_p1_poisoned : _GEN_85 ? _slots_24_io_out_uop_iw_p1_poisoned : _slots_23_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_87 ? _slots_26_io_out_uop_iw_p2_poisoned : _GEN_86 ? _slots_25_io_out_uop_iw_p2_poisoned : _GEN_85 ? _slots_24_io_out_uop_iw_p2_poisoned : _slots_23_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_87 ? _slots_26_io_out_uop_is_br : _GEN_86 ? _slots_25_io_out_uop_is_br : _GEN_85 ? _slots_24_io_out_uop_is_br : _slots_23_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_87 ? _slots_26_io_out_uop_is_jalr : _GEN_86 ? _slots_25_io_out_uop_is_jalr : _GEN_85 ? _slots_24_io_out_uop_is_jalr : _slots_23_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_87 ? _slots_26_io_out_uop_is_jal : _GEN_86 ? _slots_25_io_out_uop_is_jal : _GEN_85 ? _slots_24_io_out_uop_is_jal : _slots_23_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_87 ? _slots_26_io_out_uop_is_sfb : _GEN_86 ? _slots_25_io_out_uop_is_sfb : _GEN_85 ? _slots_24_io_out_uop_is_sfb : _slots_23_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_87 ? _slots_26_io_out_uop_br_mask : _GEN_86 ? _slots_25_io_out_uop_br_mask : _GEN_85 ? _slots_24_io_out_uop_br_mask : _slots_23_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_87 ? _slots_26_io_out_uop_br_tag : _GEN_86 ? _slots_25_io_out_uop_br_tag : _GEN_85 ? _slots_24_io_out_uop_br_tag : _slots_23_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_87 ? _slots_26_io_out_uop_ftq_idx : _GEN_86 ? _slots_25_io_out_uop_ftq_idx : _GEN_85 ? _slots_24_io_out_uop_ftq_idx : _slots_23_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_87 ? _slots_26_io_out_uop_edge_inst : _GEN_86 ? _slots_25_io_out_uop_edge_inst : _GEN_85 ? _slots_24_io_out_uop_edge_inst : _slots_23_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_87 ? _slots_26_io_out_uop_pc_lob : _GEN_86 ? _slots_25_io_out_uop_pc_lob : _GEN_85 ? _slots_24_io_out_uop_pc_lob : _slots_23_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_87 ? _slots_26_io_out_uop_taken : _GEN_86 ? _slots_25_io_out_uop_taken : _GEN_85 ? _slots_24_io_out_uop_taken : _slots_23_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_87 ? _slots_26_io_out_uop_imm_packed : _GEN_86 ? _slots_25_io_out_uop_imm_packed : _GEN_85 ? _slots_24_io_out_uop_imm_packed : _slots_23_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_87 ? _slots_26_io_out_uop_csr_addr : _GEN_86 ? _slots_25_io_out_uop_csr_addr : _GEN_85 ? _slots_24_io_out_uop_csr_addr : _slots_23_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_87 ? _slots_26_io_out_uop_rob_idx : _GEN_86 ? _slots_25_io_out_uop_rob_idx : _GEN_85 ? _slots_24_io_out_uop_rob_idx : _slots_23_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_87 ? _slots_26_io_out_uop_ldq_idx : _GEN_86 ? _slots_25_io_out_uop_ldq_idx : _GEN_85 ? _slots_24_io_out_uop_ldq_idx : _slots_23_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_87 ? _slots_26_io_out_uop_stq_idx : _GEN_86 ? _slots_25_io_out_uop_stq_idx : _GEN_85 ? _slots_24_io_out_uop_stq_idx : _slots_23_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_87 ? _slots_26_io_out_uop_rxq_idx : _GEN_86 ? _slots_25_io_out_uop_rxq_idx : _GEN_85 ? _slots_24_io_out_uop_rxq_idx : _slots_23_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_87 ? _slots_26_io_out_uop_pdst : _GEN_86 ? _slots_25_io_out_uop_pdst : _GEN_85 ? _slots_24_io_out_uop_pdst : _slots_23_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_87 ? _slots_26_io_out_uop_prs1 : _GEN_86 ? _slots_25_io_out_uop_prs1 : _GEN_85 ? _slots_24_io_out_uop_prs1 : _slots_23_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_87 ? _slots_26_io_out_uop_prs2 : _GEN_86 ? _slots_25_io_out_uop_prs2 : _GEN_85 ? _slots_24_io_out_uop_prs2 : _slots_23_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_87 ? _slots_26_io_out_uop_prs3 : _GEN_86 ? _slots_25_io_out_uop_prs3 : _GEN_85 ? _slots_24_io_out_uop_prs3 : _slots_23_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_87 ? _slots_26_io_out_uop_ppred : _GEN_86 ? _slots_25_io_out_uop_ppred : _GEN_85 ? _slots_24_io_out_uop_ppred : _slots_23_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_87 ? _slots_26_io_out_uop_prs1_busy : _GEN_86 ? _slots_25_io_out_uop_prs1_busy : _GEN_85 ? _slots_24_io_out_uop_prs1_busy : _slots_23_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_87 ? _slots_26_io_out_uop_prs2_busy : _GEN_86 ? _slots_25_io_out_uop_prs2_busy : _GEN_85 ? _slots_24_io_out_uop_prs2_busy : _slots_23_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_87 ? _slots_26_io_out_uop_prs3_busy : _GEN_86 ? _slots_25_io_out_uop_prs3_busy : _GEN_85 ? _slots_24_io_out_uop_prs3_busy : _slots_23_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_87 ? _slots_26_io_out_uop_ppred_busy : _GEN_86 ? _slots_25_io_out_uop_ppred_busy : _GEN_85 ? _slots_24_io_out_uop_ppred_busy : _slots_23_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_87 ? _slots_26_io_out_uop_stale_pdst : _GEN_86 ? _slots_25_io_out_uop_stale_pdst : _GEN_85 ? _slots_24_io_out_uop_stale_pdst : _slots_23_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_87 ? _slots_26_io_out_uop_exception : _GEN_86 ? _slots_25_io_out_uop_exception : _GEN_85 ? _slots_24_io_out_uop_exception : _slots_23_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_87 ? _slots_26_io_out_uop_exc_cause : _GEN_86 ? _slots_25_io_out_uop_exc_cause : _GEN_85 ? _slots_24_io_out_uop_exc_cause : _slots_23_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_87 ? _slots_26_io_out_uop_bypassable : _GEN_86 ? _slots_25_io_out_uop_bypassable : _GEN_85 ? _slots_24_io_out_uop_bypassable : _slots_23_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_87 ? _slots_26_io_out_uop_mem_cmd : _GEN_86 ? _slots_25_io_out_uop_mem_cmd : _GEN_85 ? _slots_24_io_out_uop_mem_cmd : _slots_23_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_87 ? _slots_26_io_out_uop_mem_size : _GEN_86 ? _slots_25_io_out_uop_mem_size : _GEN_85 ? _slots_24_io_out_uop_mem_size : _slots_23_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_87 ? _slots_26_io_out_uop_mem_signed : _GEN_86 ? _slots_25_io_out_uop_mem_signed : _GEN_85 ? _slots_24_io_out_uop_mem_signed : _slots_23_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_87 ? _slots_26_io_out_uop_is_fence : _GEN_86 ? _slots_25_io_out_uop_is_fence : _GEN_85 ? _slots_24_io_out_uop_is_fence : _slots_23_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_87 ? _slots_26_io_out_uop_is_fencei : _GEN_86 ? _slots_25_io_out_uop_is_fencei : _GEN_85 ? _slots_24_io_out_uop_is_fencei : _slots_23_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_87 ? _slots_26_io_out_uop_is_amo : _GEN_86 ? _slots_25_io_out_uop_is_amo : _GEN_85 ? _slots_24_io_out_uop_is_amo : _slots_23_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_87 ? _slots_26_io_out_uop_uses_ldq : _GEN_86 ? _slots_25_io_out_uop_uses_ldq : _GEN_85 ? _slots_24_io_out_uop_uses_ldq : _slots_23_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_87 ? _slots_26_io_out_uop_uses_stq : _GEN_86 ? _slots_25_io_out_uop_uses_stq : _GEN_85 ? _slots_24_io_out_uop_uses_stq : _slots_23_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_87 ? _slots_26_io_out_uop_is_sys_pc2epc : _GEN_86 ? _slots_25_io_out_uop_is_sys_pc2epc : _GEN_85 ? _slots_24_io_out_uop_is_sys_pc2epc : _slots_23_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_87 ? _slots_26_io_out_uop_is_unique : _GEN_86 ? _slots_25_io_out_uop_is_unique : _GEN_85 ? _slots_24_io_out_uop_is_unique : _slots_23_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_87 ? _slots_26_io_out_uop_flush_on_commit : _GEN_86 ? _slots_25_io_out_uop_flush_on_commit : _GEN_85 ? _slots_24_io_out_uop_flush_on_commit : _slots_23_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_87 ? _slots_26_io_out_uop_ldst_is_rs1 : _GEN_86 ? _slots_25_io_out_uop_ldst_is_rs1 : _GEN_85 ? _slots_24_io_out_uop_ldst_is_rs1 : _slots_23_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_87 ? _slots_26_io_out_uop_ldst : _GEN_86 ? _slots_25_io_out_uop_ldst : _GEN_85 ? _slots_24_io_out_uop_ldst : _slots_23_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_87 ? _slots_26_io_out_uop_lrs1 : _GEN_86 ? _slots_25_io_out_uop_lrs1 : _GEN_85 ? _slots_24_io_out_uop_lrs1 : _slots_23_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_87 ? _slots_26_io_out_uop_lrs2 : _GEN_86 ? _slots_25_io_out_uop_lrs2 : _GEN_85 ? _slots_24_io_out_uop_lrs2 : _slots_23_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_87 ? _slots_26_io_out_uop_lrs3 : _GEN_86 ? _slots_25_io_out_uop_lrs3 : _GEN_85 ? _slots_24_io_out_uop_lrs3 : _slots_23_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_87 ? _slots_26_io_out_uop_ldst_val : _GEN_86 ? _slots_25_io_out_uop_ldst_val : _GEN_85 ? _slots_24_io_out_uop_ldst_val : _slots_23_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_87 ? _slots_26_io_out_uop_dst_rtype : _GEN_86 ? _slots_25_io_out_uop_dst_rtype : _GEN_85 ? _slots_24_io_out_uop_dst_rtype : _slots_23_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_87 ? _slots_26_io_out_uop_lrs1_rtype : _GEN_86 ? _slots_25_io_out_uop_lrs1_rtype : _GEN_85 ? _slots_24_io_out_uop_lrs1_rtype : _slots_23_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_87 ? _slots_26_io_out_uop_lrs2_rtype : _GEN_86 ? _slots_25_io_out_uop_lrs2_rtype : _GEN_85 ? _slots_24_io_out_uop_lrs2_rtype : _slots_23_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_87 ? _slots_26_io_out_uop_frs3_en : _GEN_86 ? _slots_25_io_out_uop_frs3_en : _GEN_85 ? _slots_24_io_out_uop_frs3_en : _slots_23_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_87 ? _slots_26_io_out_uop_fp_val : _GEN_86 ? _slots_25_io_out_uop_fp_val : _GEN_85 ? _slots_24_io_out_uop_fp_val : _slots_23_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_87 ? _slots_26_io_out_uop_fp_single : _GEN_86 ? _slots_25_io_out_uop_fp_single : _GEN_85 ? _slots_24_io_out_uop_fp_single : _slots_23_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_87 ? _slots_26_io_out_uop_xcpt_pf_if : _GEN_86 ? _slots_25_io_out_uop_xcpt_pf_if : _GEN_85 ? _slots_24_io_out_uop_xcpt_pf_if : _slots_23_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_87 ? _slots_26_io_out_uop_xcpt_ae_if : _GEN_86 ? _slots_25_io_out_uop_xcpt_ae_if : _GEN_85 ? _slots_24_io_out_uop_xcpt_ae_if : _slots_23_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_87 ? _slots_26_io_out_uop_xcpt_ma_if : _GEN_86 ? _slots_25_io_out_uop_xcpt_ma_if : _GEN_85 ? _slots_24_io_out_uop_xcpt_ma_if : _slots_23_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_87 ? _slots_26_io_out_uop_bp_debug_if : _GEN_86 ? _slots_25_io_out_uop_bp_debug_if : _GEN_85 ? _slots_24_io_out_uop_bp_debug_if : _slots_23_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_87 ? _slots_26_io_out_uop_bp_xcpt_if : _GEN_86 ? _slots_25_io_out_uop_bp_xcpt_if : _GEN_85 ? _slots_24_io_out_uop_bp_xcpt_if : _slots_23_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_87 ? _slots_26_io_out_uop_debug_fsrc : _GEN_86 ? _slots_25_io_out_uop_debug_fsrc : _GEN_85 ? _slots_24_io_out_uop_debug_fsrc : _slots_23_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_87 ? _slots_26_io_out_uop_debug_tsrc : _GEN_86 ? _slots_25_io_out_uop_debug_tsrc : _GEN_85 ? _slots_24_io_out_uop_debug_tsrc : _slots_23_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_22_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_22_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_22_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_22_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_22_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_22_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_22_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_22_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_22_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_22_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_22_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_22_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_22_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_22_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_22_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_22_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_22_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_22_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_22_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_22_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_22_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_22_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_22_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_22_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_22_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_22_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_22_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_22_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_22_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_22_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_22_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_22_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_22_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_22_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_22_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_22_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_22_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_22_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_22_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_22_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_22_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_22_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_22_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_22_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_22_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_22_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_22_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_22_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_22_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_22_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_22_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_22_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_22_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_22_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_22_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_22_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_22_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_22_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_22_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_22_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_22_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_22_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_22_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_22_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_22_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_22_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_22_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_22_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_22_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_22_io_uop_uopc),
    .io_uop_inst                    (_slots_22_io_uop_inst),
    .io_uop_debug_inst              (_slots_22_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_22_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_22_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_22_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_22_io_uop_fu_code),
    .io_uop_iw_state                (_slots_22_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_22_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_22_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_22_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_22_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_22_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_22_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_22_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_22_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_22_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_22_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_22_io_uop_pc_lob),
    .io_uop_taken                   (_slots_22_io_uop_taken),
    .io_uop_imm_packed              (_slots_22_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_22_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_22_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_22_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_22_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_22_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_22_io_uop_pdst),
    .io_uop_prs1                    (_slots_22_io_uop_prs1),
    .io_uop_prs2                    (_slots_22_io_uop_prs2),
    .io_uop_prs3                    (_slots_22_io_uop_prs3),
    .io_uop_ppred                   (_slots_22_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_22_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_22_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_22_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_22_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_22_io_uop_stale_pdst),
    .io_uop_exception               (_slots_22_io_uop_exception),
    .io_uop_exc_cause               (_slots_22_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_22_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_22_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_22_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_22_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_22_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_22_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_22_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_22_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_22_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_22_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_22_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_22_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_22_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_22_io_uop_ldst),
    .io_uop_lrs1                    (_slots_22_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_22_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_22_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_22_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_22_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_22_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_22_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_22_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_22_io_uop_fp_val),
    .io_uop_fp_single               (_slots_22_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_22_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_22_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_22_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_22_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_22_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_22_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_22_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_23 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_23_io_valid),
    .io_will_be_valid               (_slots_23_io_will_be_valid),
    .io_request                     (_slots_23_io_request),
    .io_grant                       (issue_slots_23_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_22),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_23_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_90 ? _slots_27_io_out_uop_uopc : _GEN_89 ? _slots_26_io_out_uop_uopc : _GEN_88 ? _slots_25_io_out_uop_uopc : _slots_24_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_90 ? _slots_27_io_out_uop_inst : _GEN_89 ? _slots_26_io_out_uop_inst : _GEN_88 ? _slots_25_io_out_uop_inst : _slots_24_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_90 ? _slots_27_io_out_uop_debug_inst : _GEN_89 ? _slots_26_io_out_uop_debug_inst : _GEN_88 ? _slots_25_io_out_uop_debug_inst : _slots_24_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_90 ? _slots_27_io_out_uop_is_rvc : _GEN_89 ? _slots_26_io_out_uop_is_rvc : _GEN_88 ? _slots_25_io_out_uop_is_rvc : _slots_24_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_90 ? _slots_27_io_out_uop_debug_pc : _GEN_89 ? _slots_26_io_out_uop_debug_pc : _GEN_88 ? _slots_25_io_out_uop_debug_pc : _slots_24_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_90 ? _slots_27_io_out_uop_iq_type : _GEN_89 ? _slots_26_io_out_uop_iq_type : _GEN_88 ? _slots_25_io_out_uop_iq_type : _slots_24_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_90 ? _slots_27_io_out_uop_fu_code : _GEN_89 ? _slots_26_io_out_uop_fu_code : _GEN_88 ? _slots_25_io_out_uop_fu_code : _slots_24_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_90 ? _slots_27_io_out_uop_iw_state : _GEN_89 ? _slots_26_io_out_uop_iw_state : _GEN_88 ? _slots_25_io_out_uop_iw_state : _slots_24_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_90 ? _slots_27_io_out_uop_iw_p1_poisoned : _GEN_89 ? _slots_26_io_out_uop_iw_p1_poisoned : _GEN_88 ? _slots_25_io_out_uop_iw_p1_poisoned : _slots_24_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_90 ? _slots_27_io_out_uop_iw_p2_poisoned : _GEN_89 ? _slots_26_io_out_uop_iw_p2_poisoned : _GEN_88 ? _slots_25_io_out_uop_iw_p2_poisoned : _slots_24_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_90 ? _slots_27_io_out_uop_is_br : _GEN_89 ? _slots_26_io_out_uop_is_br : _GEN_88 ? _slots_25_io_out_uop_is_br : _slots_24_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_90 ? _slots_27_io_out_uop_is_jalr : _GEN_89 ? _slots_26_io_out_uop_is_jalr : _GEN_88 ? _slots_25_io_out_uop_is_jalr : _slots_24_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_90 ? _slots_27_io_out_uop_is_jal : _GEN_89 ? _slots_26_io_out_uop_is_jal : _GEN_88 ? _slots_25_io_out_uop_is_jal : _slots_24_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_90 ? _slots_27_io_out_uop_is_sfb : _GEN_89 ? _slots_26_io_out_uop_is_sfb : _GEN_88 ? _slots_25_io_out_uop_is_sfb : _slots_24_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_90 ? _slots_27_io_out_uop_br_mask : _GEN_89 ? _slots_26_io_out_uop_br_mask : _GEN_88 ? _slots_25_io_out_uop_br_mask : _slots_24_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_90 ? _slots_27_io_out_uop_br_tag : _GEN_89 ? _slots_26_io_out_uop_br_tag : _GEN_88 ? _slots_25_io_out_uop_br_tag : _slots_24_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_90 ? _slots_27_io_out_uop_ftq_idx : _GEN_89 ? _slots_26_io_out_uop_ftq_idx : _GEN_88 ? _slots_25_io_out_uop_ftq_idx : _slots_24_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_90 ? _slots_27_io_out_uop_edge_inst : _GEN_89 ? _slots_26_io_out_uop_edge_inst : _GEN_88 ? _slots_25_io_out_uop_edge_inst : _slots_24_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_90 ? _slots_27_io_out_uop_pc_lob : _GEN_89 ? _slots_26_io_out_uop_pc_lob : _GEN_88 ? _slots_25_io_out_uop_pc_lob : _slots_24_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_90 ? _slots_27_io_out_uop_taken : _GEN_89 ? _slots_26_io_out_uop_taken : _GEN_88 ? _slots_25_io_out_uop_taken : _slots_24_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_90 ? _slots_27_io_out_uop_imm_packed : _GEN_89 ? _slots_26_io_out_uop_imm_packed : _GEN_88 ? _slots_25_io_out_uop_imm_packed : _slots_24_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_90 ? _slots_27_io_out_uop_csr_addr : _GEN_89 ? _slots_26_io_out_uop_csr_addr : _GEN_88 ? _slots_25_io_out_uop_csr_addr : _slots_24_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_90 ? _slots_27_io_out_uop_rob_idx : _GEN_89 ? _slots_26_io_out_uop_rob_idx : _GEN_88 ? _slots_25_io_out_uop_rob_idx : _slots_24_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_90 ? _slots_27_io_out_uop_ldq_idx : _GEN_89 ? _slots_26_io_out_uop_ldq_idx : _GEN_88 ? _slots_25_io_out_uop_ldq_idx : _slots_24_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_90 ? _slots_27_io_out_uop_stq_idx : _GEN_89 ? _slots_26_io_out_uop_stq_idx : _GEN_88 ? _slots_25_io_out_uop_stq_idx : _slots_24_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_90 ? _slots_27_io_out_uop_rxq_idx : _GEN_89 ? _slots_26_io_out_uop_rxq_idx : _GEN_88 ? _slots_25_io_out_uop_rxq_idx : _slots_24_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_90 ? _slots_27_io_out_uop_pdst : _GEN_89 ? _slots_26_io_out_uop_pdst : _GEN_88 ? _slots_25_io_out_uop_pdst : _slots_24_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_90 ? _slots_27_io_out_uop_prs1 : _GEN_89 ? _slots_26_io_out_uop_prs1 : _GEN_88 ? _slots_25_io_out_uop_prs1 : _slots_24_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_90 ? _slots_27_io_out_uop_prs2 : _GEN_89 ? _slots_26_io_out_uop_prs2 : _GEN_88 ? _slots_25_io_out_uop_prs2 : _slots_24_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_90 ? _slots_27_io_out_uop_prs3 : _GEN_89 ? _slots_26_io_out_uop_prs3 : _GEN_88 ? _slots_25_io_out_uop_prs3 : _slots_24_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_90 ? _slots_27_io_out_uop_ppred : _GEN_89 ? _slots_26_io_out_uop_ppred : _GEN_88 ? _slots_25_io_out_uop_ppred : _slots_24_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_90 ? _slots_27_io_out_uop_prs1_busy : _GEN_89 ? _slots_26_io_out_uop_prs1_busy : _GEN_88 ? _slots_25_io_out_uop_prs1_busy : _slots_24_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_90 ? _slots_27_io_out_uop_prs2_busy : _GEN_89 ? _slots_26_io_out_uop_prs2_busy : _GEN_88 ? _slots_25_io_out_uop_prs2_busy : _slots_24_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_90 ? _slots_27_io_out_uop_prs3_busy : _GEN_89 ? _slots_26_io_out_uop_prs3_busy : _GEN_88 ? _slots_25_io_out_uop_prs3_busy : _slots_24_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_90 ? _slots_27_io_out_uop_ppred_busy : _GEN_89 ? _slots_26_io_out_uop_ppred_busy : _GEN_88 ? _slots_25_io_out_uop_ppred_busy : _slots_24_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_90 ? _slots_27_io_out_uop_stale_pdst : _GEN_89 ? _slots_26_io_out_uop_stale_pdst : _GEN_88 ? _slots_25_io_out_uop_stale_pdst : _slots_24_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_90 ? _slots_27_io_out_uop_exception : _GEN_89 ? _slots_26_io_out_uop_exception : _GEN_88 ? _slots_25_io_out_uop_exception : _slots_24_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_90 ? _slots_27_io_out_uop_exc_cause : _GEN_89 ? _slots_26_io_out_uop_exc_cause : _GEN_88 ? _slots_25_io_out_uop_exc_cause : _slots_24_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_90 ? _slots_27_io_out_uop_bypassable : _GEN_89 ? _slots_26_io_out_uop_bypassable : _GEN_88 ? _slots_25_io_out_uop_bypassable : _slots_24_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_90 ? _slots_27_io_out_uop_mem_cmd : _GEN_89 ? _slots_26_io_out_uop_mem_cmd : _GEN_88 ? _slots_25_io_out_uop_mem_cmd : _slots_24_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_90 ? _slots_27_io_out_uop_mem_size : _GEN_89 ? _slots_26_io_out_uop_mem_size : _GEN_88 ? _slots_25_io_out_uop_mem_size : _slots_24_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_90 ? _slots_27_io_out_uop_mem_signed : _GEN_89 ? _slots_26_io_out_uop_mem_signed : _GEN_88 ? _slots_25_io_out_uop_mem_signed : _slots_24_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_90 ? _slots_27_io_out_uop_is_fence : _GEN_89 ? _slots_26_io_out_uop_is_fence : _GEN_88 ? _slots_25_io_out_uop_is_fence : _slots_24_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_90 ? _slots_27_io_out_uop_is_fencei : _GEN_89 ? _slots_26_io_out_uop_is_fencei : _GEN_88 ? _slots_25_io_out_uop_is_fencei : _slots_24_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_90 ? _slots_27_io_out_uop_is_amo : _GEN_89 ? _slots_26_io_out_uop_is_amo : _GEN_88 ? _slots_25_io_out_uop_is_amo : _slots_24_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_90 ? _slots_27_io_out_uop_uses_ldq : _GEN_89 ? _slots_26_io_out_uop_uses_ldq : _GEN_88 ? _slots_25_io_out_uop_uses_ldq : _slots_24_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_90 ? _slots_27_io_out_uop_uses_stq : _GEN_89 ? _slots_26_io_out_uop_uses_stq : _GEN_88 ? _slots_25_io_out_uop_uses_stq : _slots_24_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_90 ? _slots_27_io_out_uop_is_sys_pc2epc : _GEN_89 ? _slots_26_io_out_uop_is_sys_pc2epc : _GEN_88 ? _slots_25_io_out_uop_is_sys_pc2epc : _slots_24_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_90 ? _slots_27_io_out_uop_is_unique : _GEN_89 ? _slots_26_io_out_uop_is_unique : _GEN_88 ? _slots_25_io_out_uop_is_unique : _slots_24_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_90 ? _slots_27_io_out_uop_flush_on_commit : _GEN_89 ? _slots_26_io_out_uop_flush_on_commit : _GEN_88 ? _slots_25_io_out_uop_flush_on_commit : _slots_24_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_90 ? _slots_27_io_out_uop_ldst_is_rs1 : _GEN_89 ? _slots_26_io_out_uop_ldst_is_rs1 : _GEN_88 ? _slots_25_io_out_uop_ldst_is_rs1 : _slots_24_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_90 ? _slots_27_io_out_uop_ldst : _GEN_89 ? _slots_26_io_out_uop_ldst : _GEN_88 ? _slots_25_io_out_uop_ldst : _slots_24_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_90 ? _slots_27_io_out_uop_lrs1 : _GEN_89 ? _slots_26_io_out_uop_lrs1 : _GEN_88 ? _slots_25_io_out_uop_lrs1 : _slots_24_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_90 ? _slots_27_io_out_uop_lrs2 : _GEN_89 ? _slots_26_io_out_uop_lrs2 : _GEN_88 ? _slots_25_io_out_uop_lrs2 : _slots_24_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_90 ? _slots_27_io_out_uop_lrs3 : _GEN_89 ? _slots_26_io_out_uop_lrs3 : _GEN_88 ? _slots_25_io_out_uop_lrs3 : _slots_24_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_90 ? _slots_27_io_out_uop_ldst_val : _GEN_89 ? _slots_26_io_out_uop_ldst_val : _GEN_88 ? _slots_25_io_out_uop_ldst_val : _slots_24_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_90 ? _slots_27_io_out_uop_dst_rtype : _GEN_89 ? _slots_26_io_out_uop_dst_rtype : _GEN_88 ? _slots_25_io_out_uop_dst_rtype : _slots_24_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_90 ? _slots_27_io_out_uop_lrs1_rtype : _GEN_89 ? _slots_26_io_out_uop_lrs1_rtype : _GEN_88 ? _slots_25_io_out_uop_lrs1_rtype : _slots_24_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_90 ? _slots_27_io_out_uop_lrs2_rtype : _GEN_89 ? _slots_26_io_out_uop_lrs2_rtype : _GEN_88 ? _slots_25_io_out_uop_lrs2_rtype : _slots_24_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_90 ? _slots_27_io_out_uop_frs3_en : _GEN_89 ? _slots_26_io_out_uop_frs3_en : _GEN_88 ? _slots_25_io_out_uop_frs3_en : _slots_24_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_90 ? _slots_27_io_out_uop_fp_val : _GEN_89 ? _slots_26_io_out_uop_fp_val : _GEN_88 ? _slots_25_io_out_uop_fp_val : _slots_24_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_90 ? _slots_27_io_out_uop_fp_single : _GEN_89 ? _slots_26_io_out_uop_fp_single : _GEN_88 ? _slots_25_io_out_uop_fp_single : _slots_24_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_90 ? _slots_27_io_out_uop_xcpt_pf_if : _GEN_89 ? _slots_26_io_out_uop_xcpt_pf_if : _GEN_88 ? _slots_25_io_out_uop_xcpt_pf_if : _slots_24_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_90 ? _slots_27_io_out_uop_xcpt_ae_if : _GEN_89 ? _slots_26_io_out_uop_xcpt_ae_if : _GEN_88 ? _slots_25_io_out_uop_xcpt_ae_if : _slots_24_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_90 ? _slots_27_io_out_uop_xcpt_ma_if : _GEN_89 ? _slots_26_io_out_uop_xcpt_ma_if : _GEN_88 ? _slots_25_io_out_uop_xcpt_ma_if : _slots_24_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_90 ? _slots_27_io_out_uop_bp_debug_if : _GEN_89 ? _slots_26_io_out_uop_bp_debug_if : _GEN_88 ? _slots_25_io_out_uop_bp_debug_if : _slots_24_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_90 ? _slots_27_io_out_uop_bp_xcpt_if : _GEN_89 ? _slots_26_io_out_uop_bp_xcpt_if : _GEN_88 ? _slots_25_io_out_uop_bp_xcpt_if : _slots_24_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_90 ? _slots_27_io_out_uop_debug_fsrc : _GEN_89 ? _slots_26_io_out_uop_debug_fsrc : _GEN_88 ? _slots_25_io_out_uop_debug_fsrc : _slots_24_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_90 ? _slots_27_io_out_uop_debug_tsrc : _GEN_89 ? _slots_26_io_out_uop_debug_tsrc : _GEN_88 ? _slots_25_io_out_uop_debug_tsrc : _slots_24_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_23_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_23_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_23_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_23_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_23_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_23_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_23_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_23_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_23_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_23_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_23_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_23_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_23_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_23_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_23_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_23_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_23_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_23_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_23_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_23_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_23_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_23_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_23_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_23_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_23_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_23_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_23_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_23_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_23_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_23_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_23_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_23_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_23_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_23_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_23_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_23_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_23_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_23_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_23_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_23_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_23_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_23_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_23_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_23_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_23_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_23_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_23_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_23_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_23_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_23_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_23_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_23_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_23_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_23_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_23_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_23_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_23_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_23_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_23_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_23_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_23_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_23_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_23_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_23_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_23_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_23_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_23_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_23_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_23_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_23_io_uop_uopc),
    .io_uop_inst                    (_slots_23_io_uop_inst),
    .io_uop_debug_inst              (_slots_23_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_23_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_23_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_23_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_23_io_uop_fu_code),
    .io_uop_iw_state                (_slots_23_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_23_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_23_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_23_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_23_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_23_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_23_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_23_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_23_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_23_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_23_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_23_io_uop_pc_lob),
    .io_uop_taken                   (_slots_23_io_uop_taken),
    .io_uop_imm_packed              (_slots_23_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_23_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_23_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_23_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_23_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_23_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_23_io_uop_pdst),
    .io_uop_prs1                    (_slots_23_io_uop_prs1),
    .io_uop_prs2                    (_slots_23_io_uop_prs2),
    .io_uop_prs3                    (_slots_23_io_uop_prs3),
    .io_uop_ppred                   (_slots_23_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_23_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_23_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_23_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_23_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_23_io_uop_stale_pdst),
    .io_uop_exception               (_slots_23_io_uop_exception),
    .io_uop_exc_cause               (_slots_23_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_23_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_23_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_23_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_23_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_23_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_23_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_23_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_23_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_23_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_23_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_23_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_23_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_23_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_23_io_uop_ldst),
    .io_uop_lrs1                    (_slots_23_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_23_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_23_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_23_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_23_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_23_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_23_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_23_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_23_io_uop_fp_val),
    .io_uop_fp_single               (_slots_23_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_23_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_23_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_23_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_23_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_23_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_23_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_23_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_24 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_24_io_valid),
    .io_will_be_valid               (_slots_24_io_will_be_valid),
    .io_request                     (_slots_24_io_request),
    .io_grant                       (issue_slots_24_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_23),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_24_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_93 ? _slots_28_io_out_uop_uopc : _GEN_92 ? _slots_27_io_out_uop_uopc : _GEN_91 ? _slots_26_io_out_uop_uopc : _slots_25_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_93 ? _slots_28_io_out_uop_inst : _GEN_92 ? _slots_27_io_out_uop_inst : _GEN_91 ? _slots_26_io_out_uop_inst : _slots_25_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_93 ? _slots_28_io_out_uop_debug_inst : _GEN_92 ? _slots_27_io_out_uop_debug_inst : _GEN_91 ? _slots_26_io_out_uop_debug_inst : _slots_25_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_93 ? _slots_28_io_out_uop_is_rvc : _GEN_92 ? _slots_27_io_out_uop_is_rvc : _GEN_91 ? _slots_26_io_out_uop_is_rvc : _slots_25_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_93 ? _slots_28_io_out_uop_debug_pc : _GEN_92 ? _slots_27_io_out_uop_debug_pc : _GEN_91 ? _slots_26_io_out_uop_debug_pc : _slots_25_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_93 ? _slots_28_io_out_uop_iq_type : _GEN_92 ? _slots_27_io_out_uop_iq_type : _GEN_91 ? _slots_26_io_out_uop_iq_type : _slots_25_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_93 ? _slots_28_io_out_uop_fu_code : _GEN_92 ? _slots_27_io_out_uop_fu_code : _GEN_91 ? _slots_26_io_out_uop_fu_code : _slots_25_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_93 ? _slots_28_io_out_uop_iw_state : _GEN_92 ? _slots_27_io_out_uop_iw_state : _GEN_91 ? _slots_26_io_out_uop_iw_state : _slots_25_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_93 ? _slots_28_io_out_uop_iw_p1_poisoned : _GEN_92 ? _slots_27_io_out_uop_iw_p1_poisoned : _GEN_91 ? _slots_26_io_out_uop_iw_p1_poisoned : _slots_25_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_93 ? _slots_28_io_out_uop_iw_p2_poisoned : _GEN_92 ? _slots_27_io_out_uop_iw_p2_poisoned : _GEN_91 ? _slots_26_io_out_uop_iw_p2_poisoned : _slots_25_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_93 ? _slots_28_io_out_uop_is_br : _GEN_92 ? _slots_27_io_out_uop_is_br : _GEN_91 ? _slots_26_io_out_uop_is_br : _slots_25_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_93 ? _slots_28_io_out_uop_is_jalr : _GEN_92 ? _slots_27_io_out_uop_is_jalr : _GEN_91 ? _slots_26_io_out_uop_is_jalr : _slots_25_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_93 ? _slots_28_io_out_uop_is_jal : _GEN_92 ? _slots_27_io_out_uop_is_jal : _GEN_91 ? _slots_26_io_out_uop_is_jal : _slots_25_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_93 ? _slots_28_io_out_uop_is_sfb : _GEN_92 ? _slots_27_io_out_uop_is_sfb : _GEN_91 ? _slots_26_io_out_uop_is_sfb : _slots_25_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_93 ? _slots_28_io_out_uop_br_mask : _GEN_92 ? _slots_27_io_out_uop_br_mask : _GEN_91 ? _slots_26_io_out_uop_br_mask : _slots_25_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_93 ? _slots_28_io_out_uop_br_tag : _GEN_92 ? _slots_27_io_out_uop_br_tag : _GEN_91 ? _slots_26_io_out_uop_br_tag : _slots_25_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_93 ? _slots_28_io_out_uop_ftq_idx : _GEN_92 ? _slots_27_io_out_uop_ftq_idx : _GEN_91 ? _slots_26_io_out_uop_ftq_idx : _slots_25_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_93 ? _slots_28_io_out_uop_edge_inst : _GEN_92 ? _slots_27_io_out_uop_edge_inst : _GEN_91 ? _slots_26_io_out_uop_edge_inst : _slots_25_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_93 ? _slots_28_io_out_uop_pc_lob : _GEN_92 ? _slots_27_io_out_uop_pc_lob : _GEN_91 ? _slots_26_io_out_uop_pc_lob : _slots_25_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_93 ? _slots_28_io_out_uop_taken : _GEN_92 ? _slots_27_io_out_uop_taken : _GEN_91 ? _slots_26_io_out_uop_taken : _slots_25_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_93 ? _slots_28_io_out_uop_imm_packed : _GEN_92 ? _slots_27_io_out_uop_imm_packed : _GEN_91 ? _slots_26_io_out_uop_imm_packed : _slots_25_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_93 ? _slots_28_io_out_uop_csr_addr : _GEN_92 ? _slots_27_io_out_uop_csr_addr : _GEN_91 ? _slots_26_io_out_uop_csr_addr : _slots_25_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_93 ? _slots_28_io_out_uop_rob_idx : _GEN_92 ? _slots_27_io_out_uop_rob_idx : _GEN_91 ? _slots_26_io_out_uop_rob_idx : _slots_25_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_93 ? _slots_28_io_out_uop_ldq_idx : _GEN_92 ? _slots_27_io_out_uop_ldq_idx : _GEN_91 ? _slots_26_io_out_uop_ldq_idx : _slots_25_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_93 ? _slots_28_io_out_uop_stq_idx : _GEN_92 ? _slots_27_io_out_uop_stq_idx : _GEN_91 ? _slots_26_io_out_uop_stq_idx : _slots_25_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_93 ? _slots_28_io_out_uop_rxq_idx : _GEN_92 ? _slots_27_io_out_uop_rxq_idx : _GEN_91 ? _slots_26_io_out_uop_rxq_idx : _slots_25_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_93 ? _slots_28_io_out_uop_pdst : _GEN_92 ? _slots_27_io_out_uop_pdst : _GEN_91 ? _slots_26_io_out_uop_pdst : _slots_25_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_93 ? _slots_28_io_out_uop_prs1 : _GEN_92 ? _slots_27_io_out_uop_prs1 : _GEN_91 ? _slots_26_io_out_uop_prs1 : _slots_25_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_93 ? _slots_28_io_out_uop_prs2 : _GEN_92 ? _slots_27_io_out_uop_prs2 : _GEN_91 ? _slots_26_io_out_uop_prs2 : _slots_25_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_93 ? _slots_28_io_out_uop_prs3 : _GEN_92 ? _slots_27_io_out_uop_prs3 : _GEN_91 ? _slots_26_io_out_uop_prs3 : _slots_25_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_93 ? _slots_28_io_out_uop_ppred : _GEN_92 ? _slots_27_io_out_uop_ppred : _GEN_91 ? _slots_26_io_out_uop_ppred : _slots_25_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_93 ? _slots_28_io_out_uop_prs1_busy : _GEN_92 ? _slots_27_io_out_uop_prs1_busy : _GEN_91 ? _slots_26_io_out_uop_prs1_busy : _slots_25_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_93 ? _slots_28_io_out_uop_prs2_busy : _GEN_92 ? _slots_27_io_out_uop_prs2_busy : _GEN_91 ? _slots_26_io_out_uop_prs2_busy : _slots_25_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_93 ? _slots_28_io_out_uop_prs3_busy : _GEN_92 ? _slots_27_io_out_uop_prs3_busy : _GEN_91 ? _slots_26_io_out_uop_prs3_busy : _slots_25_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_93 ? _slots_28_io_out_uop_ppred_busy : _GEN_92 ? _slots_27_io_out_uop_ppred_busy : _GEN_91 ? _slots_26_io_out_uop_ppred_busy : _slots_25_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_93 ? _slots_28_io_out_uop_stale_pdst : _GEN_92 ? _slots_27_io_out_uop_stale_pdst : _GEN_91 ? _slots_26_io_out_uop_stale_pdst : _slots_25_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_93 ? _slots_28_io_out_uop_exception : _GEN_92 ? _slots_27_io_out_uop_exception : _GEN_91 ? _slots_26_io_out_uop_exception : _slots_25_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_93 ? _slots_28_io_out_uop_exc_cause : _GEN_92 ? _slots_27_io_out_uop_exc_cause : _GEN_91 ? _slots_26_io_out_uop_exc_cause : _slots_25_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_93 ? _slots_28_io_out_uop_bypassable : _GEN_92 ? _slots_27_io_out_uop_bypassable : _GEN_91 ? _slots_26_io_out_uop_bypassable : _slots_25_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_93 ? _slots_28_io_out_uop_mem_cmd : _GEN_92 ? _slots_27_io_out_uop_mem_cmd : _GEN_91 ? _slots_26_io_out_uop_mem_cmd : _slots_25_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_93 ? _slots_28_io_out_uop_mem_size : _GEN_92 ? _slots_27_io_out_uop_mem_size : _GEN_91 ? _slots_26_io_out_uop_mem_size : _slots_25_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_93 ? _slots_28_io_out_uop_mem_signed : _GEN_92 ? _slots_27_io_out_uop_mem_signed : _GEN_91 ? _slots_26_io_out_uop_mem_signed : _slots_25_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_93 ? _slots_28_io_out_uop_is_fence : _GEN_92 ? _slots_27_io_out_uop_is_fence : _GEN_91 ? _slots_26_io_out_uop_is_fence : _slots_25_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_93 ? _slots_28_io_out_uop_is_fencei : _GEN_92 ? _slots_27_io_out_uop_is_fencei : _GEN_91 ? _slots_26_io_out_uop_is_fencei : _slots_25_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_93 ? _slots_28_io_out_uop_is_amo : _GEN_92 ? _slots_27_io_out_uop_is_amo : _GEN_91 ? _slots_26_io_out_uop_is_amo : _slots_25_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_93 ? _slots_28_io_out_uop_uses_ldq : _GEN_92 ? _slots_27_io_out_uop_uses_ldq : _GEN_91 ? _slots_26_io_out_uop_uses_ldq : _slots_25_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_93 ? _slots_28_io_out_uop_uses_stq : _GEN_92 ? _slots_27_io_out_uop_uses_stq : _GEN_91 ? _slots_26_io_out_uop_uses_stq : _slots_25_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_93 ? _slots_28_io_out_uop_is_sys_pc2epc : _GEN_92 ? _slots_27_io_out_uop_is_sys_pc2epc : _GEN_91 ? _slots_26_io_out_uop_is_sys_pc2epc : _slots_25_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_93 ? _slots_28_io_out_uop_is_unique : _GEN_92 ? _slots_27_io_out_uop_is_unique : _GEN_91 ? _slots_26_io_out_uop_is_unique : _slots_25_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_93 ? _slots_28_io_out_uop_flush_on_commit : _GEN_92 ? _slots_27_io_out_uop_flush_on_commit : _GEN_91 ? _slots_26_io_out_uop_flush_on_commit : _slots_25_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_93 ? _slots_28_io_out_uop_ldst_is_rs1 : _GEN_92 ? _slots_27_io_out_uop_ldst_is_rs1 : _GEN_91 ? _slots_26_io_out_uop_ldst_is_rs1 : _slots_25_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_93 ? _slots_28_io_out_uop_ldst : _GEN_92 ? _slots_27_io_out_uop_ldst : _GEN_91 ? _slots_26_io_out_uop_ldst : _slots_25_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_93 ? _slots_28_io_out_uop_lrs1 : _GEN_92 ? _slots_27_io_out_uop_lrs1 : _GEN_91 ? _slots_26_io_out_uop_lrs1 : _slots_25_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_93 ? _slots_28_io_out_uop_lrs2 : _GEN_92 ? _slots_27_io_out_uop_lrs2 : _GEN_91 ? _slots_26_io_out_uop_lrs2 : _slots_25_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_93 ? _slots_28_io_out_uop_lrs3 : _GEN_92 ? _slots_27_io_out_uop_lrs3 : _GEN_91 ? _slots_26_io_out_uop_lrs3 : _slots_25_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_93 ? _slots_28_io_out_uop_ldst_val : _GEN_92 ? _slots_27_io_out_uop_ldst_val : _GEN_91 ? _slots_26_io_out_uop_ldst_val : _slots_25_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_93 ? _slots_28_io_out_uop_dst_rtype : _GEN_92 ? _slots_27_io_out_uop_dst_rtype : _GEN_91 ? _slots_26_io_out_uop_dst_rtype : _slots_25_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_93 ? _slots_28_io_out_uop_lrs1_rtype : _GEN_92 ? _slots_27_io_out_uop_lrs1_rtype : _GEN_91 ? _slots_26_io_out_uop_lrs1_rtype : _slots_25_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_93 ? _slots_28_io_out_uop_lrs2_rtype : _GEN_92 ? _slots_27_io_out_uop_lrs2_rtype : _GEN_91 ? _slots_26_io_out_uop_lrs2_rtype : _slots_25_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_93 ? _slots_28_io_out_uop_frs3_en : _GEN_92 ? _slots_27_io_out_uop_frs3_en : _GEN_91 ? _slots_26_io_out_uop_frs3_en : _slots_25_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_93 ? _slots_28_io_out_uop_fp_val : _GEN_92 ? _slots_27_io_out_uop_fp_val : _GEN_91 ? _slots_26_io_out_uop_fp_val : _slots_25_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_93 ? _slots_28_io_out_uop_fp_single : _GEN_92 ? _slots_27_io_out_uop_fp_single : _GEN_91 ? _slots_26_io_out_uop_fp_single : _slots_25_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_93 ? _slots_28_io_out_uop_xcpt_pf_if : _GEN_92 ? _slots_27_io_out_uop_xcpt_pf_if : _GEN_91 ? _slots_26_io_out_uop_xcpt_pf_if : _slots_25_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_93 ? _slots_28_io_out_uop_xcpt_ae_if : _GEN_92 ? _slots_27_io_out_uop_xcpt_ae_if : _GEN_91 ? _slots_26_io_out_uop_xcpt_ae_if : _slots_25_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_93 ? _slots_28_io_out_uop_xcpt_ma_if : _GEN_92 ? _slots_27_io_out_uop_xcpt_ma_if : _GEN_91 ? _slots_26_io_out_uop_xcpt_ma_if : _slots_25_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_93 ? _slots_28_io_out_uop_bp_debug_if : _GEN_92 ? _slots_27_io_out_uop_bp_debug_if : _GEN_91 ? _slots_26_io_out_uop_bp_debug_if : _slots_25_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_93 ? _slots_28_io_out_uop_bp_xcpt_if : _GEN_92 ? _slots_27_io_out_uop_bp_xcpt_if : _GEN_91 ? _slots_26_io_out_uop_bp_xcpt_if : _slots_25_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_93 ? _slots_28_io_out_uop_debug_fsrc : _GEN_92 ? _slots_27_io_out_uop_debug_fsrc : _GEN_91 ? _slots_26_io_out_uop_debug_fsrc : _slots_25_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_93 ? _slots_28_io_out_uop_debug_tsrc : _GEN_92 ? _slots_27_io_out_uop_debug_tsrc : _GEN_91 ? _slots_26_io_out_uop_debug_tsrc : _slots_25_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_24_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_24_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_24_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_24_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_24_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_24_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_24_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_24_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_24_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_24_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_24_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_24_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_24_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_24_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_24_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_24_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_24_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_24_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_24_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_24_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_24_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_24_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_24_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_24_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_24_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_24_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_24_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_24_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_24_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_24_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_24_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_24_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_24_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_24_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_24_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_24_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_24_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_24_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_24_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_24_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_24_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_24_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_24_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_24_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_24_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_24_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_24_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_24_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_24_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_24_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_24_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_24_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_24_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_24_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_24_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_24_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_24_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_24_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_24_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_24_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_24_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_24_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_24_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_24_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_24_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_24_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_24_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_24_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_24_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_24_io_uop_uopc),
    .io_uop_inst                    (_slots_24_io_uop_inst),
    .io_uop_debug_inst              (_slots_24_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_24_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_24_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_24_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_24_io_uop_fu_code),
    .io_uop_iw_state                (_slots_24_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_24_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_24_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_24_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_24_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_24_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_24_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_24_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_24_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_24_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_24_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_24_io_uop_pc_lob),
    .io_uop_taken                   (_slots_24_io_uop_taken),
    .io_uop_imm_packed              (_slots_24_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_24_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_24_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_24_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_24_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_24_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_24_io_uop_pdst),
    .io_uop_prs1                    (_slots_24_io_uop_prs1),
    .io_uop_prs2                    (_slots_24_io_uop_prs2),
    .io_uop_prs3                    (_slots_24_io_uop_prs3),
    .io_uop_ppred                   (_slots_24_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_24_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_24_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_24_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_24_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_24_io_uop_stale_pdst),
    .io_uop_exception               (_slots_24_io_uop_exception),
    .io_uop_exc_cause               (_slots_24_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_24_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_24_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_24_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_24_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_24_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_24_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_24_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_24_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_24_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_24_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_24_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_24_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_24_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_24_io_uop_ldst),
    .io_uop_lrs1                    (_slots_24_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_24_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_24_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_24_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_24_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_24_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_24_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_24_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_24_io_uop_fp_val),
    .io_uop_fp_single               (_slots_24_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_24_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_24_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_24_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_24_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_24_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_24_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_24_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_25 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_25_io_valid),
    .io_will_be_valid               (_slots_25_io_will_be_valid),
    .io_request                     (_slots_25_io_request),
    .io_grant                       (issue_slots_25_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_24),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_25_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_96 ? _slots_29_io_out_uop_uopc : _GEN_95 ? _slots_28_io_out_uop_uopc : _GEN_94 ? _slots_27_io_out_uop_uopc : _slots_26_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_96 ? _slots_29_io_out_uop_inst : _GEN_95 ? _slots_28_io_out_uop_inst : _GEN_94 ? _slots_27_io_out_uop_inst : _slots_26_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_96 ? _slots_29_io_out_uop_debug_inst : _GEN_95 ? _slots_28_io_out_uop_debug_inst : _GEN_94 ? _slots_27_io_out_uop_debug_inst : _slots_26_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_96 ? _slots_29_io_out_uop_is_rvc : _GEN_95 ? _slots_28_io_out_uop_is_rvc : _GEN_94 ? _slots_27_io_out_uop_is_rvc : _slots_26_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_96 ? _slots_29_io_out_uop_debug_pc : _GEN_95 ? _slots_28_io_out_uop_debug_pc : _GEN_94 ? _slots_27_io_out_uop_debug_pc : _slots_26_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_96 ? _slots_29_io_out_uop_iq_type : _GEN_95 ? _slots_28_io_out_uop_iq_type : _GEN_94 ? _slots_27_io_out_uop_iq_type : _slots_26_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_96 ? _slots_29_io_out_uop_fu_code : _GEN_95 ? _slots_28_io_out_uop_fu_code : _GEN_94 ? _slots_27_io_out_uop_fu_code : _slots_26_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_96 ? _slots_29_io_out_uop_iw_state : _GEN_95 ? _slots_28_io_out_uop_iw_state : _GEN_94 ? _slots_27_io_out_uop_iw_state : _slots_26_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_96 ? _slots_29_io_out_uop_iw_p1_poisoned : _GEN_95 ? _slots_28_io_out_uop_iw_p1_poisoned : _GEN_94 ? _slots_27_io_out_uop_iw_p1_poisoned : _slots_26_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_96 ? _slots_29_io_out_uop_iw_p2_poisoned : _GEN_95 ? _slots_28_io_out_uop_iw_p2_poisoned : _GEN_94 ? _slots_27_io_out_uop_iw_p2_poisoned : _slots_26_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_96 ? _slots_29_io_out_uop_is_br : _GEN_95 ? _slots_28_io_out_uop_is_br : _GEN_94 ? _slots_27_io_out_uop_is_br : _slots_26_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_96 ? _slots_29_io_out_uop_is_jalr : _GEN_95 ? _slots_28_io_out_uop_is_jalr : _GEN_94 ? _slots_27_io_out_uop_is_jalr : _slots_26_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_96 ? _slots_29_io_out_uop_is_jal : _GEN_95 ? _slots_28_io_out_uop_is_jal : _GEN_94 ? _slots_27_io_out_uop_is_jal : _slots_26_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_96 ? _slots_29_io_out_uop_is_sfb : _GEN_95 ? _slots_28_io_out_uop_is_sfb : _GEN_94 ? _slots_27_io_out_uop_is_sfb : _slots_26_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_96 ? _slots_29_io_out_uop_br_mask : _GEN_95 ? _slots_28_io_out_uop_br_mask : _GEN_94 ? _slots_27_io_out_uop_br_mask : _slots_26_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_96 ? _slots_29_io_out_uop_br_tag : _GEN_95 ? _slots_28_io_out_uop_br_tag : _GEN_94 ? _slots_27_io_out_uop_br_tag : _slots_26_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_96 ? _slots_29_io_out_uop_ftq_idx : _GEN_95 ? _slots_28_io_out_uop_ftq_idx : _GEN_94 ? _slots_27_io_out_uop_ftq_idx : _slots_26_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_96 ? _slots_29_io_out_uop_edge_inst : _GEN_95 ? _slots_28_io_out_uop_edge_inst : _GEN_94 ? _slots_27_io_out_uop_edge_inst : _slots_26_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_96 ? _slots_29_io_out_uop_pc_lob : _GEN_95 ? _slots_28_io_out_uop_pc_lob : _GEN_94 ? _slots_27_io_out_uop_pc_lob : _slots_26_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_96 ? _slots_29_io_out_uop_taken : _GEN_95 ? _slots_28_io_out_uop_taken : _GEN_94 ? _slots_27_io_out_uop_taken : _slots_26_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_96 ? _slots_29_io_out_uop_imm_packed : _GEN_95 ? _slots_28_io_out_uop_imm_packed : _GEN_94 ? _slots_27_io_out_uop_imm_packed : _slots_26_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_96 ? _slots_29_io_out_uop_csr_addr : _GEN_95 ? _slots_28_io_out_uop_csr_addr : _GEN_94 ? _slots_27_io_out_uop_csr_addr : _slots_26_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_96 ? _slots_29_io_out_uop_rob_idx : _GEN_95 ? _slots_28_io_out_uop_rob_idx : _GEN_94 ? _slots_27_io_out_uop_rob_idx : _slots_26_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_96 ? _slots_29_io_out_uop_ldq_idx : _GEN_95 ? _slots_28_io_out_uop_ldq_idx : _GEN_94 ? _slots_27_io_out_uop_ldq_idx : _slots_26_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_96 ? _slots_29_io_out_uop_stq_idx : _GEN_95 ? _slots_28_io_out_uop_stq_idx : _GEN_94 ? _slots_27_io_out_uop_stq_idx : _slots_26_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_96 ? _slots_29_io_out_uop_rxq_idx : _GEN_95 ? _slots_28_io_out_uop_rxq_idx : _GEN_94 ? _slots_27_io_out_uop_rxq_idx : _slots_26_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_96 ? _slots_29_io_out_uop_pdst : _GEN_95 ? _slots_28_io_out_uop_pdst : _GEN_94 ? _slots_27_io_out_uop_pdst : _slots_26_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_96 ? _slots_29_io_out_uop_prs1 : _GEN_95 ? _slots_28_io_out_uop_prs1 : _GEN_94 ? _slots_27_io_out_uop_prs1 : _slots_26_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_96 ? _slots_29_io_out_uop_prs2 : _GEN_95 ? _slots_28_io_out_uop_prs2 : _GEN_94 ? _slots_27_io_out_uop_prs2 : _slots_26_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_96 ? _slots_29_io_out_uop_prs3 : _GEN_95 ? _slots_28_io_out_uop_prs3 : _GEN_94 ? _slots_27_io_out_uop_prs3 : _slots_26_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_96 ? _slots_29_io_out_uop_ppred : _GEN_95 ? _slots_28_io_out_uop_ppred : _GEN_94 ? _slots_27_io_out_uop_ppred : _slots_26_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_96 ? _slots_29_io_out_uop_prs1_busy : _GEN_95 ? _slots_28_io_out_uop_prs1_busy : _GEN_94 ? _slots_27_io_out_uop_prs1_busy : _slots_26_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_96 ? _slots_29_io_out_uop_prs2_busy : _GEN_95 ? _slots_28_io_out_uop_prs2_busy : _GEN_94 ? _slots_27_io_out_uop_prs2_busy : _slots_26_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_96 ? _slots_29_io_out_uop_prs3_busy : _GEN_95 ? _slots_28_io_out_uop_prs3_busy : _GEN_94 ? _slots_27_io_out_uop_prs3_busy : _slots_26_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_96 ? _slots_29_io_out_uop_ppred_busy : _GEN_95 ? _slots_28_io_out_uop_ppred_busy : _GEN_94 ? _slots_27_io_out_uop_ppred_busy : _slots_26_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_96 ? _slots_29_io_out_uop_stale_pdst : _GEN_95 ? _slots_28_io_out_uop_stale_pdst : _GEN_94 ? _slots_27_io_out_uop_stale_pdst : _slots_26_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_96 ? _slots_29_io_out_uop_exception : _GEN_95 ? _slots_28_io_out_uop_exception : _GEN_94 ? _slots_27_io_out_uop_exception : _slots_26_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_96 ? _slots_29_io_out_uop_exc_cause : _GEN_95 ? _slots_28_io_out_uop_exc_cause : _GEN_94 ? _slots_27_io_out_uop_exc_cause : _slots_26_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_96 ? _slots_29_io_out_uop_bypassable : _GEN_95 ? _slots_28_io_out_uop_bypassable : _GEN_94 ? _slots_27_io_out_uop_bypassable : _slots_26_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_96 ? _slots_29_io_out_uop_mem_cmd : _GEN_95 ? _slots_28_io_out_uop_mem_cmd : _GEN_94 ? _slots_27_io_out_uop_mem_cmd : _slots_26_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_96 ? _slots_29_io_out_uop_mem_size : _GEN_95 ? _slots_28_io_out_uop_mem_size : _GEN_94 ? _slots_27_io_out_uop_mem_size : _slots_26_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_96 ? _slots_29_io_out_uop_mem_signed : _GEN_95 ? _slots_28_io_out_uop_mem_signed : _GEN_94 ? _slots_27_io_out_uop_mem_signed : _slots_26_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_96 ? _slots_29_io_out_uop_is_fence : _GEN_95 ? _slots_28_io_out_uop_is_fence : _GEN_94 ? _slots_27_io_out_uop_is_fence : _slots_26_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_96 ? _slots_29_io_out_uop_is_fencei : _GEN_95 ? _slots_28_io_out_uop_is_fencei : _GEN_94 ? _slots_27_io_out_uop_is_fencei : _slots_26_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_96 ? _slots_29_io_out_uop_is_amo : _GEN_95 ? _slots_28_io_out_uop_is_amo : _GEN_94 ? _slots_27_io_out_uop_is_amo : _slots_26_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_96 ? _slots_29_io_out_uop_uses_ldq : _GEN_95 ? _slots_28_io_out_uop_uses_ldq : _GEN_94 ? _slots_27_io_out_uop_uses_ldq : _slots_26_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_96 ? _slots_29_io_out_uop_uses_stq : _GEN_95 ? _slots_28_io_out_uop_uses_stq : _GEN_94 ? _slots_27_io_out_uop_uses_stq : _slots_26_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_96 ? _slots_29_io_out_uop_is_sys_pc2epc : _GEN_95 ? _slots_28_io_out_uop_is_sys_pc2epc : _GEN_94 ? _slots_27_io_out_uop_is_sys_pc2epc : _slots_26_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_96 ? _slots_29_io_out_uop_is_unique : _GEN_95 ? _slots_28_io_out_uop_is_unique : _GEN_94 ? _slots_27_io_out_uop_is_unique : _slots_26_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_96 ? _slots_29_io_out_uop_flush_on_commit : _GEN_95 ? _slots_28_io_out_uop_flush_on_commit : _GEN_94 ? _slots_27_io_out_uop_flush_on_commit : _slots_26_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_96 ? _slots_29_io_out_uop_ldst_is_rs1 : _GEN_95 ? _slots_28_io_out_uop_ldst_is_rs1 : _GEN_94 ? _slots_27_io_out_uop_ldst_is_rs1 : _slots_26_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_96 ? _slots_29_io_out_uop_ldst : _GEN_95 ? _slots_28_io_out_uop_ldst : _GEN_94 ? _slots_27_io_out_uop_ldst : _slots_26_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_96 ? _slots_29_io_out_uop_lrs1 : _GEN_95 ? _slots_28_io_out_uop_lrs1 : _GEN_94 ? _slots_27_io_out_uop_lrs1 : _slots_26_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_96 ? _slots_29_io_out_uop_lrs2 : _GEN_95 ? _slots_28_io_out_uop_lrs2 : _GEN_94 ? _slots_27_io_out_uop_lrs2 : _slots_26_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_96 ? _slots_29_io_out_uop_lrs3 : _GEN_95 ? _slots_28_io_out_uop_lrs3 : _GEN_94 ? _slots_27_io_out_uop_lrs3 : _slots_26_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_96 ? _slots_29_io_out_uop_ldst_val : _GEN_95 ? _slots_28_io_out_uop_ldst_val : _GEN_94 ? _slots_27_io_out_uop_ldst_val : _slots_26_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_96 ? _slots_29_io_out_uop_dst_rtype : _GEN_95 ? _slots_28_io_out_uop_dst_rtype : _GEN_94 ? _slots_27_io_out_uop_dst_rtype : _slots_26_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_96 ? _slots_29_io_out_uop_lrs1_rtype : _GEN_95 ? _slots_28_io_out_uop_lrs1_rtype : _GEN_94 ? _slots_27_io_out_uop_lrs1_rtype : _slots_26_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_96 ? _slots_29_io_out_uop_lrs2_rtype : _GEN_95 ? _slots_28_io_out_uop_lrs2_rtype : _GEN_94 ? _slots_27_io_out_uop_lrs2_rtype : _slots_26_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_96 ? _slots_29_io_out_uop_frs3_en : _GEN_95 ? _slots_28_io_out_uop_frs3_en : _GEN_94 ? _slots_27_io_out_uop_frs3_en : _slots_26_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_96 ? _slots_29_io_out_uop_fp_val : _GEN_95 ? _slots_28_io_out_uop_fp_val : _GEN_94 ? _slots_27_io_out_uop_fp_val : _slots_26_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_96 ? _slots_29_io_out_uop_fp_single : _GEN_95 ? _slots_28_io_out_uop_fp_single : _GEN_94 ? _slots_27_io_out_uop_fp_single : _slots_26_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_96 ? _slots_29_io_out_uop_xcpt_pf_if : _GEN_95 ? _slots_28_io_out_uop_xcpt_pf_if : _GEN_94 ? _slots_27_io_out_uop_xcpt_pf_if : _slots_26_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_96 ? _slots_29_io_out_uop_xcpt_ae_if : _GEN_95 ? _slots_28_io_out_uop_xcpt_ae_if : _GEN_94 ? _slots_27_io_out_uop_xcpt_ae_if : _slots_26_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_96 ? _slots_29_io_out_uop_xcpt_ma_if : _GEN_95 ? _slots_28_io_out_uop_xcpt_ma_if : _GEN_94 ? _slots_27_io_out_uop_xcpt_ma_if : _slots_26_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_96 ? _slots_29_io_out_uop_bp_debug_if : _GEN_95 ? _slots_28_io_out_uop_bp_debug_if : _GEN_94 ? _slots_27_io_out_uop_bp_debug_if : _slots_26_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_96 ? _slots_29_io_out_uop_bp_xcpt_if : _GEN_95 ? _slots_28_io_out_uop_bp_xcpt_if : _GEN_94 ? _slots_27_io_out_uop_bp_xcpt_if : _slots_26_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_96 ? _slots_29_io_out_uop_debug_fsrc : _GEN_95 ? _slots_28_io_out_uop_debug_fsrc : _GEN_94 ? _slots_27_io_out_uop_debug_fsrc : _slots_26_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_96 ? _slots_29_io_out_uop_debug_tsrc : _GEN_95 ? _slots_28_io_out_uop_debug_tsrc : _GEN_94 ? _slots_27_io_out_uop_debug_tsrc : _slots_26_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_25_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_25_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_25_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_25_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_25_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_25_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_25_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_25_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_25_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_25_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_25_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_25_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_25_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_25_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_25_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_25_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_25_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_25_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_25_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_25_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_25_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_25_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_25_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_25_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_25_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_25_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_25_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_25_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_25_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_25_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_25_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_25_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_25_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_25_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_25_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_25_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_25_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_25_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_25_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_25_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_25_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_25_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_25_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_25_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_25_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_25_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_25_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_25_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_25_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_25_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_25_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_25_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_25_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_25_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_25_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_25_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_25_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_25_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_25_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_25_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_25_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_25_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_25_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_25_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_25_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_25_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_25_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_25_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_25_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_25_io_uop_uopc),
    .io_uop_inst                    (_slots_25_io_uop_inst),
    .io_uop_debug_inst              (_slots_25_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_25_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_25_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_25_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_25_io_uop_fu_code),
    .io_uop_iw_state                (_slots_25_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_25_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_25_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_25_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_25_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_25_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_25_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_25_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_25_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_25_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_25_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_25_io_uop_pc_lob),
    .io_uop_taken                   (_slots_25_io_uop_taken),
    .io_uop_imm_packed              (_slots_25_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_25_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_25_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_25_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_25_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_25_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_25_io_uop_pdst),
    .io_uop_prs1                    (_slots_25_io_uop_prs1),
    .io_uop_prs2                    (_slots_25_io_uop_prs2),
    .io_uop_prs3                    (_slots_25_io_uop_prs3),
    .io_uop_ppred                   (_slots_25_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_25_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_25_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_25_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_25_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_25_io_uop_stale_pdst),
    .io_uop_exception               (_slots_25_io_uop_exception),
    .io_uop_exc_cause               (_slots_25_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_25_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_25_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_25_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_25_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_25_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_25_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_25_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_25_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_25_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_25_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_25_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_25_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_25_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_25_io_uop_ldst),
    .io_uop_lrs1                    (_slots_25_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_25_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_25_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_25_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_25_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_25_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_25_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_25_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_25_io_uop_fp_val),
    .io_uop_fp_single               (_slots_25_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_25_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_25_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_25_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_25_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_25_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_25_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_25_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_26 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_26_io_valid),
    .io_will_be_valid               (_slots_26_io_will_be_valid),
    .io_request                     (_slots_26_io_request),
    .io_grant                       (issue_slots_26_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_25),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_26_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_99 ? _slots_30_io_out_uop_uopc : _GEN_98 ? _slots_29_io_out_uop_uopc : _GEN_97 ? _slots_28_io_out_uop_uopc : _slots_27_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_99 ? _slots_30_io_out_uop_inst : _GEN_98 ? _slots_29_io_out_uop_inst : _GEN_97 ? _slots_28_io_out_uop_inst : _slots_27_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_99 ? _slots_30_io_out_uop_debug_inst : _GEN_98 ? _slots_29_io_out_uop_debug_inst : _GEN_97 ? _slots_28_io_out_uop_debug_inst : _slots_27_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_99 ? _slots_30_io_out_uop_is_rvc : _GEN_98 ? _slots_29_io_out_uop_is_rvc : _GEN_97 ? _slots_28_io_out_uop_is_rvc : _slots_27_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_99 ? _slots_30_io_out_uop_debug_pc : _GEN_98 ? _slots_29_io_out_uop_debug_pc : _GEN_97 ? _slots_28_io_out_uop_debug_pc : _slots_27_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_99 ? _slots_30_io_out_uop_iq_type : _GEN_98 ? _slots_29_io_out_uop_iq_type : _GEN_97 ? _slots_28_io_out_uop_iq_type : _slots_27_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_99 ? _slots_30_io_out_uop_fu_code : _GEN_98 ? _slots_29_io_out_uop_fu_code : _GEN_97 ? _slots_28_io_out_uop_fu_code : _slots_27_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_99 ? _slots_30_io_out_uop_iw_state : _GEN_98 ? _slots_29_io_out_uop_iw_state : _GEN_97 ? _slots_28_io_out_uop_iw_state : _slots_27_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_99 ? _slots_30_io_out_uop_iw_p1_poisoned : _GEN_98 ? _slots_29_io_out_uop_iw_p1_poisoned : _GEN_97 ? _slots_28_io_out_uop_iw_p1_poisoned : _slots_27_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_99 ? _slots_30_io_out_uop_iw_p2_poisoned : _GEN_98 ? _slots_29_io_out_uop_iw_p2_poisoned : _GEN_97 ? _slots_28_io_out_uop_iw_p2_poisoned : _slots_27_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_99 ? _slots_30_io_out_uop_is_br : _GEN_98 ? _slots_29_io_out_uop_is_br : _GEN_97 ? _slots_28_io_out_uop_is_br : _slots_27_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_99 ? _slots_30_io_out_uop_is_jalr : _GEN_98 ? _slots_29_io_out_uop_is_jalr : _GEN_97 ? _slots_28_io_out_uop_is_jalr : _slots_27_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_99 ? _slots_30_io_out_uop_is_jal : _GEN_98 ? _slots_29_io_out_uop_is_jal : _GEN_97 ? _slots_28_io_out_uop_is_jal : _slots_27_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_99 ? _slots_30_io_out_uop_is_sfb : _GEN_98 ? _slots_29_io_out_uop_is_sfb : _GEN_97 ? _slots_28_io_out_uop_is_sfb : _slots_27_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_99 ? _slots_30_io_out_uop_br_mask : _GEN_98 ? _slots_29_io_out_uop_br_mask : _GEN_97 ? _slots_28_io_out_uop_br_mask : _slots_27_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_99 ? _slots_30_io_out_uop_br_tag : _GEN_98 ? _slots_29_io_out_uop_br_tag : _GEN_97 ? _slots_28_io_out_uop_br_tag : _slots_27_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_99 ? _slots_30_io_out_uop_ftq_idx : _GEN_98 ? _slots_29_io_out_uop_ftq_idx : _GEN_97 ? _slots_28_io_out_uop_ftq_idx : _slots_27_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_99 ? _slots_30_io_out_uop_edge_inst : _GEN_98 ? _slots_29_io_out_uop_edge_inst : _GEN_97 ? _slots_28_io_out_uop_edge_inst : _slots_27_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_99 ? _slots_30_io_out_uop_pc_lob : _GEN_98 ? _slots_29_io_out_uop_pc_lob : _GEN_97 ? _slots_28_io_out_uop_pc_lob : _slots_27_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_99 ? _slots_30_io_out_uop_taken : _GEN_98 ? _slots_29_io_out_uop_taken : _GEN_97 ? _slots_28_io_out_uop_taken : _slots_27_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_99 ? _slots_30_io_out_uop_imm_packed : _GEN_98 ? _slots_29_io_out_uop_imm_packed : _GEN_97 ? _slots_28_io_out_uop_imm_packed : _slots_27_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_99 ? _slots_30_io_out_uop_csr_addr : _GEN_98 ? _slots_29_io_out_uop_csr_addr : _GEN_97 ? _slots_28_io_out_uop_csr_addr : _slots_27_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_99 ? _slots_30_io_out_uop_rob_idx : _GEN_98 ? _slots_29_io_out_uop_rob_idx : _GEN_97 ? _slots_28_io_out_uop_rob_idx : _slots_27_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_99 ? _slots_30_io_out_uop_ldq_idx : _GEN_98 ? _slots_29_io_out_uop_ldq_idx : _GEN_97 ? _slots_28_io_out_uop_ldq_idx : _slots_27_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_99 ? _slots_30_io_out_uop_stq_idx : _GEN_98 ? _slots_29_io_out_uop_stq_idx : _GEN_97 ? _slots_28_io_out_uop_stq_idx : _slots_27_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_99 ? _slots_30_io_out_uop_rxq_idx : _GEN_98 ? _slots_29_io_out_uop_rxq_idx : _GEN_97 ? _slots_28_io_out_uop_rxq_idx : _slots_27_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_99 ? _slots_30_io_out_uop_pdst : _GEN_98 ? _slots_29_io_out_uop_pdst : _GEN_97 ? _slots_28_io_out_uop_pdst : _slots_27_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_99 ? _slots_30_io_out_uop_prs1 : _GEN_98 ? _slots_29_io_out_uop_prs1 : _GEN_97 ? _slots_28_io_out_uop_prs1 : _slots_27_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_99 ? _slots_30_io_out_uop_prs2 : _GEN_98 ? _slots_29_io_out_uop_prs2 : _GEN_97 ? _slots_28_io_out_uop_prs2 : _slots_27_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_99 ? _slots_30_io_out_uop_prs3 : _GEN_98 ? _slots_29_io_out_uop_prs3 : _GEN_97 ? _slots_28_io_out_uop_prs3 : _slots_27_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_99 ? _slots_30_io_out_uop_ppred : _GEN_98 ? _slots_29_io_out_uop_ppred : _GEN_97 ? _slots_28_io_out_uop_ppred : _slots_27_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_99 ? _slots_30_io_out_uop_prs1_busy : _GEN_98 ? _slots_29_io_out_uop_prs1_busy : _GEN_97 ? _slots_28_io_out_uop_prs1_busy : _slots_27_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_99 ? _slots_30_io_out_uop_prs2_busy : _GEN_98 ? _slots_29_io_out_uop_prs2_busy : _GEN_97 ? _slots_28_io_out_uop_prs2_busy : _slots_27_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_99 ? _slots_30_io_out_uop_prs3_busy : _GEN_98 ? _slots_29_io_out_uop_prs3_busy : _GEN_97 ? _slots_28_io_out_uop_prs3_busy : _slots_27_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_99 ? _slots_30_io_out_uop_ppred_busy : _GEN_98 ? _slots_29_io_out_uop_ppred_busy : _GEN_97 ? _slots_28_io_out_uop_ppred_busy : _slots_27_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_99 ? _slots_30_io_out_uop_stale_pdst : _GEN_98 ? _slots_29_io_out_uop_stale_pdst : _GEN_97 ? _slots_28_io_out_uop_stale_pdst : _slots_27_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_99 ? _slots_30_io_out_uop_exception : _GEN_98 ? _slots_29_io_out_uop_exception : _GEN_97 ? _slots_28_io_out_uop_exception : _slots_27_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_99 ? _slots_30_io_out_uop_exc_cause : _GEN_98 ? _slots_29_io_out_uop_exc_cause : _GEN_97 ? _slots_28_io_out_uop_exc_cause : _slots_27_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_99 ? _slots_30_io_out_uop_bypassable : _GEN_98 ? _slots_29_io_out_uop_bypassable : _GEN_97 ? _slots_28_io_out_uop_bypassable : _slots_27_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_99 ? _slots_30_io_out_uop_mem_cmd : _GEN_98 ? _slots_29_io_out_uop_mem_cmd : _GEN_97 ? _slots_28_io_out_uop_mem_cmd : _slots_27_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_99 ? _slots_30_io_out_uop_mem_size : _GEN_98 ? _slots_29_io_out_uop_mem_size : _GEN_97 ? _slots_28_io_out_uop_mem_size : _slots_27_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_99 ? _slots_30_io_out_uop_mem_signed : _GEN_98 ? _slots_29_io_out_uop_mem_signed : _GEN_97 ? _slots_28_io_out_uop_mem_signed : _slots_27_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_99 ? _slots_30_io_out_uop_is_fence : _GEN_98 ? _slots_29_io_out_uop_is_fence : _GEN_97 ? _slots_28_io_out_uop_is_fence : _slots_27_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_99 ? _slots_30_io_out_uop_is_fencei : _GEN_98 ? _slots_29_io_out_uop_is_fencei : _GEN_97 ? _slots_28_io_out_uop_is_fencei : _slots_27_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_99 ? _slots_30_io_out_uop_is_amo : _GEN_98 ? _slots_29_io_out_uop_is_amo : _GEN_97 ? _slots_28_io_out_uop_is_amo : _slots_27_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_99 ? _slots_30_io_out_uop_uses_ldq : _GEN_98 ? _slots_29_io_out_uop_uses_ldq : _GEN_97 ? _slots_28_io_out_uop_uses_ldq : _slots_27_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_99 ? _slots_30_io_out_uop_uses_stq : _GEN_98 ? _slots_29_io_out_uop_uses_stq : _GEN_97 ? _slots_28_io_out_uop_uses_stq : _slots_27_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_99 ? _slots_30_io_out_uop_is_sys_pc2epc : _GEN_98 ? _slots_29_io_out_uop_is_sys_pc2epc : _GEN_97 ? _slots_28_io_out_uop_is_sys_pc2epc : _slots_27_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_99 ? _slots_30_io_out_uop_is_unique : _GEN_98 ? _slots_29_io_out_uop_is_unique : _GEN_97 ? _slots_28_io_out_uop_is_unique : _slots_27_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_99 ? _slots_30_io_out_uop_flush_on_commit : _GEN_98 ? _slots_29_io_out_uop_flush_on_commit : _GEN_97 ? _slots_28_io_out_uop_flush_on_commit : _slots_27_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_99 ? _slots_30_io_out_uop_ldst_is_rs1 : _GEN_98 ? _slots_29_io_out_uop_ldst_is_rs1 : _GEN_97 ? _slots_28_io_out_uop_ldst_is_rs1 : _slots_27_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_99 ? _slots_30_io_out_uop_ldst : _GEN_98 ? _slots_29_io_out_uop_ldst : _GEN_97 ? _slots_28_io_out_uop_ldst : _slots_27_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_99 ? _slots_30_io_out_uop_lrs1 : _GEN_98 ? _slots_29_io_out_uop_lrs1 : _GEN_97 ? _slots_28_io_out_uop_lrs1 : _slots_27_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_99 ? _slots_30_io_out_uop_lrs2 : _GEN_98 ? _slots_29_io_out_uop_lrs2 : _GEN_97 ? _slots_28_io_out_uop_lrs2 : _slots_27_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_99 ? _slots_30_io_out_uop_lrs3 : _GEN_98 ? _slots_29_io_out_uop_lrs3 : _GEN_97 ? _slots_28_io_out_uop_lrs3 : _slots_27_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_99 ? _slots_30_io_out_uop_ldst_val : _GEN_98 ? _slots_29_io_out_uop_ldst_val : _GEN_97 ? _slots_28_io_out_uop_ldst_val : _slots_27_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_99 ? _slots_30_io_out_uop_dst_rtype : _GEN_98 ? _slots_29_io_out_uop_dst_rtype : _GEN_97 ? _slots_28_io_out_uop_dst_rtype : _slots_27_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_99 ? _slots_30_io_out_uop_lrs1_rtype : _GEN_98 ? _slots_29_io_out_uop_lrs1_rtype : _GEN_97 ? _slots_28_io_out_uop_lrs1_rtype : _slots_27_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_99 ? _slots_30_io_out_uop_lrs2_rtype : _GEN_98 ? _slots_29_io_out_uop_lrs2_rtype : _GEN_97 ? _slots_28_io_out_uop_lrs2_rtype : _slots_27_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_99 ? _slots_30_io_out_uop_frs3_en : _GEN_98 ? _slots_29_io_out_uop_frs3_en : _GEN_97 ? _slots_28_io_out_uop_frs3_en : _slots_27_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_99 ? _slots_30_io_out_uop_fp_val : _GEN_98 ? _slots_29_io_out_uop_fp_val : _GEN_97 ? _slots_28_io_out_uop_fp_val : _slots_27_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_99 ? _slots_30_io_out_uop_fp_single : _GEN_98 ? _slots_29_io_out_uop_fp_single : _GEN_97 ? _slots_28_io_out_uop_fp_single : _slots_27_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_99 ? _slots_30_io_out_uop_xcpt_pf_if : _GEN_98 ? _slots_29_io_out_uop_xcpt_pf_if : _GEN_97 ? _slots_28_io_out_uop_xcpt_pf_if : _slots_27_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_99 ? _slots_30_io_out_uop_xcpt_ae_if : _GEN_98 ? _slots_29_io_out_uop_xcpt_ae_if : _GEN_97 ? _slots_28_io_out_uop_xcpt_ae_if : _slots_27_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_99 ? _slots_30_io_out_uop_xcpt_ma_if : _GEN_98 ? _slots_29_io_out_uop_xcpt_ma_if : _GEN_97 ? _slots_28_io_out_uop_xcpt_ma_if : _slots_27_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_99 ? _slots_30_io_out_uop_bp_debug_if : _GEN_98 ? _slots_29_io_out_uop_bp_debug_if : _GEN_97 ? _slots_28_io_out_uop_bp_debug_if : _slots_27_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_99 ? _slots_30_io_out_uop_bp_xcpt_if : _GEN_98 ? _slots_29_io_out_uop_bp_xcpt_if : _GEN_97 ? _slots_28_io_out_uop_bp_xcpt_if : _slots_27_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_99 ? _slots_30_io_out_uop_debug_fsrc : _GEN_98 ? _slots_29_io_out_uop_debug_fsrc : _GEN_97 ? _slots_28_io_out_uop_debug_fsrc : _slots_27_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_99 ? _slots_30_io_out_uop_debug_tsrc : _GEN_98 ? _slots_29_io_out_uop_debug_tsrc : _GEN_97 ? _slots_28_io_out_uop_debug_tsrc : _slots_27_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_26_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_26_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_26_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_26_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_26_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_26_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_26_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_26_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_26_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_26_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_26_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_26_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_26_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_26_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_26_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_26_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_26_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_26_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_26_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_26_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_26_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_26_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_26_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_26_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_26_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_26_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_26_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_26_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_26_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_26_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_26_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_26_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_26_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_26_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_26_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_26_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_26_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_26_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_26_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_26_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_26_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_26_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_26_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_26_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_26_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_26_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_26_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_26_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_26_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_26_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_26_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_26_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_26_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_26_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_26_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_26_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_26_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_26_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_26_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_26_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_26_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_26_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_26_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_26_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_26_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_26_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_26_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_26_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_26_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_26_io_uop_uopc),
    .io_uop_inst                    (_slots_26_io_uop_inst),
    .io_uop_debug_inst              (_slots_26_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_26_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_26_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_26_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_26_io_uop_fu_code),
    .io_uop_iw_state                (_slots_26_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_26_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_26_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_26_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_26_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_26_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_26_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_26_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_26_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_26_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_26_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_26_io_uop_pc_lob),
    .io_uop_taken                   (_slots_26_io_uop_taken),
    .io_uop_imm_packed              (_slots_26_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_26_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_26_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_26_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_26_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_26_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_26_io_uop_pdst),
    .io_uop_prs1                    (_slots_26_io_uop_prs1),
    .io_uop_prs2                    (_slots_26_io_uop_prs2),
    .io_uop_prs3                    (_slots_26_io_uop_prs3),
    .io_uop_ppred                   (_slots_26_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_26_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_26_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_26_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_26_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_26_io_uop_stale_pdst),
    .io_uop_exception               (_slots_26_io_uop_exception),
    .io_uop_exc_cause               (_slots_26_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_26_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_26_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_26_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_26_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_26_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_26_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_26_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_26_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_26_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_26_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_26_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_26_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_26_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_26_io_uop_ldst),
    .io_uop_lrs1                    (_slots_26_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_26_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_26_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_26_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_26_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_26_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_26_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_26_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_26_io_uop_fp_val),
    .io_uop_fp_single               (_slots_26_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_26_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_26_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_26_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_26_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_26_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_26_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_26_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_27 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_27_io_valid),
    .io_will_be_valid               (_slots_27_io_will_be_valid),
    .io_request                     (_slots_27_io_request),
    .io_grant                       (issue_slots_27_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_26),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_27_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_102 ? _slots_31_io_out_uop_uopc : _GEN_101 ? _slots_30_io_out_uop_uopc : _GEN_100 ? _slots_29_io_out_uop_uopc : _slots_28_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_102 ? _slots_31_io_out_uop_inst : _GEN_101 ? _slots_30_io_out_uop_inst : _GEN_100 ? _slots_29_io_out_uop_inst : _slots_28_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_102 ? _slots_31_io_out_uop_debug_inst : _GEN_101 ? _slots_30_io_out_uop_debug_inst : _GEN_100 ? _slots_29_io_out_uop_debug_inst : _slots_28_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_102 ? _slots_31_io_out_uop_is_rvc : _GEN_101 ? _slots_30_io_out_uop_is_rvc : _GEN_100 ? _slots_29_io_out_uop_is_rvc : _slots_28_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_102 ? _slots_31_io_out_uop_debug_pc : _GEN_101 ? _slots_30_io_out_uop_debug_pc : _GEN_100 ? _slots_29_io_out_uop_debug_pc : _slots_28_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_102 ? _slots_31_io_out_uop_iq_type : _GEN_101 ? _slots_30_io_out_uop_iq_type : _GEN_100 ? _slots_29_io_out_uop_iq_type : _slots_28_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_102 ? _slots_31_io_out_uop_fu_code : _GEN_101 ? _slots_30_io_out_uop_fu_code : _GEN_100 ? _slots_29_io_out_uop_fu_code : _slots_28_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_102 ? _slots_31_io_out_uop_iw_state : _GEN_101 ? _slots_30_io_out_uop_iw_state : _GEN_100 ? _slots_29_io_out_uop_iw_state : _slots_28_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_102 ? _slots_31_io_out_uop_iw_p1_poisoned : _GEN_101 ? _slots_30_io_out_uop_iw_p1_poisoned : _GEN_100 ? _slots_29_io_out_uop_iw_p1_poisoned : _slots_28_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_102 ? _slots_31_io_out_uop_iw_p2_poisoned : _GEN_101 ? _slots_30_io_out_uop_iw_p2_poisoned : _GEN_100 ? _slots_29_io_out_uop_iw_p2_poisoned : _slots_28_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_102 ? _slots_31_io_out_uop_is_br : _GEN_101 ? _slots_30_io_out_uop_is_br : _GEN_100 ? _slots_29_io_out_uop_is_br : _slots_28_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_102 ? _slots_31_io_out_uop_is_jalr : _GEN_101 ? _slots_30_io_out_uop_is_jalr : _GEN_100 ? _slots_29_io_out_uop_is_jalr : _slots_28_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_102 ? _slots_31_io_out_uop_is_jal : _GEN_101 ? _slots_30_io_out_uop_is_jal : _GEN_100 ? _slots_29_io_out_uop_is_jal : _slots_28_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_102 ? _slots_31_io_out_uop_is_sfb : _GEN_101 ? _slots_30_io_out_uop_is_sfb : _GEN_100 ? _slots_29_io_out_uop_is_sfb : _slots_28_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_102 ? _slots_31_io_out_uop_br_mask : _GEN_101 ? _slots_30_io_out_uop_br_mask : _GEN_100 ? _slots_29_io_out_uop_br_mask : _slots_28_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_102 ? _slots_31_io_out_uop_br_tag : _GEN_101 ? _slots_30_io_out_uop_br_tag : _GEN_100 ? _slots_29_io_out_uop_br_tag : _slots_28_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_102 ? _slots_31_io_out_uop_ftq_idx : _GEN_101 ? _slots_30_io_out_uop_ftq_idx : _GEN_100 ? _slots_29_io_out_uop_ftq_idx : _slots_28_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_102 ? _slots_31_io_out_uop_edge_inst : _GEN_101 ? _slots_30_io_out_uop_edge_inst : _GEN_100 ? _slots_29_io_out_uop_edge_inst : _slots_28_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_102 ? _slots_31_io_out_uop_pc_lob : _GEN_101 ? _slots_30_io_out_uop_pc_lob : _GEN_100 ? _slots_29_io_out_uop_pc_lob : _slots_28_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_102 ? _slots_31_io_out_uop_taken : _GEN_101 ? _slots_30_io_out_uop_taken : _GEN_100 ? _slots_29_io_out_uop_taken : _slots_28_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_102 ? _slots_31_io_out_uop_imm_packed : _GEN_101 ? _slots_30_io_out_uop_imm_packed : _GEN_100 ? _slots_29_io_out_uop_imm_packed : _slots_28_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_102 ? _slots_31_io_out_uop_csr_addr : _GEN_101 ? _slots_30_io_out_uop_csr_addr : _GEN_100 ? _slots_29_io_out_uop_csr_addr : _slots_28_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_102 ? _slots_31_io_out_uop_rob_idx : _GEN_101 ? _slots_30_io_out_uop_rob_idx : _GEN_100 ? _slots_29_io_out_uop_rob_idx : _slots_28_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_102 ? _slots_31_io_out_uop_ldq_idx : _GEN_101 ? _slots_30_io_out_uop_ldq_idx : _GEN_100 ? _slots_29_io_out_uop_ldq_idx : _slots_28_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_102 ? _slots_31_io_out_uop_stq_idx : _GEN_101 ? _slots_30_io_out_uop_stq_idx : _GEN_100 ? _slots_29_io_out_uop_stq_idx : _slots_28_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_102 ? _slots_31_io_out_uop_rxq_idx : _GEN_101 ? _slots_30_io_out_uop_rxq_idx : _GEN_100 ? _slots_29_io_out_uop_rxq_idx : _slots_28_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_102 ? _slots_31_io_out_uop_pdst : _GEN_101 ? _slots_30_io_out_uop_pdst : _GEN_100 ? _slots_29_io_out_uop_pdst : _slots_28_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_102 ? _slots_31_io_out_uop_prs1 : _GEN_101 ? _slots_30_io_out_uop_prs1 : _GEN_100 ? _slots_29_io_out_uop_prs1 : _slots_28_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_102 ? _slots_31_io_out_uop_prs2 : _GEN_101 ? _slots_30_io_out_uop_prs2 : _GEN_100 ? _slots_29_io_out_uop_prs2 : _slots_28_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_102 ? _slots_31_io_out_uop_prs3 : _GEN_101 ? _slots_30_io_out_uop_prs3 : _GEN_100 ? _slots_29_io_out_uop_prs3 : _slots_28_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_102 ? _slots_31_io_out_uop_ppred : _GEN_101 ? _slots_30_io_out_uop_ppred : _GEN_100 ? _slots_29_io_out_uop_ppred : _slots_28_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_102 ? _slots_31_io_out_uop_prs1_busy : _GEN_101 ? _slots_30_io_out_uop_prs1_busy : _GEN_100 ? _slots_29_io_out_uop_prs1_busy : _slots_28_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_102 ? _slots_31_io_out_uop_prs2_busy : _GEN_101 ? _slots_30_io_out_uop_prs2_busy : _GEN_100 ? _slots_29_io_out_uop_prs2_busy : _slots_28_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_102 ? _slots_31_io_out_uop_prs3_busy : _GEN_101 ? _slots_30_io_out_uop_prs3_busy : _GEN_100 ? _slots_29_io_out_uop_prs3_busy : _slots_28_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_102 ? _slots_31_io_out_uop_ppred_busy : _GEN_101 ? _slots_30_io_out_uop_ppred_busy : _GEN_100 ? _slots_29_io_out_uop_ppred_busy : _slots_28_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_102 ? _slots_31_io_out_uop_stale_pdst : _GEN_101 ? _slots_30_io_out_uop_stale_pdst : _GEN_100 ? _slots_29_io_out_uop_stale_pdst : _slots_28_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_102 ? _slots_31_io_out_uop_exception : _GEN_101 ? _slots_30_io_out_uop_exception : _GEN_100 ? _slots_29_io_out_uop_exception : _slots_28_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_102 ? _slots_31_io_out_uop_exc_cause : _GEN_101 ? _slots_30_io_out_uop_exc_cause : _GEN_100 ? _slots_29_io_out_uop_exc_cause : _slots_28_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_102 ? _slots_31_io_out_uop_bypassable : _GEN_101 ? _slots_30_io_out_uop_bypassable : _GEN_100 ? _slots_29_io_out_uop_bypassable : _slots_28_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_102 ? _slots_31_io_out_uop_mem_cmd : _GEN_101 ? _slots_30_io_out_uop_mem_cmd : _GEN_100 ? _slots_29_io_out_uop_mem_cmd : _slots_28_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_102 ? _slots_31_io_out_uop_mem_size : _GEN_101 ? _slots_30_io_out_uop_mem_size : _GEN_100 ? _slots_29_io_out_uop_mem_size : _slots_28_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_102 ? _slots_31_io_out_uop_mem_signed : _GEN_101 ? _slots_30_io_out_uop_mem_signed : _GEN_100 ? _slots_29_io_out_uop_mem_signed : _slots_28_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_102 ? _slots_31_io_out_uop_is_fence : _GEN_101 ? _slots_30_io_out_uop_is_fence : _GEN_100 ? _slots_29_io_out_uop_is_fence : _slots_28_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_102 ? _slots_31_io_out_uop_is_fencei : _GEN_101 ? _slots_30_io_out_uop_is_fencei : _GEN_100 ? _slots_29_io_out_uop_is_fencei : _slots_28_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_102 ? _slots_31_io_out_uop_is_amo : _GEN_101 ? _slots_30_io_out_uop_is_amo : _GEN_100 ? _slots_29_io_out_uop_is_amo : _slots_28_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_102 ? _slots_31_io_out_uop_uses_ldq : _GEN_101 ? _slots_30_io_out_uop_uses_ldq : _GEN_100 ? _slots_29_io_out_uop_uses_ldq : _slots_28_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_102 ? _slots_31_io_out_uop_uses_stq : _GEN_101 ? _slots_30_io_out_uop_uses_stq : _GEN_100 ? _slots_29_io_out_uop_uses_stq : _slots_28_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_102 ? _slots_31_io_out_uop_is_sys_pc2epc : _GEN_101 ? _slots_30_io_out_uop_is_sys_pc2epc : _GEN_100 ? _slots_29_io_out_uop_is_sys_pc2epc : _slots_28_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_102 ? _slots_31_io_out_uop_is_unique : _GEN_101 ? _slots_30_io_out_uop_is_unique : _GEN_100 ? _slots_29_io_out_uop_is_unique : _slots_28_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_102 ? _slots_31_io_out_uop_flush_on_commit : _GEN_101 ? _slots_30_io_out_uop_flush_on_commit : _GEN_100 ? _slots_29_io_out_uop_flush_on_commit : _slots_28_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_102 ? _slots_31_io_out_uop_ldst_is_rs1 : _GEN_101 ? _slots_30_io_out_uop_ldst_is_rs1 : _GEN_100 ? _slots_29_io_out_uop_ldst_is_rs1 : _slots_28_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_102 ? _slots_31_io_out_uop_ldst : _GEN_101 ? _slots_30_io_out_uop_ldst : _GEN_100 ? _slots_29_io_out_uop_ldst : _slots_28_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_102 ? _slots_31_io_out_uop_lrs1 : _GEN_101 ? _slots_30_io_out_uop_lrs1 : _GEN_100 ? _slots_29_io_out_uop_lrs1 : _slots_28_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_102 ? _slots_31_io_out_uop_lrs2 : _GEN_101 ? _slots_30_io_out_uop_lrs2 : _GEN_100 ? _slots_29_io_out_uop_lrs2 : _slots_28_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_102 ? _slots_31_io_out_uop_lrs3 : _GEN_101 ? _slots_30_io_out_uop_lrs3 : _GEN_100 ? _slots_29_io_out_uop_lrs3 : _slots_28_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_102 ? _slots_31_io_out_uop_ldst_val : _GEN_101 ? _slots_30_io_out_uop_ldst_val : _GEN_100 ? _slots_29_io_out_uop_ldst_val : _slots_28_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_102 ? _slots_31_io_out_uop_dst_rtype : _GEN_101 ? _slots_30_io_out_uop_dst_rtype : _GEN_100 ? _slots_29_io_out_uop_dst_rtype : _slots_28_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_102 ? _slots_31_io_out_uop_lrs1_rtype : _GEN_101 ? _slots_30_io_out_uop_lrs1_rtype : _GEN_100 ? _slots_29_io_out_uop_lrs1_rtype : _slots_28_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_102 ? _slots_31_io_out_uop_lrs2_rtype : _GEN_101 ? _slots_30_io_out_uop_lrs2_rtype : _GEN_100 ? _slots_29_io_out_uop_lrs2_rtype : _slots_28_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_102 ? _slots_31_io_out_uop_frs3_en : _GEN_101 ? _slots_30_io_out_uop_frs3_en : _GEN_100 ? _slots_29_io_out_uop_frs3_en : _slots_28_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_102 ? _slots_31_io_out_uop_fp_val : _GEN_101 ? _slots_30_io_out_uop_fp_val : _GEN_100 ? _slots_29_io_out_uop_fp_val : _slots_28_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_102 ? _slots_31_io_out_uop_fp_single : _GEN_101 ? _slots_30_io_out_uop_fp_single : _GEN_100 ? _slots_29_io_out_uop_fp_single : _slots_28_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_102 ? _slots_31_io_out_uop_xcpt_pf_if : _GEN_101 ? _slots_30_io_out_uop_xcpt_pf_if : _GEN_100 ? _slots_29_io_out_uop_xcpt_pf_if : _slots_28_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_102 ? _slots_31_io_out_uop_xcpt_ae_if : _GEN_101 ? _slots_30_io_out_uop_xcpt_ae_if : _GEN_100 ? _slots_29_io_out_uop_xcpt_ae_if : _slots_28_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_102 ? _slots_31_io_out_uop_xcpt_ma_if : _GEN_101 ? _slots_30_io_out_uop_xcpt_ma_if : _GEN_100 ? _slots_29_io_out_uop_xcpt_ma_if : _slots_28_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_102 ? _slots_31_io_out_uop_bp_debug_if : _GEN_101 ? _slots_30_io_out_uop_bp_debug_if : _GEN_100 ? _slots_29_io_out_uop_bp_debug_if : _slots_28_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_102 ? _slots_31_io_out_uop_bp_xcpt_if : _GEN_101 ? _slots_30_io_out_uop_bp_xcpt_if : _GEN_100 ? _slots_29_io_out_uop_bp_xcpt_if : _slots_28_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_102 ? _slots_31_io_out_uop_debug_fsrc : _GEN_101 ? _slots_30_io_out_uop_debug_fsrc : _GEN_100 ? _slots_29_io_out_uop_debug_fsrc : _slots_28_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_102 ? _slots_31_io_out_uop_debug_tsrc : _GEN_101 ? _slots_30_io_out_uop_debug_tsrc : _GEN_100 ? _slots_29_io_out_uop_debug_tsrc : _slots_28_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_27_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_27_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_27_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_27_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_27_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_27_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_27_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_27_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_27_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_27_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_27_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_27_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_27_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_27_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_27_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_27_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_27_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_27_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_27_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_27_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_27_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_27_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_27_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_27_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_27_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_27_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_27_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_27_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_27_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_27_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_27_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_27_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_27_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_27_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_27_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_27_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_27_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_27_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_27_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_27_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_27_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_27_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_27_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_27_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_27_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_27_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_27_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_27_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_27_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_27_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_27_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_27_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_27_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_27_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_27_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_27_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_27_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_27_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_27_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_27_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_27_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_27_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_27_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_27_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_27_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_27_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_27_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_27_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_27_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_27_io_uop_uopc),
    .io_uop_inst                    (_slots_27_io_uop_inst),
    .io_uop_debug_inst              (_slots_27_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_27_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_27_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_27_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_27_io_uop_fu_code),
    .io_uop_iw_state                (_slots_27_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_27_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_27_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_27_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_27_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_27_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_27_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_27_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_27_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_27_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_27_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_27_io_uop_pc_lob),
    .io_uop_taken                   (_slots_27_io_uop_taken),
    .io_uop_imm_packed              (_slots_27_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_27_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_27_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_27_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_27_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_27_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_27_io_uop_pdst),
    .io_uop_prs1                    (_slots_27_io_uop_prs1),
    .io_uop_prs2                    (_slots_27_io_uop_prs2),
    .io_uop_prs3                    (_slots_27_io_uop_prs3),
    .io_uop_ppred                   (_slots_27_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_27_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_27_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_27_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_27_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_27_io_uop_stale_pdst),
    .io_uop_exception               (_slots_27_io_uop_exception),
    .io_uop_exc_cause               (_slots_27_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_27_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_27_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_27_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_27_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_27_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_27_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_27_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_27_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_27_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_27_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_27_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_27_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_27_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_27_io_uop_ldst),
    .io_uop_lrs1                    (_slots_27_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_27_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_27_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_27_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_27_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_27_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_27_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_27_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_27_io_uop_fp_val),
    .io_uop_fp_single               (_slots_27_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_27_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_27_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_27_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_27_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_27_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_27_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_27_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_28 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_28_io_valid),
    .io_will_be_valid               (_slots_28_io_will_be_valid),
    .io_request                     (_slots_28_io_request),
    .io_grant                       (issue_slots_28_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_27),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_28_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_105 ? _slots_32_io_out_uop_uopc : _GEN_104 ? _slots_31_io_out_uop_uopc : _GEN_103 ? _slots_30_io_out_uop_uopc : _slots_29_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_105 ? _slots_32_io_out_uop_inst : _GEN_104 ? _slots_31_io_out_uop_inst : _GEN_103 ? _slots_30_io_out_uop_inst : _slots_29_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_105 ? _slots_32_io_out_uop_debug_inst : _GEN_104 ? _slots_31_io_out_uop_debug_inst : _GEN_103 ? _slots_30_io_out_uop_debug_inst : _slots_29_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_105 ? _slots_32_io_out_uop_is_rvc : _GEN_104 ? _slots_31_io_out_uop_is_rvc : _GEN_103 ? _slots_30_io_out_uop_is_rvc : _slots_29_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_105 ? _slots_32_io_out_uop_debug_pc : _GEN_104 ? _slots_31_io_out_uop_debug_pc : _GEN_103 ? _slots_30_io_out_uop_debug_pc : _slots_29_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_105 ? _slots_32_io_out_uop_iq_type : _GEN_104 ? _slots_31_io_out_uop_iq_type : _GEN_103 ? _slots_30_io_out_uop_iq_type : _slots_29_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_105 ? _slots_32_io_out_uop_fu_code : _GEN_104 ? _slots_31_io_out_uop_fu_code : _GEN_103 ? _slots_30_io_out_uop_fu_code : _slots_29_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_105 ? _slots_32_io_out_uop_iw_state : _GEN_104 ? _slots_31_io_out_uop_iw_state : _GEN_103 ? _slots_30_io_out_uop_iw_state : _slots_29_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_105 ? _slots_32_io_out_uop_iw_p1_poisoned : _GEN_104 ? _slots_31_io_out_uop_iw_p1_poisoned : _GEN_103 ? _slots_30_io_out_uop_iw_p1_poisoned : _slots_29_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_105 ? _slots_32_io_out_uop_iw_p2_poisoned : _GEN_104 ? _slots_31_io_out_uop_iw_p2_poisoned : _GEN_103 ? _slots_30_io_out_uop_iw_p2_poisoned : _slots_29_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_105 ? _slots_32_io_out_uop_is_br : _GEN_104 ? _slots_31_io_out_uop_is_br : _GEN_103 ? _slots_30_io_out_uop_is_br : _slots_29_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_105 ? _slots_32_io_out_uop_is_jalr : _GEN_104 ? _slots_31_io_out_uop_is_jalr : _GEN_103 ? _slots_30_io_out_uop_is_jalr : _slots_29_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_105 ? _slots_32_io_out_uop_is_jal : _GEN_104 ? _slots_31_io_out_uop_is_jal : _GEN_103 ? _slots_30_io_out_uop_is_jal : _slots_29_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_105 ? _slots_32_io_out_uop_is_sfb : _GEN_104 ? _slots_31_io_out_uop_is_sfb : _GEN_103 ? _slots_30_io_out_uop_is_sfb : _slots_29_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_105 ? _slots_32_io_out_uop_br_mask : _GEN_104 ? _slots_31_io_out_uop_br_mask : _GEN_103 ? _slots_30_io_out_uop_br_mask : _slots_29_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_105 ? _slots_32_io_out_uop_br_tag : _GEN_104 ? _slots_31_io_out_uop_br_tag : _GEN_103 ? _slots_30_io_out_uop_br_tag : _slots_29_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_105 ? _slots_32_io_out_uop_ftq_idx : _GEN_104 ? _slots_31_io_out_uop_ftq_idx : _GEN_103 ? _slots_30_io_out_uop_ftq_idx : _slots_29_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_105 ? _slots_32_io_out_uop_edge_inst : _GEN_104 ? _slots_31_io_out_uop_edge_inst : _GEN_103 ? _slots_30_io_out_uop_edge_inst : _slots_29_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_105 ? _slots_32_io_out_uop_pc_lob : _GEN_104 ? _slots_31_io_out_uop_pc_lob : _GEN_103 ? _slots_30_io_out_uop_pc_lob : _slots_29_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_105 ? _slots_32_io_out_uop_taken : _GEN_104 ? _slots_31_io_out_uop_taken : _GEN_103 ? _slots_30_io_out_uop_taken : _slots_29_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_105 ? _slots_32_io_out_uop_imm_packed : _GEN_104 ? _slots_31_io_out_uop_imm_packed : _GEN_103 ? _slots_30_io_out_uop_imm_packed : _slots_29_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_105 ? _slots_32_io_out_uop_csr_addr : _GEN_104 ? _slots_31_io_out_uop_csr_addr : _GEN_103 ? _slots_30_io_out_uop_csr_addr : _slots_29_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_105 ? _slots_32_io_out_uop_rob_idx : _GEN_104 ? _slots_31_io_out_uop_rob_idx : _GEN_103 ? _slots_30_io_out_uop_rob_idx : _slots_29_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_105 ? _slots_32_io_out_uop_ldq_idx : _GEN_104 ? _slots_31_io_out_uop_ldq_idx : _GEN_103 ? _slots_30_io_out_uop_ldq_idx : _slots_29_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_105 ? _slots_32_io_out_uop_stq_idx : _GEN_104 ? _slots_31_io_out_uop_stq_idx : _GEN_103 ? _slots_30_io_out_uop_stq_idx : _slots_29_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_105 ? _slots_32_io_out_uop_rxq_idx : _GEN_104 ? _slots_31_io_out_uop_rxq_idx : _GEN_103 ? _slots_30_io_out_uop_rxq_idx : _slots_29_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_105 ? _slots_32_io_out_uop_pdst : _GEN_104 ? _slots_31_io_out_uop_pdst : _GEN_103 ? _slots_30_io_out_uop_pdst : _slots_29_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_105 ? _slots_32_io_out_uop_prs1 : _GEN_104 ? _slots_31_io_out_uop_prs1 : _GEN_103 ? _slots_30_io_out_uop_prs1 : _slots_29_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_105 ? _slots_32_io_out_uop_prs2 : _GEN_104 ? _slots_31_io_out_uop_prs2 : _GEN_103 ? _slots_30_io_out_uop_prs2 : _slots_29_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_105 ? _slots_32_io_out_uop_prs3 : _GEN_104 ? _slots_31_io_out_uop_prs3 : _GEN_103 ? _slots_30_io_out_uop_prs3 : _slots_29_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_105 ? _slots_32_io_out_uop_ppred : _GEN_104 ? _slots_31_io_out_uop_ppred : _GEN_103 ? _slots_30_io_out_uop_ppred : _slots_29_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_105 ? _slots_32_io_out_uop_prs1_busy : _GEN_104 ? _slots_31_io_out_uop_prs1_busy : _GEN_103 ? _slots_30_io_out_uop_prs1_busy : _slots_29_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_105 ? _slots_32_io_out_uop_prs2_busy : _GEN_104 ? _slots_31_io_out_uop_prs2_busy : _GEN_103 ? _slots_30_io_out_uop_prs2_busy : _slots_29_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_105 ? _slots_32_io_out_uop_prs3_busy : _GEN_104 ? _slots_31_io_out_uop_prs3_busy : _GEN_103 ? _slots_30_io_out_uop_prs3_busy : _slots_29_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_105 ? _slots_32_io_out_uop_ppred_busy : _GEN_104 ? _slots_31_io_out_uop_ppred_busy : _GEN_103 ? _slots_30_io_out_uop_ppred_busy : _slots_29_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_105 ? _slots_32_io_out_uop_stale_pdst : _GEN_104 ? _slots_31_io_out_uop_stale_pdst : _GEN_103 ? _slots_30_io_out_uop_stale_pdst : _slots_29_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_105 ? _slots_32_io_out_uop_exception : _GEN_104 ? _slots_31_io_out_uop_exception : _GEN_103 ? _slots_30_io_out_uop_exception : _slots_29_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_105 ? _slots_32_io_out_uop_exc_cause : _GEN_104 ? _slots_31_io_out_uop_exc_cause : _GEN_103 ? _slots_30_io_out_uop_exc_cause : _slots_29_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_105 ? _slots_32_io_out_uop_bypassable : _GEN_104 ? _slots_31_io_out_uop_bypassable : _GEN_103 ? _slots_30_io_out_uop_bypassable : _slots_29_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_105 ? _slots_32_io_out_uop_mem_cmd : _GEN_104 ? _slots_31_io_out_uop_mem_cmd : _GEN_103 ? _slots_30_io_out_uop_mem_cmd : _slots_29_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_105 ? _slots_32_io_out_uop_mem_size : _GEN_104 ? _slots_31_io_out_uop_mem_size : _GEN_103 ? _slots_30_io_out_uop_mem_size : _slots_29_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_105 ? _slots_32_io_out_uop_mem_signed : _GEN_104 ? _slots_31_io_out_uop_mem_signed : _GEN_103 ? _slots_30_io_out_uop_mem_signed : _slots_29_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_105 ? _slots_32_io_out_uop_is_fence : _GEN_104 ? _slots_31_io_out_uop_is_fence : _GEN_103 ? _slots_30_io_out_uop_is_fence : _slots_29_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_105 ? _slots_32_io_out_uop_is_fencei : _GEN_104 ? _slots_31_io_out_uop_is_fencei : _GEN_103 ? _slots_30_io_out_uop_is_fencei : _slots_29_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_105 ? _slots_32_io_out_uop_is_amo : _GEN_104 ? _slots_31_io_out_uop_is_amo : _GEN_103 ? _slots_30_io_out_uop_is_amo : _slots_29_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_105 ? _slots_32_io_out_uop_uses_ldq : _GEN_104 ? _slots_31_io_out_uop_uses_ldq : _GEN_103 ? _slots_30_io_out_uop_uses_ldq : _slots_29_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_105 ? _slots_32_io_out_uop_uses_stq : _GEN_104 ? _slots_31_io_out_uop_uses_stq : _GEN_103 ? _slots_30_io_out_uop_uses_stq : _slots_29_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_105 ? _slots_32_io_out_uop_is_sys_pc2epc : _GEN_104 ? _slots_31_io_out_uop_is_sys_pc2epc : _GEN_103 ? _slots_30_io_out_uop_is_sys_pc2epc : _slots_29_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_105 ? _slots_32_io_out_uop_is_unique : _GEN_104 ? _slots_31_io_out_uop_is_unique : _GEN_103 ? _slots_30_io_out_uop_is_unique : _slots_29_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_105 ? _slots_32_io_out_uop_flush_on_commit : _GEN_104 ? _slots_31_io_out_uop_flush_on_commit : _GEN_103 ? _slots_30_io_out_uop_flush_on_commit : _slots_29_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_105 ? _slots_32_io_out_uop_ldst_is_rs1 : _GEN_104 ? _slots_31_io_out_uop_ldst_is_rs1 : _GEN_103 ? _slots_30_io_out_uop_ldst_is_rs1 : _slots_29_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_105 ? _slots_32_io_out_uop_ldst : _GEN_104 ? _slots_31_io_out_uop_ldst : _GEN_103 ? _slots_30_io_out_uop_ldst : _slots_29_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_105 ? _slots_32_io_out_uop_lrs1 : _GEN_104 ? _slots_31_io_out_uop_lrs1 : _GEN_103 ? _slots_30_io_out_uop_lrs1 : _slots_29_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_105 ? _slots_32_io_out_uop_lrs2 : _GEN_104 ? _slots_31_io_out_uop_lrs2 : _GEN_103 ? _slots_30_io_out_uop_lrs2 : _slots_29_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_105 ? _slots_32_io_out_uop_lrs3 : _GEN_104 ? _slots_31_io_out_uop_lrs3 : _GEN_103 ? _slots_30_io_out_uop_lrs3 : _slots_29_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_105 ? _slots_32_io_out_uop_ldst_val : _GEN_104 ? _slots_31_io_out_uop_ldst_val : _GEN_103 ? _slots_30_io_out_uop_ldst_val : _slots_29_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_105 ? _slots_32_io_out_uop_dst_rtype : _GEN_104 ? _slots_31_io_out_uop_dst_rtype : _GEN_103 ? _slots_30_io_out_uop_dst_rtype : _slots_29_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_105 ? _slots_32_io_out_uop_lrs1_rtype : _GEN_104 ? _slots_31_io_out_uop_lrs1_rtype : _GEN_103 ? _slots_30_io_out_uop_lrs1_rtype : _slots_29_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_105 ? _slots_32_io_out_uop_lrs2_rtype : _GEN_104 ? _slots_31_io_out_uop_lrs2_rtype : _GEN_103 ? _slots_30_io_out_uop_lrs2_rtype : _slots_29_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_105 ? _slots_32_io_out_uop_frs3_en : _GEN_104 ? _slots_31_io_out_uop_frs3_en : _GEN_103 ? _slots_30_io_out_uop_frs3_en : _slots_29_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_105 ? _slots_32_io_out_uop_fp_val : _GEN_104 ? _slots_31_io_out_uop_fp_val : _GEN_103 ? _slots_30_io_out_uop_fp_val : _slots_29_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_105 ? _slots_32_io_out_uop_fp_single : _GEN_104 ? _slots_31_io_out_uop_fp_single : _GEN_103 ? _slots_30_io_out_uop_fp_single : _slots_29_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_105 ? _slots_32_io_out_uop_xcpt_pf_if : _GEN_104 ? _slots_31_io_out_uop_xcpt_pf_if : _GEN_103 ? _slots_30_io_out_uop_xcpt_pf_if : _slots_29_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_105 ? _slots_32_io_out_uop_xcpt_ae_if : _GEN_104 ? _slots_31_io_out_uop_xcpt_ae_if : _GEN_103 ? _slots_30_io_out_uop_xcpt_ae_if : _slots_29_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_105 ? _slots_32_io_out_uop_xcpt_ma_if : _GEN_104 ? _slots_31_io_out_uop_xcpt_ma_if : _GEN_103 ? _slots_30_io_out_uop_xcpt_ma_if : _slots_29_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_105 ? _slots_32_io_out_uop_bp_debug_if : _GEN_104 ? _slots_31_io_out_uop_bp_debug_if : _GEN_103 ? _slots_30_io_out_uop_bp_debug_if : _slots_29_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_105 ? _slots_32_io_out_uop_bp_xcpt_if : _GEN_104 ? _slots_31_io_out_uop_bp_xcpt_if : _GEN_103 ? _slots_30_io_out_uop_bp_xcpt_if : _slots_29_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_105 ? _slots_32_io_out_uop_debug_fsrc : _GEN_104 ? _slots_31_io_out_uop_debug_fsrc : _GEN_103 ? _slots_30_io_out_uop_debug_fsrc : _slots_29_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_105 ? _slots_32_io_out_uop_debug_tsrc : _GEN_104 ? _slots_31_io_out_uop_debug_tsrc : _GEN_103 ? _slots_30_io_out_uop_debug_tsrc : _slots_29_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_28_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_28_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_28_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_28_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_28_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_28_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_28_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_28_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_28_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_28_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_28_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_28_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_28_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_28_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_28_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_28_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_28_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_28_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_28_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_28_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_28_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_28_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_28_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_28_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_28_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_28_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_28_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_28_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_28_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_28_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_28_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_28_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_28_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_28_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_28_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_28_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_28_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_28_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_28_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_28_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_28_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_28_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_28_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_28_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_28_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_28_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_28_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_28_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_28_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_28_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_28_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_28_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_28_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_28_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_28_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_28_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_28_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_28_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_28_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_28_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_28_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_28_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_28_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_28_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_28_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_28_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_28_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_28_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_28_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_28_io_uop_uopc),
    .io_uop_inst                    (_slots_28_io_uop_inst),
    .io_uop_debug_inst              (_slots_28_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_28_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_28_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_28_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_28_io_uop_fu_code),
    .io_uop_iw_state                (_slots_28_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_28_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_28_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_28_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_28_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_28_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_28_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_28_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_28_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_28_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_28_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_28_io_uop_pc_lob),
    .io_uop_taken                   (_slots_28_io_uop_taken),
    .io_uop_imm_packed              (_slots_28_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_28_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_28_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_28_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_28_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_28_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_28_io_uop_pdst),
    .io_uop_prs1                    (_slots_28_io_uop_prs1),
    .io_uop_prs2                    (_slots_28_io_uop_prs2),
    .io_uop_prs3                    (_slots_28_io_uop_prs3),
    .io_uop_ppred                   (_slots_28_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_28_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_28_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_28_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_28_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_28_io_uop_stale_pdst),
    .io_uop_exception               (_slots_28_io_uop_exception),
    .io_uop_exc_cause               (_slots_28_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_28_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_28_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_28_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_28_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_28_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_28_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_28_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_28_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_28_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_28_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_28_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_28_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_28_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_28_io_uop_ldst),
    .io_uop_lrs1                    (_slots_28_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_28_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_28_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_28_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_28_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_28_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_28_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_28_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_28_io_uop_fp_val),
    .io_uop_fp_single               (_slots_28_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_28_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_28_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_28_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_28_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_28_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_28_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_28_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_29 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_29_io_valid),
    .io_will_be_valid               (_slots_29_io_will_be_valid),
    .io_request                     (_slots_29_io_request),
    .io_grant                       (issue_slots_29_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_28),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_29_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_108 ? _slots_33_io_out_uop_uopc : _GEN_107 ? _slots_32_io_out_uop_uopc : _GEN_106 ? _slots_31_io_out_uop_uopc : _slots_30_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_108 ? _slots_33_io_out_uop_inst : _GEN_107 ? _slots_32_io_out_uop_inst : _GEN_106 ? _slots_31_io_out_uop_inst : _slots_30_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_108 ? _slots_33_io_out_uop_debug_inst : _GEN_107 ? _slots_32_io_out_uop_debug_inst : _GEN_106 ? _slots_31_io_out_uop_debug_inst : _slots_30_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_108 ? _slots_33_io_out_uop_is_rvc : _GEN_107 ? _slots_32_io_out_uop_is_rvc : _GEN_106 ? _slots_31_io_out_uop_is_rvc : _slots_30_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_108 ? _slots_33_io_out_uop_debug_pc : _GEN_107 ? _slots_32_io_out_uop_debug_pc : _GEN_106 ? _slots_31_io_out_uop_debug_pc : _slots_30_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_108 ? _slots_33_io_out_uop_iq_type : _GEN_107 ? _slots_32_io_out_uop_iq_type : _GEN_106 ? _slots_31_io_out_uop_iq_type : _slots_30_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_108 ? _slots_33_io_out_uop_fu_code : _GEN_107 ? _slots_32_io_out_uop_fu_code : _GEN_106 ? _slots_31_io_out_uop_fu_code : _slots_30_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_108 ? _slots_33_io_out_uop_iw_state : _GEN_107 ? _slots_32_io_out_uop_iw_state : _GEN_106 ? _slots_31_io_out_uop_iw_state : _slots_30_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_108 ? _slots_33_io_out_uop_iw_p1_poisoned : _GEN_107 ? _slots_32_io_out_uop_iw_p1_poisoned : _GEN_106 ? _slots_31_io_out_uop_iw_p1_poisoned : _slots_30_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_108 ? _slots_33_io_out_uop_iw_p2_poisoned : _GEN_107 ? _slots_32_io_out_uop_iw_p2_poisoned : _GEN_106 ? _slots_31_io_out_uop_iw_p2_poisoned : _slots_30_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_108 ? _slots_33_io_out_uop_is_br : _GEN_107 ? _slots_32_io_out_uop_is_br : _GEN_106 ? _slots_31_io_out_uop_is_br : _slots_30_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_108 ? _slots_33_io_out_uop_is_jalr : _GEN_107 ? _slots_32_io_out_uop_is_jalr : _GEN_106 ? _slots_31_io_out_uop_is_jalr : _slots_30_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_108 ? _slots_33_io_out_uop_is_jal : _GEN_107 ? _slots_32_io_out_uop_is_jal : _GEN_106 ? _slots_31_io_out_uop_is_jal : _slots_30_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_108 ? _slots_33_io_out_uop_is_sfb : _GEN_107 ? _slots_32_io_out_uop_is_sfb : _GEN_106 ? _slots_31_io_out_uop_is_sfb : _slots_30_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_108 ? _slots_33_io_out_uop_br_mask : _GEN_107 ? _slots_32_io_out_uop_br_mask : _GEN_106 ? _slots_31_io_out_uop_br_mask : _slots_30_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_108 ? _slots_33_io_out_uop_br_tag : _GEN_107 ? _slots_32_io_out_uop_br_tag : _GEN_106 ? _slots_31_io_out_uop_br_tag : _slots_30_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_108 ? _slots_33_io_out_uop_ftq_idx : _GEN_107 ? _slots_32_io_out_uop_ftq_idx : _GEN_106 ? _slots_31_io_out_uop_ftq_idx : _slots_30_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_108 ? _slots_33_io_out_uop_edge_inst : _GEN_107 ? _slots_32_io_out_uop_edge_inst : _GEN_106 ? _slots_31_io_out_uop_edge_inst : _slots_30_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_108 ? _slots_33_io_out_uop_pc_lob : _GEN_107 ? _slots_32_io_out_uop_pc_lob : _GEN_106 ? _slots_31_io_out_uop_pc_lob : _slots_30_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_108 ? _slots_33_io_out_uop_taken : _GEN_107 ? _slots_32_io_out_uop_taken : _GEN_106 ? _slots_31_io_out_uop_taken : _slots_30_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_108 ? _slots_33_io_out_uop_imm_packed : _GEN_107 ? _slots_32_io_out_uop_imm_packed : _GEN_106 ? _slots_31_io_out_uop_imm_packed : _slots_30_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_108 ? _slots_33_io_out_uop_csr_addr : _GEN_107 ? _slots_32_io_out_uop_csr_addr : _GEN_106 ? _slots_31_io_out_uop_csr_addr : _slots_30_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_108 ? _slots_33_io_out_uop_rob_idx : _GEN_107 ? _slots_32_io_out_uop_rob_idx : _GEN_106 ? _slots_31_io_out_uop_rob_idx : _slots_30_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_108 ? _slots_33_io_out_uop_ldq_idx : _GEN_107 ? _slots_32_io_out_uop_ldq_idx : _GEN_106 ? _slots_31_io_out_uop_ldq_idx : _slots_30_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_108 ? _slots_33_io_out_uop_stq_idx : _GEN_107 ? _slots_32_io_out_uop_stq_idx : _GEN_106 ? _slots_31_io_out_uop_stq_idx : _slots_30_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_108 ? _slots_33_io_out_uop_rxq_idx : _GEN_107 ? _slots_32_io_out_uop_rxq_idx : _GEN_106 ? _slots_31_io_out_uop_rxq_idx : _slots_30_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_108 ? _slots_33_io_out_uop_pdst : _GEN_107 ? _slots_32_io_out_uop_pdst : _GEN_106 ? _slots_31_io_out_uop_pdst : _slots_30_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_108 ? _slots_33_io_out_uop_prs1 : _GEN_107 ? _slots_32_io_out_uop_prs1 : _GEN_106 ? _slots_31_io_out_uop_prs1 : _slots_30_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_108 ? _slots_33_io_out_uop_prs2 : _GEN_107 ? _slots_32_io_out_uop_prs2 : _GEN_106 ? _slots_31_io_out_uop_prs2 : _slots_30_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_108 ? _slots_33_io_out_uop_prs3 : _GEN_107 ? _slots_32_io_out_uop_prs3 : _GEN_106 ? _slots_31_io_out_uop_prs3 : _slots_30_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_108 ? _slots_33_io_out_uop_ppred : _GEN_107 ? _slots_32_io_out_uop_ppred : _GEN_106 ? _slots_31_io_out_uop_ppred : _slots_30_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_108 ? _slots_33_io_out_uop_prs1_busy : _GEN_107 ? _slots_32_io_out_uop_prs1_busy : _GEN_106 ? _slots_31_io_out_uop_prs1_busy : _slots_30_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_108 ? _slots_33_io_out_uop_prs2_busy : _GEN_107 ? _slots_32_io_out_uop_prs2_busy : _GEN_106 ? _slots_31_io_out_uop_prs2_busy : _slots_30_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_108 ? _slots_33_io_out_uop_prs3_busy : _GEN_107 ? _slots_32_io_out_uop_prs3_busy : _GEN_106 ? _slots_31_io_out_uop_prs3_busy : _slots_30_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_108 ? _slots_33_io_out_uop_ppred_busy : _GEN_107 ? _slots_32_io_out_uop_ppred_busy : _GEN_106 ? _slots_31_io_out_uop_ppred_busy : _slots_30_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_108 ? _slots_33_io_out_uop_stale_pdst : _GEN_107 ? _slots_32_io_out_uop_stale_pdst : _GEN_106 ? _slots_31_io_out_uop_stale_pdst : _slots_30_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_108 ? _slots_33_io_out_uop_exception : _GEN_107 ? _slots_32_io_out_uop_exception : _GEN_106 ? _slots_31_io_out_uop_exception : _slots_30_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_108 ? _slots_33_io_out_uop_exc_cause : _GEN_107 ? _slots_32_io_out_uop_exc_cause : _GEN_106 ? _slots_31_io_out_uop_exc_cause : _slots_30_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_108 ? _slots_33_io_out_uop_bypassable : _GEN_107 ? _slots_32_io_out_uop_bypassable : _GEN_106 ? _slots_31_io_out_uop_bypassable : _slots_30_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_108 ? _slots_33_io_out_uop_mem_cmd : _GEN_107 ? _slots_32_io_out_uop_mem_cmd : _GEN_106 ? _slots_31_io_out_uop_mem_cmd : _slots_30_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_108 ? _slots_33_io_out_uop_mem_size : _GEN_107 ? _slots_32_io_out_uop_mem_size : _GEN_106 ? _slots_31_io_out_uop_mem_size : _slots_30_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_108 ? _slots_33_io_out_uop_mem_signed : _GEN_107 ? _slots_32_io_out_uop_mem_signed : _GEN_106 ? _slots_31_io_out_uop_mem_signed : _slots_30_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_108 ? _slots_33_io_out_uop_is_fence : _GEN_107 ? _slots_32_io_out_uop_is_fence : _GEN_106 ? _slots_31_io_out_uop_is_fence : _slots_30_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_108 ? _slots_33_io_out_uop_is_fencei : _GEN_107 ? _slots_32_io_out_uop_is_fencei : _GEN_106 ? _slots_31_io_out_uop_is_fencei : _slots_30_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_108 ? _slots_33_io_out_uop_is_amo : _GEN_107 ? _slots_32_io_out_uop_is_amo : _GEN_106 ? _slots_31_io_out_uop_is_amo : _slots_30_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_108 ? _slots_33_io_out_uop_uses_ldq : _GEN_107 ? _slots_32_io_out_uop_uses_ldq : _GEN_106 ? _slots_31_io_out_uop_uses_ldq : _slots_30_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_108 ? _slots_33_io_out_uop_uses_stq : _GEN_107 ? _slots_32_io_out_uop_uses_stq : _GEN_106 ? _slots_31_io_out_uop_uses_stq : _slots_30_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_108 ? _slots_33_io_out_uop_is_sys_pc2epc : _GEN_107 ? _slots_32_io_out_uop_is_sys_pc2epc : _GEN_106 ? _slots_31_io_out_uop_is_sys_pc2epc : _slots_30_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_108 ? _slots_33_io_out_uop_is_unique : _GEN_107 ? _slots_32_io_out_uop_is_unique : _GEN_106 ? _slots_31_io_out_uop_is_unique : _slots_30_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_108 ? _slots_33_io_out_uop_flush_on_commit : _GEN_107 ? _slots_32_io_out_uop_flush_on_commit : _GEN_106 ? _slots_31_io_out_uop_flush_on_commit : _slots_30_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_108 ? _slots_33_io_out_uop_ldst_is_rs1 : _GEN_107 ? _slots_32_io_out_uop_ldst_is_rs1 : _GEN_106 ? _slots_31_io_out_uop_ldst_is_rs1 : _slots_30_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_108 ? _slots_33_io_out_uop_ldst : _GEN_107 ? _slots_32_io_out_uop_ldst : _GEN_106 ? _slots_31_io_out_uop_ldst : _slots_30_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_108 ? _slots_33_io_out_uop_lrs1 : _GEN_107 ? _slots_32_io_out_uop_lrs1 : _GEN_106 ? _slots_31_io_out_uop_lrs1 : _slots_30_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_108 ? _slots_33_io_out_uop_lrs2 : _GEN_107 ? _slots_32_io_out_uop_lrs2 : _GEN_106 ? _slots_31_io_out_uop_lrs2 : _slots_30_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_108 ? _slots_33_io_out_uop_lrs3 : _GEN_107 ? _slots_32_io_out_uop_lrs3 : _GEN_106 ? _slots_31_io_out_uop_lrs3 : _slots_30_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_108 ? _slots_33_io_out_uop_ldst_val : _GEN_107 ? _slots_32_io_out_uop_ldst_val : _GEN_106 ? _slots_31_io_out_uop_ldst_val : _slots_30_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_108 ? _slots_33_io_out_uop_dst_rtype : _GEN_107 ? _slots_32_io_out_uop_dst_rtype : _GEN_106 ? _slots_31_io_out_uop_dst_rtype : _slots_30_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_108 ? _slots_33_io_out_uop_lrs1_rtype : _GEN_107 ? _slots_32_io_out_uop_lrs1_rtype : _GEN_106 ? _slots_31_io_out_uop_lrs1_rtype : _slots_30_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_108 ? _slots_33_io_out_uop_lrs2_rtype : _GEN_107 ? _slots_32_io_out_uop_lrs2_rtype : _GEN_106 ? _slots_31_io_out_uop_lrs2_rtype : _slots_30_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_108 ? _slots_33_io_out_uop_frs3_en : _GEN_107 ? _slots_32_io_out_uop_frs3_en : _GEN_106 ? _slots_31_io_out_uop_frs3_en : _slots_30_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_108 ? _slots_33_io_out_uop_fp_val : _GEN_107 ? _slots_32_io_out_uop_fp_val : _GEN_106 ? _slots_31_io_out_uop_fp_val : _slots_30_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_108 ? _slots_33_io_out_uop_fp_single : _GEN_107 ? _slots_32_io_out_uop_fp_single : _GEN_106 ? _slots_31_io_out_uop_fp_single : _slots_30_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_108 ? _slots_33_io_out_uop_xcpt_pf_if : _GEN_107 ? _slots_32_io_out_uop_xcpt_pf_if : _GEN_106 ? _slots_31_io_out_uop_xcpt_pf_if : _slots_30_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_108 ? _slots_33_io_out_uop_xcpt_ae_if : _GEN_107 ? _slots_32_io_out_uop_xcpt_ae_if : _GEN_106 ? _slots_31_io_out_uop_xcpt_ae_if : _slots_30_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_108 ? _slots_33_io_out_uop_xcpt_ma_if : _GEN_107 ? _slots_32_io_out_uop_xcpt_ma_if : _GEN_106 ? _slots_31_io_out_uop_xcpt_ma_if : _slots_30_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_108 ? _slots_33_io_out_uop_bp_debug_if : _GEN_107 ? _slots_32_io_out_uop_bp_debug_if : _GEN_106 ? _slots_31_io_out_uop_bp_debug_if : _slots_30_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_108 ? _slots_33_io_out_uop_bp_xcpt_if : _GEN_107 ? _slots_32_io_out_uop_bp_xcpt_if : _GEN_106 ? _slots_31_io_out_uop_bp_xcpt_if : _slots_30_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_108 ? _slots_33_io_out_uop_debug_fsrc : _GEN_107 ? _slots_32_io_out_uop_debug_fsrc : _GEN_106 ? _slots_31_io_out_uop_debug_fsrc : _slots_30_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_108 ? _slots_33_io_out_uop_debug_tsrc : _GEN_107 ? _slots_32_io_out_uop_debug_tsrc : _GEN_106 ? _slots_31_io_out_uop_debug_tsrc : _slots_30_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_29_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_29_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_29_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_29_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_29_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_29_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_29_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_29_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_29_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_29_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_29_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_29_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_29_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_29_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_29_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_29_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_29_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_29_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_29_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_29_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_29_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_29_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_29_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_29_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_29_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_29_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_29_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_29_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_29_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_29_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_29_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_29_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_29_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_29_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_29_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_29_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_29_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_29_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_29_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_29_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_29_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_29_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_29_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_29_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_29_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_29_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_29_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_29_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_29_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_29_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_29_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_29_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_29_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_29_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_29_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_29_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_29_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_29_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_29_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_29_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_29_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_29_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_29_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_29_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_29_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_29_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_29_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_29_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_29_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_29_io_uop_uopc),
    .io_uop_inst                    (_slots_29_io_uop_inst),
    .io_uop_debug_inst              (_slots_29_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_29_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_29_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_29_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_29_io_uop_fu_code),
    .io_uop_iw_state                (_slots_29_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_29_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_29_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_29_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_29_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_29_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_29_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_29_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_29_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_29_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_29_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_29_io_uop_pc_lob),
    .io_uop_taken                   (_slots_29_io_uop_taken),
    .io_uop_imm_packed              (_slots_29_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_29_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_29_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_29_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_29_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_29_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_29_io_uop_pdst),
    .io_uop_prs1                    (_slots_29_io_uop_prs1),
    .io_uop_prs2                    (_slots_29_io_uop_prs2),
    .io_uop_prs3                    (_slots_29_io_uop_prs3),
    .io_uop_ppred                   (_slots_29_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_29_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_29_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_29_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_29_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_29_io_uop_stale_pdst),
    .io_uop_exception               (_slots_29_io_uop_exception),
    .io_uop_exc_cause               (_slots_29_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_29_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_29_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_29_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_29_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_29_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_29_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_29_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_29_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_29_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_29_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_29_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_29_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_29_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_29_io_uop_ldst),
    .io_uop_lrs1                    (_slots_29_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_29_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_29_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_29_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_29_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_29_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_29_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_29_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_29_io_uop_fp_val),
    .io_uop_fp_single               (_slots_29_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_29_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_29_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_29_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_29_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_29_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_29_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_29_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_30 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_30_io_valid),
    .io_will_be_valid               (_slots_30_io_will_be_valid),
    .io_request                     (_slots_30_io_request),
    .io_grant                       (issue_slots_30_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_29),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_30_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_111 ? _slots_34_io_out_uop_uopc : _GEN_110 ? _slots_33_io_out_uop_uopc : _GEN_109 ? _slots_32_io_out_uop_uopc : _slots_31_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_111 ? _slots_34_io_out_uop_inst : _GEN_110 ? _slots_33_io_out_uop_inst : _GEN_109 ? _slots_32_io_out_uop_inst : _slots_31_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_111 ? _slots_34_io_out_uop_debug_inst : _GEN_110 ? _slots_33_io_out_uop_debug_inst : _GEN_109 ? _slots_32_io_out_uop_debug_inst : _slots_31_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_111 ? _slots_34_io_out_uop_is_rvc : _GEN_110 ? _slots_33_io_out_uop_is_rvc : _GEN_109 ? _slots_32_io_out_uop_is_rvc : _slots_31_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_111 ? _slots_34_io_out_uop_debug_pc : _GEN_110 ? _slots_33_io_out_uop_debug_pc : _GEN_109 ? _slots_32_io_out_uop_debug_pc : _slots_31_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_111 ? _slots_34_io_out_uop_iq_type : _GEN_110 ? _slots_33_io_out_uop_iq_type : _GEN_109 ? _slots_32_io_out_uop_iq_type : _slots_31_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_111 ? _slots_34_io_out_uop_fu_code : _GEN_110 ? _slots_33_io_out_uop_fu_code : _GEN_109 ? _slots_32_io_out_uop_fu_code : _slots_31_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_111 ? _slots_34_io_out_uop_iw_state : _GEN_110 ? _slots_33_io_out_uop_iw_state : _GEN_109 ? _slots_32_io_out_uop_iw_state : _slots_31_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_111 ? _slots_34_io_out_uop_iw_p1_poisoned : _GEN_110 ? _slots_33_io_out_uop_iw_p1_poisoned : _GEN_109 ? _slots_32_io_out_uop_iw_p1_poisoned : _slots_31_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_111 ? _slots_34_io_out_uop_iw_p2_poisoned : _GEN_110 ? _slots_33_io_out_uop_iw_p2_poisoned : _GEN_109 ? _slots_32_io_out_uop_iw_p2_poisoned : _slots_31_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_111 ? _slots_34_io_out_uop_is_br : _GEN_110 ? _slots_33_io_out_uop_is_br : _GEN_109 ? _slots_32_io_out_uop_is_br : _slots_31_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_111 ? _slots_34_io_out_uop_is_jalr : _GEN_110 ? _slots_33_io_out_uop_is_jalr : _GEN_109 ? _slots_32_io_out_uop_is_jalr : _slots_31_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_111 ? _slots_34_io_out_uop_is_jal : _GEN_110 ? _slots_33_io_out_uop_is_jal : _GEN_109 ? _slots_32_io_out_uop_is_jal : _slots_31_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_111 ? _slots_34_io_out_uop_is_sfb : _GEN_110 ? _slots_33_io_out_uop_is_sfb : _GEN_109 ? _slots_32_io_out_uop_is_sfb : _slots_31_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_111 ? _slots_34_io_out_uop_br_mask : _GEN_110 ? _slots_33_io_out_uop_br_mask : _GEN_109 ? _slots_32_io_out_uop_br_mask : _slots_31_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_111 ? _slots_34_io_out_uop_br_tag : _GEN_110 ? _slots_33_io_out_uop_br_tag : _GEN_109 ? _slots_32_io_out_uop_br_tag : _slots_31_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_111 ? _slots_34_io_out_uop_ftq_idx : _GEN_110 ? _slots_33_io_out_uop_ftq_idx : _GEN_109 ? _slots_32_io_out_uop_ftq_idx : _slots_31_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_111 ? _slots_34_io_out_uop_edge_inst : _GEN_110 ? _slots_33_io_out_uop_edge_inst : _GEN_109 ? _slots_32_io_out_uop_edge_inst : _slots_31_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_111 ? _slots_34_io_out_uop_pc_lob : _GEN_110 ? _slots_33_io_out_uop_pc_lob : _GEN_109 ? _slots_32_io_out_uop_pc_lob : _slots_31_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_111 ? _slots_34_io_out_uop_taken : _GEN_110 ? _slots_33_io_out_uop_taken : _GEN_109 ? _slots_32_io_out_uop_taken : _slots_31_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_111 ? _slots_34_io_out_uop_imm_packed : _GEN_110 ? _slots_33_io_out_uop_imm_packed : _GEN_109 ? _slots_32_io_out_uop_imm_packed : _slots_31_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_111 ? _slots_34_io_out_uop_csr_addr : _GEN_110 ? _slots_33_io_out_uop_csr_addr : _GEN_109 ? _slots_32_io_out_uop_csr_addr : _slots_31_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_111 ? _slots_34_io_out_uop_rob_idx : _GEN_110 ? _slots_33_io_out_uop_rob_idx : _GEN_109 ? _slots_32_io_out_uop_rob_idx : _slots_31_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_111 ? _slots_34_io_out_uop_ldq_idx : _GEN_110 ? _slots_33_io_out_uop_ldq_idx : _GEN_109 ? _slots_32_io_out_uop_ldq_idx : _slots_31_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_111 ? _slots_34_io_out_uop_stq_idx : _GEN_110 ? _slots_33_io_out_uop_stq_idx : _GEN_109 ? _slots_32_io_out_uop_stq_idx : _slots_31_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_111 ? _slots_34_io_out_uop_rxq_idx : _GEN_110 ? _slots_33_io_out_uop_rxq_idx : _GEN_109 ? _slots_32_io_out_uop_rxq_idx : _slots_31_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_111 ? _slots_34_io_out_uop_pdst : _GEN_110 ? _slots_33_io_out_uop_pdst : _GEN_109 ? _slots_32_io_out_uop_pdst : _slots_31_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_111 ? _slots_34_io_out_uop_prs1 : _GEN_110 ? _slots_33_io_out_uop_prs1 : _GEN_109 ? _slots_32_io_out_uop_prs1 : _slots_31_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_111 ? _slots_34_io_out_uop_prs2 : _GEN_110 ? _slots_33_io_out_uop_prs2 : _GEN_109 ? _slots_32_io_out_uop_prs2 : _slots_31_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_111 ? _slots_34_io_out_uop_prs3 : _GEN_110 ? _slots_33_io_out_uop_prs3 : _GEN_109 ? _slots_32_io_out_uop_prs3 : _slots_31_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_111 ? _slots_34_io_out_uop_ppred : _GEN_110 ? _slots_33_io_out_uop_ppred : _GEN_109 ? _slots_32_io_out_uop_ppred : _slots_31_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_111 ? _slots_34_io_out_uop_prs1_busy : _GEN_110 ? _slots_33_io_out_uop_prs1_busy : _GEN_109 ? _slots_32_io_out_uop_prs1_busy : _slots_31_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_111 ? _slots_34_io_out_uop_prs2_busy : _GEN_110 ? _slots_33_io_out_uop_prs2_busy : _GEN_109 ? _slots_32_io_out_uop_prs2_busy : _slots_31_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_111 ? _slots_34_io_out_uop_prs3_busy : _GEN_110 ? _slots_33_io_out_uop_prs3_busy : _GEN_109 ? _slots_32_io_out_uop_prs3_busy : _slots_31_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_111 ? _slots_34_io_out_uop_ppred_busy : _GEN_110 ? _slots_33_io_out_uop_ppred_busy : _GEN_109 ? _slots_32_io_out_uop_ppred_busy : _slots_31_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_111 ? _slots_34_io_out_uop_stale_pdst : _GEN_110 ? _slots_33_io_out_uop_stale_pdst : _GEN_109 ? _slots_32_io_out_uop_stale_pdst : _slots_31_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_111 ? _slots_34_io_out_uop_exception : _GEN_110 ? _slots_33_io_out_uop_exception : _GEN_109 ? _slots_32_io_out_uop_exception : _slots_31_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_111 ? _slots_34_io_out_uop_exc_cause : _GEN_110 ? _slots_33_io_out_uop_exc_cause : _GEN_109 ? _slots_32_io_out_uop_exc_cause : _slots_31_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_111 ? _slots_34_io_out_uop_bypassable : _GEN_110 ? _slots_33_io_out_uop_bypassable : _GEN_109 ? _slots_32_io_out_uop_bypassable : _slots_31_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_111 ? _slots_34_io_out_uop_mem_cmd : _GEN_110 ? _slots_33_io_out_uop_mem_cmd : _GEN_109 ? _slots_32_io_out_uop_mem_cmd : _slots_31_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_111 ? _slots_34_io_out_uop_mem_size : _GEN_110 ? _slots_33_io_out_uop_mem_size : _GEN_109 ? _slots_32_io_out_uop_mem_size : _slots_31_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_111 ? _slots_34_io_out_uop_mem_signed : _GEN_110 ? _slots_33_io_out_uop_mem_signed : _GEN_109 ? _slots_32_io_out_uop_mem_signed : _slots_31_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_111 ? _slots_34_io_out_uop_is_fence : _GEN_110 ? _slots_33_io_out_uop_is_fence : _GEN_109 ? _slots_32_io_out_uop_is_fence : _slots_31_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_111 ? _slots_34_io_out_uop_is_fencei : _GEN_110 ? _slots_33_io_out_uop_is_fencei : _GEN_109 ? _slots_32_io_out_uop_is_fencei : _slots_31_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_111 ? _slots_34_io_out_uop_is_amo : _GEN_110 ? _slots_33_io_out_uop_is_amo : _GEN_109 ? _slots_32_io_out_uop_is_amo : _slots_31_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_111 ? _slots_34_io_out_uop_uses_ldq : _GEN_110 ? _slots_33_io_out_uop_uses_ldq : _GEN_109 ? _slots_32_io_out_uop_uses_ldq : _slots_31_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_111 ? _slots_34_io_out_uop_uses_stq : _GEN_110 ? _slots_33_io_out_uop_uses_stq : _GEN_109 ? _slots_32_io_out_uop_uses_stq : _slots_31_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_111 ? _slots_34_io_out_uop_is_sys_pc2epc : _GEN_110 ? _slots_33_io_out_uop_is_sys_pc2epc : _GEN_109 ? _slots_32_io_out_uop_is_sys_pc2epc : _slots_31_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_111 ? _slots_34_io_out_uop_is_unique : _GEN_110 ? _slots_33_io_out_uop_is_unique : _GEN_109 ? _slots_32_io_out_uop_is_unique : _slots_31_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_111 ? _slots_34_io_out_uop_flush_on_commit : _GEN_110 ? _slots_33_io_out_uop_flush_on_commit : _GEN_109 ? _slots_32_io_out_uop_flush_on_commit : _slots_31_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_111 ? _slots_34_io_out_uop_ldst_is_rs1 : _GEN_110 ? _slots_33_io_out_uop_ldst_is_rs1 : _GEN_109 ? _slots_32_io_out_uop_ldst_is_rs1 : _slots_31_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_111 ? _slots_34_io_out_uop_ldst : _GEN_110 ? _slots_33_io_out_uop_ldst : _GEN_109 ? _slots_32_io_out_uop_ldst : _slots_31_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_111 ? _slots_34_io_out_uop_lrs1 : _GEN_110 ? _slots_33_io_out_uop_lrs1 : _GEN_109 ? _slots_32_io_out_uop_lrs1 : _slots_31_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_111 ? _slots_34_io_out_uop_lrs2 : _GEN_110 ? _slots_33_io_out_uop_lrs2 : _GEN_109 ? _slots_32_io_out_uop_lrs2 : _slots_31_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_111 ? _slots_34_io_out_uop_lrs3 : _GEN_110 ? _slots_33_io_out_uop_lrs3 : _GEN_109 ? _slots_32_io_out_uop_lrs3 : _slots_31_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_111 ? _slots_34_io_out_uop_ldst_val : _GEN_110 ? _slots_33_io_out_uop_ldst_val : _GEN_109 ? _slots_32_io_out_uop_ldst_val : _slots_31_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_111 ? _slots_34_io_out_uop_dst_rtype : _GEN_110 ? _slots_33_io_out_uop_dst_rtype : _GEN_109 ? _slots_32_io_out_uop_dst_rtype : _slots_31_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_111 ? _slots_34_io_out_uop_lrs1_rtype : _GEN_110 ? _slots_33_io_out_uop_lrs1_rtype : _GEN_109 ? _slots_32_io_out_uop_lrs1_rtype : _slots_31_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_111 ? _slots_34_io_out_uop_lrs2_rtype : _GEN_110 ? _slots_33_io_out_uop_lrs2_rtype : _GEN_109 ? _slots_32_io_out_uop_lrs2_rtype : _slots_31_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_111 ? _slots_34_io_out_uop_frs3_en : _GEN_110 ? _slots_33_io_out_uop_frs3_en : _GEN_109 ? _slots_32_io_out_uop_frs3_en : _slots_31_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_111 ? _slots_34_io_out_uop_fp_val : _GEN_110 ? _slots_33_io_out_uop_fp_val : _GEN_109 ? _slots_32_io_out_uop_fp_val : _slots_31_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_111 ? _slots_34_io_out_uop_fp_single : _GEN_110 ? _slots_33_io_out_uop_fp_single : _GEN_109 ? _slots_32_io_out_uop_fp_single : _slots_31_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_111 ? _slots_34_io_out_uop_xcpt_pf_if : _GEN_110 ? _slots_33_io_out_uop_xcpt_pf_if : _GEN_109 ? _slots_32_io_out_uop_xcpt_pf_if : _slots_31_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_111 ? _slots_34_io_out_uop_xcpt_ae_if : _GEN_110 ? _slots_33_io_out_uop_xcpt_ae_if : _GEN_109 ? _slots_32_io_out_uop_xcpt_ae_if : _slots_31_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_111 ? _slots_34_io_out_uop_xcpt_ma_if : _GEN_110 ? _slots_33_io_out_uop_xcpt_ma_if : _GEN_109 ? _slots_32_io_out_uop_xcpt_ma_if : _slots_31_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_111 ? _slots_34_io_out_uop_bp_debug_if : _GEN_110 ? _slots_33_io_out_uop_bp_debug_if : _GEN_109 ? _slots_32_io_out_uop_bp_debug_if : _slots_31_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_111 ? _slots_34_io_out_uop_bp_xcpt_if : _GEN_110 ? _slots_33_io_out_uop_bp_xcpt_if : _GEN_109 ? _slots_32_io_out_uop_bp_xcpt_if : _slots_31_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_111 ? _slots_34_io_out_uop_debug_fsrc : _GEN_110 ? _slots_33_io_out_uop_debug_fsrc : _GEN_109 ? _slots_32_io_out_uop_debug_fsrc : _slots_31_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_111 ? _slots_34_io_out_uop_debug_tsrc : _GEN_110 ? _slots_33_io_out_uop_debug_tsrc : _GEN_109 ? _slots_32_io_out_uop_debug_tsrc : _slots_31_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_30_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_30_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_30_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_30_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_30_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_30_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_30_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_30_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_30_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_30_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_30_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_30_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_30_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_30_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_30_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_30_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_30_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_30_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_30_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_30_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_30_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_30_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_30_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_30_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_30_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_30_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_30_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_30_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_30_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_30_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_30_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_30_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_30_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_30_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_30_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_30_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_30_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_30_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_30_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_30_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_30_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_30_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_30_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_30_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_30_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_30_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_30_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_30_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_30_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_30_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_30_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_30_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_30_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_30_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_30_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_30_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_30_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_30_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_30_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_30_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_30_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_30_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_30_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_30_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_30_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_30_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_30_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_30_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_30_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_30_io_uop_uopc),
    .io_uop_inst                    (_slots_30_io_uop_inst),
    .io_uop_debug_inst              (_slots_30_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_30_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_30_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_30_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_30_io_uop_fu_code),
    .io_uop_iw_state                (_slots_30_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_30_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_30_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_30_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_30_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_30_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_30_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_30_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_30_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_30_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_30_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_30_io_uop_pc_lob),
    .io_uop_taken                   (_slots_30_io_uop_taken),
    .io_uop_imm_packed              (_slots_30_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_30_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_30_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_30_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_30_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_30_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_30_io_uop_pdst),
    .io_uop_prs1                    (_slots_30_io_uop_prs1),
    .io_uop_prs2                    (_slots_30_io_uop_prs2),
    .io_uop_prs3                    (_slots_30_io_uop_prs3),
    .io_uop_ppred                   (_slots_30_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_30_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_30_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_30_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_30_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_30_io_uop_stale_pdst),
    .io_uop_exception               (_slots_30_io_uop_exception),
    .io_uop_exc_cause               (_slots_30_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_30_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_30_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_30_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_30_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_30_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_30_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_30_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_30_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_30_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_30_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_30_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_30_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_30_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_30_io_uop_ldst),
    .io_uop_lrs1                    (_slots_30_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_30_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_30_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_30_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_30_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_30_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_30_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_30_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_30_io_uop_fp_val),
    .io_uop_fp_single               (_slots_30_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_30_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_30_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_30_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_30_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_30_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_30_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_30_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_31 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_31_io_valid),
    .io_will_be_valid               (_slots_31_io_will_be_valid),
    .io_request                     (_slots_31_io_request),
    .io_grant                       (issue_slots_31_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_30),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_31_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_114 ? _slots_35_io_out_uop_uopc : _GEN_113 ? _slots_34_io_out_uop_uopc : _GEN_112 ? _slots_33_io_out_uop_uopc : _slots_32_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_114 ? _slots_35_io_out_uop_inst : _GEN_113 ? _slots_34_io_out_uop_inst : _GEN_112 ? _slots_33_io_out_uop_inst : _slots_32_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_114 ? _slots_35_io_out_uop_debug_inst : _GEN_113 ? _slots_34_io_out_uop_debug_inst : _GEN_112 ? _slots_33_io_out_uop_debug_inst : _slots_32_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_114 ? _slots_35_io_out_uop_is_rvc : _GEN_113 ? _slots_34_io_out_uop_is_rvc : _GEN_112 ? _slots_33_io_out_uop_is_rvc : _slots_32_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_114 ? _slots_35_io_out_uop_debug_pc : _GEN_113 ? _slots_34_io_out_uop_debug_pc : _GEN_112 ? _slots_33_io_out_uop_debug_pc : _slots_32_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_114 ? _slots_35_io_out_uop_iq_type : _GEN_113 ? _slots_34_io_out_uop_iq_type : _GEN_112 ? _slots_33_io_out_uop_iq_type : _slots_32_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_114 ? _slots_35_io_out_uop_fu_code : _GEN_113 ? _slots_34_io_out_uop_fu_code : _GEN_112 ? _slots_33_io_out_uop_fu_code : _slots_32_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_114 ? _slots_35_io_out_uop_iw_state : _GEN_113 ? _slots_34_io_out_uop_iw_state : _GEN_112 ? _slots_33_io_out_uop_iw_state : _slots_32_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_114 ? _slots_35_io_out_uop_iw_p1_poisoned : _GEN_113 ? _slots_34_io_out_uop_iw_p1_poisoned : _GEN_112 ? _slots_33_io_out_uop_iw_p1_poisoned : _slots_32_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_114 ? _slots_35_io_out_uop_iw_p2_poisoned : _GEN_113 ? _slots_34_io_out_uop_iw_p2_poisoned : _GEN_112 ? _slots_33_io_out_uop_iw_p2_poisoned : _slots_32_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_114 ? _slots_35_io_out_uop_is_br : _GEN_113 ? _slots_34_io_out_uop_is_br : _GEN_112 ? _slots_33_io_out_uop_is_br : _slots_32_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_114 ? _slots_35_io_out_uop_is_jalr : _GEN_113 ? _slots_34_io_out_uop_is_jalr : _GEN_112 ? _slots_33_io_out_uop_is_jalr : _slots_32_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_114 ? _slots_35_io_out_uop_is_jal : _GEN_113 ? _slots_34_io_out_uop_is_jal : _GEN_112 ? _slots_33_io_out_uop_is_jal : _slots_32_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_114 ? _slots_35_io_out_uop_is_sfb : _GEN_113 ? _slots_34_io_out_uop_is_sfb : _GEN_112 ? _slots_33_io_out_uop_is_sfb : _slots_32_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_114 ? _slots_35_io_out_uop_br_mask : _GEN_113 ? _slots_34_io_out_uop_br_mask : _GEN_112 ? _slots_33_io_out_uop_br_mask : _slots_32_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_114 ? _slots_35_io_out_uop_br_tag : _GEN_113 ? _slots_34_io_out_uop_br_tag : _GEN_112 ? _slots_33_io_out_uop_br_tag : _slots_32_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_114 ? _slots_35_io_out_uop_ftq_idx : _GEN_113 ? _slots_34_io_out_uop_ftq_idx : _GEN_112 ? _slots_33_io_out_uop_ftq_idx : _slots_32_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_114 ? _slots_35_io_out_uop_edge_inst : _GEN_113 ? _slots_34_io_out_uop_edge_inst : _GEN_112 ? _slots_33_io_out_uop_edge_inst : _slots_32_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_114 ? _slots_35_io_out_uop_pc_lob : _GEN_113 ? _slots_34_io_out_uop_pc_lob : _GEN_112 ? _slots_33_io_out_uop_pc_lob : _slots_32_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_114 ? _slots_35_io_out_uop_taken : _GEN_113 ? _slots_34_io_out_uop_taken : _GEN_112 ? _slots_33_io_out_uop_taken : _slots_32_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_114 ? _slots_35_io_out_uop_imm_packed : _GEN_113 ? _slots_34_io_out_uop_imm_packed : _GEN_112 ? _slots_33_io_out_uop_imm_packed : _slots_32_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_114 ? _slots_35_io_out_uop_csr_addr : _GEN_113 ? _slots_34_io_out_uop_csr_addr : _GEN_112 ? _slots_33_io_out_uop_csr_addr : _slots_32_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_114 ? _slots_35_io_out_uop_rob_idx : _GEN_113 ? _slots_34_io_out_uop_rob_idx : _GEN_112 ? _slots_33_io_out_uop_rob_idx : _slots_32_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_114 ? _slots_35_io_out_uop_ldq_idx : _GEN_113 ? _slots_34_io_out_uop_ldq_idx : _GEN_112 ? _slots_33_io_out_uop_ldq_idx : _slots_32_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_114 ? _slots_35_io_out_uop_stq_idx : _GEN_113 ? _slots_34_io_out_uop_stq_idx : _GEN_112 ? _slots_33_io_out_uop_stq_idx : _slots_32_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_114 ? _slots_35_io_out_uop_rxq_idx : _GEN_113 ? _slots_34_io_out_uop_rxq_idx : _GEN_112 ? _slots_33_io_out_uop_rxq_idx : _slots_32_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_114 ? _slots_35_io_out_uop_pdst : _GEN_113 ? _slots_34_io_out_uop_pdst : _GEN_112 ? _slots_33_io_out_uop_pdst : _slots_32_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_114 ? _slots_35_io_out_uop_prs1 : _GEN_113 ? _slots_34_io_out_uop_prs1 : _GEN_112 ? _slots_33_io_out_uop_prs1 : _slots_32_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_114 ? _slots_35_io_out_uop_prs2 : _GEN_113 ? _slots_34_io_out_uop_prs2 : _GEN_112 ? _slots_33_io_out_uop_prs2 : _slots_32_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_114 ? _slots_35_io_out_uop_prs3 : _GEN_113 ? _slots_34_io_out_uop_prs3 : _GEN_112 ? _slots_33_io_out_uop_prs3 : _slots_32_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_114 ? _slots_35_io_out_uop_ppred : _GEN_113 ? _slots_34_io_out_uop_ppred : _GEN_112 ? _slots_33_io_out_uop_ppred : _slots_32_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_114 ? _slots_35_io_out_uop_prs1_busy : _GEN_113 ? _slots_34_io_out_uop_prs1_busy : _GEN_112 ? _slots_33_io_out_uop_prs1_busy : _slots_32_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_114 ? _slots_35_io_out_uop_prs2_busy : _GEN_113 ? _slots_34_io_out_uop_prs2_busy : _GEN_112 ? _slots_33_io_out_uop_prs2_busy : _slots_32_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_114 ? _slots_35_io_out_uop_prs3_busy : _GEN_113 ? _slots_34_io_out_uop_prs3_busy : _GEN_112 ? _slots_33_io_out_uop_prs3_busy : _slots_32_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_114 ? _slots_35_io_out_uop_ppred_busy : _GEN_113 ? _slots_34_io_out_uop_ppred_busy : _GEN_112 ? _slots_33_io_out_uop_ppred_busy : _slots_32_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_114 ? _slots_35_io_out_uop_stale_pdst : _GEN_113 ? _slots_34_io_out_uop_stale_pdst : _GEN_112 ? _slots_33_io_out_uop_stale_pdst : _slots_32_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_114 ? _slots_35_io_out_uop_exception : _GEN_113 ? _slots_34_io_out_uop_exception : _GEN_112 ? _slots_33_io_out_uop_exception : _slots_32_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_114 ? _slots_35_io_out_uop_exc_cause : _GEN_113 ? _slots_34_io_out_uop_exc_cause : _GEN_112 ? _slots_33_io_out_uop_exc_cause : _slots_32_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_114 ? _slots_35_io_out_uop_bypassable : _GEN_113 ? _slots_34_io_out_uop_bypassable : _GEN_112 ? _slots_33_io_out_uop_bypassable : _slots_32_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_114 ? _slots_35_io_out_uop_mem_cmd : _GEN_113 ? _slots_34_io_out_uop_mem_cmd : _GEN_112 ? _slots_33_io_out_uop_mem_cmd : _slots_32_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_114 ? _slots_35_io_out_uop_mem_size : _GEN_113 ? _slots_34_io_out_uop_mem_size : _GEN_112 ? _slots_33_io_out_uop_mem_size : _slots_32_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_114 ? _slots_35_io_out_uop_mem_signed : _GEN_113 ? _slots_34_io_out_uop_mem_signed : _GEN_112 ? _slots_33_io_out_uop_mem_signed : _slots_32_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_114 ? _slots_35_io_out_uop_is_fence : _GEN_113 ? _slots_34_io_out_uop_is_fence : _GEN_112 ? _slots_33_io_out_uop_is_fence : _slots_32_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_114 ? _slots_35_io_out_uop_is_fencei : _GEN_113 ? _slots_34_io_out_uop_is_fencei : _GEN_112 ? _slots_33_io_out_uop_is_fencei : _slots_32_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_114 ? _slots_35_io_out_uop_is_amo : _GEN_113 ? _slots_34_io_out_uop_is_amo : _GEN_112 ? _slots_33_io_out_uop_is_amo : _slots_32_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_114 ? _slots_35_io_out_uop_uses_ldq : _GEN_113 ? _slots_34_io_out_uop_uses_ldq : _GEN_112 ? _slots_33_io_out_uop_uses_ldq : _slots_32_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_114 ? _slots_35_io_out_uop_uses_stq : _GEN_113 ? _slots_34_io_out_uop_uses_stq : _GEN_112 ? _slots_33_io_out_uop_uses_stq : _slots_32_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_114 ? _slots_35_io_out_uop_is_sys_pc2epc : _GEN_113 ? _slots_34_io_out_uop_is_sys_pc2epc : _GEN_112 ? _slots_33_io_out_uop_is_sys_pc2epc : _slots_32_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_114 ? _slots_35_io_out_uop_is_unique : _GEN_113 ? _slots_34_io_out_uop_is_unique : _GEN_112 ? _slots_33_io_out_uop_is_unique : _slots_32_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_114 ? _slots_35_io_out_uop_flush_on_commit : _GEN_113 ? _slots_34_io_out_uop_flush_on_commit : _GEN_112 ? _slots_33_io_out_uop_flush_on_commit : _slots_32_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_114 ? _slots_35_io_out_uop_ldst_is_rs1 : _GEN_113 ? _slots_34_io_out_uop_ldst_is_rs1 : _GEN_112 ? _slots_33_io_out_uop_ldst_is_rs1 : _slots_32_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_114 ? _slots_35_io_out_uop_ldst : _GEN_113 ? _slots_34_io_out_uop_ldst : _GEN_112 ? _slots_33_io_out_uop_ldst : _slots_32_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_114 ? _slots_35_io_out_uop_lrs1 : _GEN_113 ? _slots_34_io_out_uop_lrs1 : _GEN_112 ? _slots_33_io_out_uop_lrs1 : _slots_32_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_114 ? _slots_35_io_out_uop_lrs2 : _GEN_113 ? _slots_34_io_out_uop_lrs2 : _GEN_112 ? _slots_33_io_out_uop_lrs2 : _slots_32_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_114 ? _slots_35_io_out_uop_lrs3 : _GEN_113 ? _slots_34_io_out_uop_lrs3 : _GEN_112 ? _slots_33_io_out_uop_lrs3 : _slots_32_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_114 ? _slots_35_io_out_uop_ldst_val : _GEN_113 ? _slots_34_io_out_uop_ldst_val : _GEN_112 ? _slots_33_io_out_uop_ldst_val : _slots_32_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_114 ? _slots_35_io_out_uop_dst_rtype : _GEN_113 ? _slots_34_io_out_uop_dst_rtype : _GEN_112 ? _slots_33_io_out_uop_dst_rtype : _slots_32_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_114 ? _slots_35_io_out_uop_lrs1_rtype : _GEN_113 ? _slots_34_io_out_uop_lrs1_rtype : _GEN_112 ? _slots_33_io_out_uop_lrs1_rtype : _slots_32_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_114 ? _slots_35_io_out_uop_lrs2_rtype : _GEN_113 ? _slots_34_io_out_uop_lrs2_rtype : _GEN_112 ? _slots_33_io_out_uop_lrs2_rtype : _slots_32_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_114 ? _slots_35_io_out_uop_frs3_en : _GEN_113 ? _slots_34_io_out_uop_frs3_en : _GEN_112 ? _slots_33_io_out_uop_frs3_en : _slots_32_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_114 ? _slots_35_io_out_uop_fp_val : _GEN_113 ? _slots_34_io_out_uop_fp_val : _GEN_112 ? _slots_33_io_out_uop_fp_val : _slots_32_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_114 ? _slots_35_io_out_uop_fp_single : _GEN_113 ? _slots_34_io_out_uop_fp_single : _GEN_112 ? _slots_33_io_out_uop_fp_single : _slots_32_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_114 ? _slots_35_io_out_uop_xcpt_pf_if : _GEN_113 ? _slots_34_io_out_uop_xcpt_pf_if : _GEN_112 ? _slots_33_io_out_uop_xcpt_pf_if : _slots_32_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_114 ? _slots_35_io_out_uop_xcpt_ae_if : _GEN_113 ? _slots_34_io_out_uop_xcpt_ae_if : _GEN_112 ? _slots_33_io_out_uop_xcpt_ae_if : _slots_32_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_114 ? _slots_35_io_out_uop_xcpt_ma_if : _GEN_113 ? _slots_34_io_out_uop_xcpt_ma_if : _GEN_112 ? _slots_33_io_out_uop_xcpt_ma_if : _slots_32_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_114 ? _slots_35_io_out_uop_bp_debug_if : _GEN_113 ? _slots_34_io_out_uop_bp_debug_if : _GEN_112 ? _slots_33_io_out_uop_bp_debug_if : _slots_32_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_114 ? _slots_35_io_out_uop_bp_xcpt_if : _GEN_113 ? _slots_34_io_out_uop_bp_xcpt_if : _GEN_112 ? _slots_33_io_out_uop_bp_xcpt_if : _slots_32_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_114 ? _slots_35_io_out_uop_debug_fsrc : _GEN_113 ? _slots_34_io_out_uop_debug_fsrc : _GEN_112 ? _slots_33_io_out_uop_debug_fsrc : _slots_32_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_114 ? _slots_35_io_out_uop_debug_tsrc : _GEN_113 ? _slots_34_io_out_uop_debug_tsrc : _GEN_112 ? _slots_33_io_out_uop_debug_tsrc : _slots_32_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_31_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_31_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_31_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_31_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_31_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_31_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_31_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_31_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_31_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_31_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_31_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_31_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_31_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_31_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_31_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_31_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_31_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_31_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_31_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_31_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_31_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_31_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_31_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_31_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_31_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_31_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_31_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_31_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_31_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_31_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_31_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_31_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_31_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_31_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_31_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_31_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_31_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_31_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_31_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_31_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_31_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_31_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_31_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_31_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_31_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_31_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_31_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_31_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_31_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_31_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_31_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_31_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_31_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_31_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_31_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_31_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_31_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_31_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_31_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_31_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_31_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_31_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_31_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_31_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_31_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_31_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_31_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_31_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_31_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_31_io_uop_uopc),
    .io_uop_inst                    (_slots_31_io_uop_inst),
    .io_uop_debug_inst              (_slots_31_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_31_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_31_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_31_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_31_io_uop_fu_code),
    .io_uop_iw_state                (_slots_31_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_31_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_31_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_31_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_31_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_31_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_31_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_31_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_31_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_31_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_31_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_31_io_uop_pc_lob),
    .io_uop_taken                   (_slots_31_io_uop_taken),
    .io_uop_imm_packed              (_slots_31_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_31_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_31_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_31_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_31_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_31_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_31_io_uop_pdst),
    .io_uop_prs1                    (_slots_31_io_uop_prs1),
    .io_uop_prs2                    (_slots_31_io_uop_prs2),
    .io_uop_prs3                    (_slots_31_io_uop_prs3),
    .io_uop_ppred                   (_slots_31_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_31_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_31_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_31_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_31_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_31_io_uop_stale_pdst),
    .io_uop_exception               (_slots_31_io_uop_exception),
    .io_uop_exc_cause               (_slots_31_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_31_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_31_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_31_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_31_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_31_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_31_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_31_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_31_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_31_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_31_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_31_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_31_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_31_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_31_io_uop_ldst),
    .io_uop_lrs1                    (_slots_31_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_31_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_31_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_31_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_31_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_31_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_31_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_31_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_31_io_uop_fp_val),
    .io_uop_fp_single               (_slots_31_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_31_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_31_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_31_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_31_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_31_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_31_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_31_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_32 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_32_io_valid),
    .io_will_be_valid               (_slots_32_io_will_be_valid),
    .io_request                     (_slots_32_io_request),
    .io_grant                       (issue_slots_32_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_31),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_32_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_117 ? _slots_36_io_out_uop_uopc : _GEN_116 ? _slots_35_io_out_uop_uopc : _GEN_115 ? _slots_34_io_out_uop_uopc : _slots_33_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_117 ? _slots_36_io_out_uop_inst : _GEN_116 ? _slots_35_io_out_uop_inst : _GEN_115 ? _slots_34_io_out_uop_inst : _slots_33_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_117 ? _slots_36_io_out_uop_debug_inst : _GEN_116 ? _slots_35_io_out_uop_debug_inst : _GEN_115 ? _slots_34_io_out_uop_debug_inst : _slots_33_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_117 ? _slots_36_io_out_uop_is_rvc : _GEN_116 ? _slots_35_io_out_uop_is_rvc : _GEN_115 ? _slots_34_io_out_uop_is_rvc : _slots_33_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_117 ? _slots_36_io_out_uop_debug_pc : _GEN_116 ? _slots_35_io_out_uop_debug_pc : _GEN_115 ? _slots_34_io_out_uop_debug_pc : _slots_33_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_117 ? _slots_36_io_out_uop_iq_type : _GEN_116 ? _slots_35_io_out_uop_iq_type : _GEN_115 ? _slots_34_io_out_uop_iq_type : _slots_33_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_117 ? _slots_36_io_out_uop_fu_code : _GEN_116 ? _slots_35_io_out_uop_fu_code : _GEN_115 ? _slots_34_io_out_uop_fu_code : _slots_33_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_117 ? _slots_36_io_out_uop_iw_state : _GEN_116 ? _slots_35_io_out_uop_iw_state : _GEN_115 ? _slots_34_io_out_uop_iw_state : _slots_33_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_117 ? _slots_36_io_out_uop_iw_p1_poisoned : _GEN_116 ? _slots_35_io_out_uop_iw_p1_poisoned : _GEN_115 ? _slots_34_io_out_uop_iw_p1_poisoned : _slots_33_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_117 ? _slots_36_io_out_uop_iw_p2_poisoned : _GEN_116 ? _slots_35_io_out_uop_iw_p2_poisoned : _GEN_115 ? _slots_34_io_out_uop_iw_p2_poisoned : _slots_33_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_117 ? _slots_36_io_out_uop_is_br : _GEN_116 ? _slots_35_io_out_uop_is_br : _GEN_115 ? _slots_34_io_out_uop_is_br : _slots_33_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_117 ? _slots_36_io_out_uop_is_jalr : _GEN_116 ? _slots_35_io_out_uop_is_jalr : _GEN_115 ? _slots_34_io_out_uop_is_jalr : _slots_33_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_117 ? _slots_36_io_out_uop_is_jal : _GEN_116 ? _slots_35_io_out_uop_is_jal : _GEN_115 ? _slots_34_io_out_uop_is_jal : _slots_33_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_117 ? _slots_36_io_out_uop_is_sfb : _GEN_116 ? _slots_35_io_out_uop_is_sfb : _GEN_115 ? _slots_34_io_out_uop_is_sfb : _slots_33_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_117 ? _slots_36_io_out_uop_br_mask : _GEN_116 ? _slots_35_io_out_uop_br_mask : _GEN_115 ? _slots_34_io_out_uop_br_mask : _slots_33_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_117 ? _slots_36_io_out_uop_br_tag : _GEN_116 ? _slots_35_io_out_uop_br_tag : _GEN_115 ? _slots_34_io_out_uop_br_tag : _slots_33_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_117 ? _slots_36_io_out_uop_ftq_idx : _GEN_116 ? _slots_35_io_out_uop_ftq_idx : _GEN_115 ? _slots_34_io_out_uop_ftq_idx : _slots_33_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_117 ? _slots_36_io_out_uop_edge_inst : _GEN_116 ? _slots_35_io_out_uop_edge_inst : _GEN_115 ? _slots_34_io_out_uop_edge_inst : _slots_33_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_117 ? _slots_36_io_out_uop_pc_lob : _GEN_116 ? _slots_35_io_out_uop_pc_lob : _GEN_115 ? _slots_34_io_out_uop_pc_lob : _slots_33_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_117 ? _slots_36_io_out_uop_taken : _GEN_116 ? _slots_35_io_out_uop_taken : _GEN_115 ? _slots_34_io_out_uop_taken : _slots_33_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_117 ? _slots_36_io_out_uop_imm_packed : _GEN_116 ? _slots_35_io_out_uop_imm_packed : _GEN_115 ? _slots_34_io_out_uop_imm_packed : _slots_33_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_117 ? _slots_36_io_out_uop_csr_addr : _GEN_116 ? _slots_35_io_out_uop_csr_addr : _GEN_115 ? _slots_34_io_out_uop_csr_addr : _slots_33_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_117 ? _slots_36_io_out_uop_rob_idx : _GEN_116 ? _slots_35_io_out_uop_rob_idx : _GEN_115 ? _slots_34_io_out_uop_rob_idx : _slots_33_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_117 ? _slots_36_io_out_uop_ldq_idx : _GEN_116 ? _slots_35_io_out_uop_ldq_idx : _GEN_115 ? _slots_34_io_out_uop_ldq_idx : _slots_33_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_117 ? _slots_36_io_out_uop_stq_idx : _GEN_116 ? _slots_35_io_out_uop_stq_idx : _GEN_115 ? _slots_34_io_out_uop_stq_idx : _slots_33_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_117 ? _slots_36_io_out_uop_rxq_idx : _GEN_116 ? _slots_35_io_out_uop_rxq_idx : _GEN_115 ? _slots_34_io_out_uop_rxq_idx : _slots_33_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_117 ? _slots_36_io_out_uop_pdst : _GEN_116 ? _slots_35_io_out_uop_pdst : _GEN_115 ? _slots_34_io_out_uop_pdst : _slots_33_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_117 ? _slots_36_io_out_uop_prs1 : _GEN_116 ? _slots_35_io_out_uop_prs1 : _GEN_115 ? _slots_34_io_out_uop_prs1 : _slots_33_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_117 ? _slots_36_io_out_uop_prs2 : _GEN_116 ? _slots_35_io_out_uop_prs2 : _GEN_115 ? _slots_34_io_out_uop_prs2 : _slots_33_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_117 ? _slots_36_io_out_uop_prs3 : _GEN_116 ? _slots_35_io_out_uop_prs3 : _GEN_115 ? _slots_34_io_out_uop_prs3 : _slots_33_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_117 ? _slots_36_io_out_uop_ppred : _GEN_116 ? _slots_35_io_out_uop_ppred : _GEN_115 ? _slots_34_io_out_uop_ppred : _slots_33_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_117 ? _slots_36_io_out_uop_prs1_busy : _GEN_116 ? _slots_35_io_out_uop_prs1_busy : _GEN_115 ? _slots_34_io_out_uop_prs1_busy : _slots_33_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_117 ? _slots_36_io_out_uop_prs2_busy : _GEN_116 ? _slots_35_io_out_uop_prs2_busy : _GEN_115 ? _slots_34_io_out_uop_prs2_busy : _slots_33_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_117 ? _slots_36_io_out_uop_prs3_busy : _GEN_116 ? _slots_35_io_out_uop_prs3_busy : _GEN_115 ? _slots_34_io_out_uop_prs3_busy : _slots_33_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_117 ? _slots_36_io_out_uop_ppred_busy : _GEN_116 ? _slots_35_io_out_uop_ppred_busy : _GEN_115 ? _slots_34_io_out_uop_ppred_busy : _slots_33_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_117 ? _slots_36_io_out_uop_stale_pdst : _GEN_116 ? _slots_35_io_out_uop_stale_pdst : _GEN_115 ? _slots_34_io_out_uop_stale_pdst : _slots_33_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_117 ? _slots_36_io_out_uop_exception : _GEN_116 ? _slots_35_io_out_uop_exception : _GEN_115 ? _slots_34_io_out_uop_exception : _slots_33_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_117 ? _slots_36_io_out_uop_exc_cause : _GEN_116 ? _slots_35_io_out_uop_exc_cause : _GEN_115 ? _slots_34_io_out_uop_exc_cause : _slots_33_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_117 ? _slots_36_io_out_uop_bypassable : _GEN_116 ? _slots_35_io_out_uop_bypassable : _GEN_115 ? _slots_34_io_out_uop_bypassable : _slots_33_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_117 ? _slots_36_io_out_uop_mem_cmd : _GEN_116 ? _slots_35_io_out_uop_mem_cmd : _GEN_115 ? _slots_34_io_out_uop_mem_cmd : _slots_33_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_117 ? _slots_36_io_out_uop_mem_size : _GEN_116 ? _slots_35_io_out_uop_mem_size : _GEN_115 ? _slots_34_io_out_uop_mem_size : _slots_33_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_117 ? _slots_36_io_out_uop_mem_signed : _GEN_116 ? _slots_35_io_out_uop_mem_signed : _GEN_115 ? _slots_34_io_out_uop_mem_signed : _slots_33_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_117 ? _slots_36_io_out_uop_is_fence : _GEN_116 ? _slots_35_io_out_uop_is_fence : _GEN_115 ? _slots_34_io_out_uop_is_fence : _slots_33_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_117 ? _slots_36_io_out_uop_is_fencei : _GEN_116 ? _slots_35_io_out_uop_is_fencei : _GEN_115 ? _slots_34_io_out_uop_is_fencei : _slots_33_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_117 ? _slots_36_io_out_uop_is_amo : _GEN_116 ? _slots_35_io_out_uop_is_amo : _GEN_115 ? _slots_34_io_out_uop_is_amo : _slots_33_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_117 ? _slots_36_io_out_uop_uses_ldq : _GEN_116 ? _slots_35_io_out_uop_uses_ldq : _GEN_115 ? _slots_34_io_out_uop_uses_ldq : _slots_33_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_117 ? _slots_36_io_out_uop_uses_stq : _GEN_116 ? _slots_35_io_out_uop_uses_stq : _GEN_115 ? _slots_34_io_out_uop_uses_stq : _slots_33_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_117 ? _slots_36_io_out_uop_is_sys_pc2epc : _GEN_116 ? _slots_35_io_out_uop_is_sys_pc2epc : _GEN_115 ? _slots_34_io_out_uop_is_sys_pc2epc : _slots_33_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_117 ? _slots_36_io_out_uop_is_unique : _GEN_116 ? _slots_35_io_out_uop_is_unique : _GEN_115 ? _slots_34_io_out_uop_is_unique : _slots_33_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_117 ? _slots_36_io_out_uop_flush_on_commit : _GEN_116 ? _slots_35_io_out_uop_flush_on_commit : _GEN_115 ? _slots_34_io_out_uop_flush_on_commit : _slots_33_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_117 ? _slots_36_io_out_uop_ldst_is_rs1 : _GEN_116 ? _slots_35_io_out_uop_ldst_is_rs1 : _GEN_115 ? _slots_34_io_out_uop_ldst_is_rs1 : _slots_33_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_117 ? _slots_36_io_out_uop_ldst : _GEN_116 ? _slots_35_io_out_uop_ldst : _GEN_115 ? _slots_34_io_out_uop_ldst : _slots_33_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_117 ? _slots_36_io_out_uop_lrs1 : _GEN_116 ? _slots_35_io_out_uop_lrs1 : _GEN_115 ? _slots_34_io_out_uop_lrs1 : _slots_33_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_117 ? _slots_36_io_out_uop_lrs2 : _GEN_116 ? _slots_35_io_out_uop_lrs2 : _GEN_115 ? _slots_34_io_out_uop_lrs2 : _slots_33_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_117 ? _slots_36_io_out_uop_lrs3 : _GEN_116 ? _slots_35_io_out_uop_lrs3 : _GEN_115 ? _slots_34_io_out_uop_lrs3 : _slots_33_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_117 ? _slots_36_io_out_uop_ldst_val : _GEN_116 ? _slots_35_io_out_uop_ldst_val : _GEN_115 ? _slots_34_io_out_uop_ldst_val : _slots_33_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_117 ? _slots_36_io_out_uop_dst_rtype : _GEN_116 ? _slots_35_io_out_uop_dst_rtype : _GEN_115 ? _slots_34_io_out_uop_dst_rtype : _slots_33_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_117 ? _slots_36_io_out_uop_lrs1_rtype : _GEN_116 ? _slots_35_io_out_uop_lrs1_rtype : _GEN_115 ? _slots_34_io_out_uop_lrs1_rtype : _slots_33_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_117 ? _slots_36_io_out_uop_lrs2_rtype : _GEN_116 ? _slots_35_io_out_uop_lrs2_rtype : _GEN_115 ? _slots_34_io_out_uop_lrs2_rtype : _slots_33_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_117 ? _slots_36_io_out_uop_frs3_en : _GEN_116 ? _slots_35_io_out_uop_frs3_en : _GEN_115 ? _slots_34_io_out_uop_frs3_en : _slots_33_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_117 ? _slots_36_io_out_uop_fp_val : _GEN_116 ? _slots_35_io_out_uop_fp_val : _GEN_115 ? _slots_34_io_out_uop_fp_val : _slots_33_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_117 ? _slots_36_io_out_uop_fp_single : _GEN_116 ? _slots_35_io_out_uop_fp_single : _GEN_115 ? _slots_34_io_out_uop_fp_single : _slots_33_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_117 ? _slots_36_io_out_uop_xcpt_pf_if : _GEN_116 ? _slots_35_io_out_uop_xcpt_pf_if : _GEN_115 ? _slots_34_io_out_uop_xcpt_pf_if : _slots_33_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_117 ? _slots_36_io_out_uop_xcpt_ae_if : _GEN_116 ? _slots_35_io_out_uop_xcpt_ae_if : _GEN_115 ? _slots_34_io_out_uop_xcpt_ae_if : _slots_33_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_117 ? _slots_36_io_out_uop_xcpt_ma_if : _GEN_116 ? _slots_35_io_out_uop_xcpt_ma_if : _GEN_115 ? _slots_34_io_out_uop_xcpt_ma_if : _slots_33_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_117 ? _slots_36_io_out_uop_bp_debug_if : _GEN_116 ? _slots_35_io_out_uop_bp_debug_if : _GEN_115 ? _slots_34_io_out_uop_bp_debug_if : _slots_33_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_117 ? _slots_36_io_out_uop_bp_xcpt_if : _GEN_116 ? _slots_35_io_out_uop_bp_xcpt_if : _GEN_115 ? _slots_34_io_out_uop_bp_xcpt_if : _slots_33_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_117 ? _slots_36_io_out_uop_debug_fsrc : _GEN_116 ? _slots_35_io_out_uop_debug_fsrc : _GEN_115 ? _slots_34_io_out_uop_debug_fsrc : _slots_33_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_117 ? _slots_36_io_out_uop_debug_tsrc : _GEN_116 ? _slots_35_io_out_uop_debug_tsrc : _GEN_115 ? _slots_34_io_out_uop_debug_tsrc : _slots_33_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_32_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_32_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_32_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_32_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_32_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_32_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_32_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_32_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_32_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_32_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_32_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_32_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_32_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_32_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_32_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_32_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_32_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_32_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_32_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_32_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_32_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_32_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_32_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_32_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_32_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_32_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_32_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_32_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_32_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_32_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_32_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_32_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_32_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_32_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_32_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_32_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_32_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_32_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_32_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_32_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_32_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_32_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_32_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_32_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_32_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_32_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_32_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_32_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_32_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_32_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_32_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_32_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_32_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_32_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_32_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_32_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_32_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_32_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_32_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_32_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_32_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_32_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_32_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_32_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_32_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_32_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_32_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_32_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_32_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_32_io_uop_uopc),
    .io_uop_inst                    (_slots_32_io_uop_inst),
    .io_uop_debug_inst              (_slots_32_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_32_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_32_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_32_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_32_io_uop_fu_code),
    .io_uop_iw_state                (_slots_32_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_32_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_32_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_32_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_32_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_32_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_32_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_32_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_32_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_32_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_32_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_32_io_uop_pc_lob),
    .io_uop_taken                   (_slots_32_io_uop_taken),
    .io_uop_imm_packed              (_slots_32_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_32_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_32_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_32_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_32_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_32_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_32_io_uop_pdst),
    .io_uop_prs1                    (_slots_32_io_uop_prs1),
    .io_uop_prs2                    (_slots_32_io_uop_prs2),
    .io_uop_prs3                    (_slots_32_io_uop_prs3),
    .io_uop_ppred                   (_slots_32_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_32_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_32_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_32_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_32_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_32_io_uop_stale_pdst),
    .io_uop_exception               (_slots_32_io_uop_exception),
    .io_uop_exc_cause               (_slots_32_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_32_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_32_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_32_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_32_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_32_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_32_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_32_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_32_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_32_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_32_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_32_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_32_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_32_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_32_io_uop_ldst),
    .io_uop_lrs1                    (_slots_32_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_32_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_32_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_32_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_32_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_32_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_32_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_32_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_32_io_uop_fp_val),
    .io_uop_fp_single               (_slots_32_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_32_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_32_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_32_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_32_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_32_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_32_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_32_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_33 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_33_io_valid),
    .io_will_be_valid               (_slots_33_io_will_be_valid),
    .io_request                     (_slots_33_io_request),
    .io_grant                       (issue_slots_33_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_32),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_33_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_120 ? _slots_37_io_out_uop_uopc : _GEN_119 ? _slots_36_io_out_uop_uopc : _GEN_118 ? _slots_35_io_out_uop_uopc : _slots_34_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_120 ? _slots_37_io_out_uop_inst : _GEN_119 ? _slots_36_io_out_uop_inst : _GEN_118 ? _slots_35_io_out_uop_inst : _slots_34_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_120 ? _slots_37_io_out_uop_debug_inst : _GEN_119 ? _slots_36_io_out_uop_debug_inst : _GEN_118 ? _slots_35_io_out_uop_debug_inst : _slots_34_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_120 ? _slots_37_io_out_uop_is_rvc : _GEN_119 ? _slots_36_io_out_uop_is_rvc : _GEN_118 ? _slots_35_io_out_uop_is_rvc : _slots_34_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_120 ? _slots_37_io_out_uop_debug_pc : _GEN_119 ? _slots_36_io_out_uop_debug_pc : _GEN_118 ? _slots_35_io_out_uop_debug_pc : _slots_34_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_120 ? _slots_37_io_out_uop_iq_type : _GEN_119 ? _slots_36_io_out_uop_iq_type : _GEN_118 ? _slots_35_io_out_uop_iq_type : _slots_34_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_120 ? _slots_37_io_out_uop_fu_code : _GEN_119 ? _slots_36_io_out_uop_fu_code : _GEN_118 ? _slots_35_io_out_uop_fu_code : _slots_34_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_120 ? _slots_37_io_out_uop_iw_state : _GEN_119 ? _slots_36_io_out_uop_iw_state : _GEN_118 ? _slots_35_io_out_uop_iw_state : _slots_34_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_120 ? _slots_37_io_out_uop_iw_p1_poisoned : _GEN_119 ? _slots_36_io_out_uop_iw_p1_poisoned : _GEN_118 ? _slots_35_io_out_uop_iw_p1_poisoned : _slots_34_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_120 ? _slots_37_io_out_uop_iw_p2_poisoned : _GEN_119 ? _slots_36_io_out_uop_iw_p2_poisoned : _GEN_118 ? _slots_35_io_out_uop_iw_p2_poisoned : _slots_34_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_120 ? _slots_37_io_out_uop_is_br : _GEN_119 ? _slots_36_io_out_uop_is_br : _GEN_118 ? _slots_35_io_out_uop_is_br : _slots_34_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_120 ? _slots_37_io_out_uop_is_jalr : _GEN_119 ? _slots_36_io_out_uop_is_jalr : _GEN_118 ? _slots_35_io_out_uop_is_jalr : _slots_34_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_120 ? _slots_37_io_out_uop_is_jal : _GEN_119 ? _slots_36_io_out_uop_is_jal : _GEN_118 ? _slots_35_io_out_uop_is_jal : _slots_34_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_120 ? _slots_37_io_out_uop_is_sfb : _GEN_119 ? _slots_36_io_out_uop_is_sfb : _GEN_118 ? _slots_35_io_out_uop_is_sfb : _slots_34_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_120 ? _slots_37_io_out_uop_br_mask : _GEN_119 ? _slots_36_io_out_uop_br_mask : _GEN_118 ? _slots_35_io_out_uop_br_mask : _slots_34_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_120 ? _slots_37_io_out_uop_br_tag : _GEN_119 ? _slots_36_io_out_uop_br_tag : _GEN_118 ? _slots_35_io_out_uop_br_tag : _slots_34_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_120 ? _slots_37_io_out_uop_ftq_idx : _GEN_119 ? _slots_36_io_out_uop_ftq_idx : _GEN_118 ? _slots_35_io_out_uop_ftq_idx : _slots_34_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_120 ? _slots_37_io_out_uop_edge_inst : _GEN_119 ? _slots_36_io_out_uop_edge_inst : _GEN_118 ? _slots_35_io_out_uop_edge_inst : _slots_34_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_120 ? _slots_37_io_out_uop_pc_lob : _GEN_119 ? _slots_36_io_out_uop_pc_lob : _GEN_118 ? _slots_35_io_out_uop_pc_lob : _slots_34_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_120 ? _slots_37_io_out_uop_taken : _GEN_119 ? _slots_36_io_out_uop_taken : _GEN_118 ? _slots_35_io_out_uop_taken : _slots_34_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_120 ? _slots_37_io_out_uop_imm_packed : _GEN_119 ? _slots_36_io_out_uop_imm_packed : _GEN_118 ? _slots_35_io_out_uop_imm_packed : _slots_34_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_120 ? _slots_37_io_out_uop_csr_addr : _GEN_119 ? _slots_36_io_out_uop_csr_addr : _GEN_118 ? _slots_35_io_out_uop_csr_addr : _slots_34_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_120 ? _slots_37_io_out_uop_rob_idx : _GEN_119 ? _slots_36_io_out_uop_rob_idx : _GEN_118 ? _slots_35_io_out_uop_rob_idx : _slots_34_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_120 ? _slots_37_io_out_uop_ldq_idx : _GEN_119 ? _slots_36_io_out_uop_ldq_idx : _GEN_118 ? _slots_35_io_out_uop_ldq_idx : _slots_34_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_120 ? _slots_37_io_out_uop_stq_idx : _GEN_119 ? _slots_36_io_out_uop_stq_idx : _GEN_118 ? _slots_35_io_out_uop_stq_idx : _slots_34_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_120 ? _slots_37_io_out_uop_rxq_idx : _GEN_119 ? _slots_36_io_out_uop_rxq_idx : _GEN_118 ? _slots_35_io_out_uop_rxq_idx : _slots_34_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_120 ? _slots_37_io_out_uop_pdst : _GEN_119 ? _slots_36_io_out_uop_pdst : _GEN_118 ? _slots_35_io_out_uop_pdst : _slots_34_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_120 ? _slots_37_io_out_uop_prs1 : _GEN_119 ? _slots_36_io_out_uop_prs1 : _GEN_118 ? _slots_35_io_out_uop_prs1 : _slots_34_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_120 ? _slots_37_io_out_uop_prs2 : _GEN_119 ? _slots_36_io_out_uop_prs2 : _GEN_118 ? _slots_35_io_out_uop_prs2 : _slots_34_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_120 ? _slots_37_io_out_uop_prs3 : _GEN_119 ? _slots_36_io_out_uop_prs3 : _GEN_118 ? _slots_35_io_out_uop_prs3 : _slots_34_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_120 ? _slots_37_io_out_uop_ppred : _GEN_119 ? _slots_36_io_out_uop_ppred : _GEN_118 ? _slots_35_io_out_uop_ppred : _slots_34_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_120 ? _slots_37_io_out_uop_prs1_busy : _GEN_119 ? _slots_36_io_out_uop_prs1_busy : _GEN_118 ? _slots_35_io_out_uop_prs1_busy : _slots_34_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_120 ? _slots_37_io_out_uop_prs2_busy : _GEN_119 ? _slots_36_io_out_uop_prs2_busy : _GEN_118 ? _slots_35_io_out_uop_prs2_busy : _slots_34_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_120 ? _slots_37_io_out_uop_prs3_busy : _GEN_119 ? _slots_36_io_out_uop_prs3_busy : _GEN_118 ? _slots_35_io_out_uop_prs3_busy : _slots_34_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_120 ? _slots_37_io_out_uop_ppred_busy : _GEN_119 ? _slots_36_io_out_uop_ppred_busy : _GEN_118 ? _slots_35_io_out_uop_ppred_busy : _slots_34_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_120 ? _slots_37_io_out_uop_stale_pdst : _GEN_119 ? _slots_36_io_out_uop_stale_pdst : _GEN_118 ? _slots_35_io_out_uop_stale_pdst : _slots_34_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_120 ? _slots_37_io_out_uop_exception : _GEN_119 ? _slots_36_io_out_uop_exception : _GEN_118 ? _slots_35_io_out_uop_exception : _slots_34_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_120 ? _slots_37_io_out_uop_exc_cause : _GEN_119 ? _slots_36_io_out_uop_exc_cause : _GEN_118 ? _slots_35_io_out_uop_exc_cause : _slots_34_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_120 ? _slots_37_io_out_uop_bypassable : _GEN_119 ? _slots_36_io_out_uop_bypassable : _GEN_118 ? _slots_35_io_out_uop_bypassable : _slots_34_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_120 ? _slots_37_io_out_uop_mem_cmd : _GEN_119 ? _slots_36_io_out_uop_mem_cmd : _GEN_118 ? _slots_35_io_out_uop_mem_cmd : _slots_34_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_120 ? _slots_37_io_out_uop_mem_size : _GEN_119 ? _slots_36_io_out_uop_mem_size : _GEN_118 ? _slots_35_io_out_uop_mem_size : _slots_34_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_120 ? _slots_37_io_out_uop_mem_signed : _GEN_119 ? _slots_36_io_out_uop_mem_signed : _GEN_118 ? _slots_35_io_out_uop_mem_signed : _slots_34_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_120 ? _slots_37_io_out_uop_is_fence : _GEN_119 ? _slots_36_io_out_uop_is_fence : _GEN_118 ? _slots_35_io_out_uop_is_fence : _slots_34_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_120 ? _slots_37_io_out_uop_is_fencei : _GEN_119 ? _slots_36_io_out_uop_is_fencei : _GEN_118 ? _slots_35_io_out_uop_is_fencei : _slots_34_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_120 ? _slots_37_io_out_uop_is_amo : _GEN_119 ? _slots_36_io_out_uop_is_amo : _GEN_118 ? _slots_35_io_out_uop_is_amo : _slots_34_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_120 ? _slots_37_io_out_uop_uses_ldq : _GEN_119 ? _slots_36_io_out_uop_uses_ldq : _GEN_118 ? _slots_35_io_out_uop_uses_ldq : _slots_34_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_120 ? _slots_37_io_out_uop_uses_stq : _GEN_119 ? _slots_36_io_out_uop_uses_stq : _GEN_118 ? _slots_35_io_out_uop_uses_stq : _slots_34_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_120 ? _slots_37_io_out_uop_is_sys_pc2epc : _GEN_119 ? _slots_36_io_out_uop_is_sys_pc2epc : _GEN_118 ? _slots_35_io_out_uop_is_sys_pc2epc : _slots_34_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_120 ? _slots_37_io_out_uop_is_unique : _GEN_119 ? _slots_36_io_out_uop_is_unique : _GEN_118 ? _slots_35_io_out_uop_is_unique : _slots_34_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_120 ? _slots_37_io_out_uop_flush_on_commit : _GEN_119 ? _slots_36_io_out_uop_flush_on_commit : _GEN_118 ? _slots_35_io_out_uop_flush_on_commit : _slots_34_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_120 ? _slots_37_io_out_uop_ldst_is_rs1 : _GEN_119 ? _slots_36_io_out_uop_ldst_is_rs1 : _GEN_118 ? _slots_35_io_out_uop_ldst_is_rs1 : _slots_34_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_120 ? _slots_37_io_out_uop_ldst : _GEN_119 ? _slots_36_io_out_uop_ldst : _GEN_118 ? _slots_35_io_out_uop_ldst : _slots_34_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_120 ? _slots_37_io_out_uop_lrs1 : _GEN_119 ? _slots_36_io_out_uop_lrs1 : _GEN_118 ? _slots_35_io_out_uop_lrs1 : _slots_34_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_120 ? _slots_37_io_out_uop_lrs2 : _GEN_119 ? _slots_36_io_out_uop_lrs2 : _GEN_118 ? _slots_35_io_out_uop_lrs2 : _slots_34_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_120 ? _slots_37_io_out_uop_lrs3 : _GEN_119 ? _slots_36_io_out_uop_lrs3 : _GEN_118 ? _slots_35_io_out_uop_lrs3 : _slots_34_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_120 ? _slots_37_io_out_uop_ldst_val : _GEN_119 ? _slots_36_io_out_uop_ldst_val : _GEN_118 ? _slots_35_io_out_uop_ldst_val : _slots_34_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_120 ? _slots_37_io_out_uop_dst_rtype : _GEN_119 ? _slots_36_io_out_uop_dst_rtype : _GEN_118 ? _slots_35_io_out_uop_dst_rtype : _slots_34_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_120 ? _slots_37_io_out_uop_lrs1_rtype : _GEN_119 ? _slots_36_io_out_uop_lrs1_rtype : _GEN_118 ? _slots_35_io_out_uop_lrs1_rtype : _slots_34_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_120 ? _slots_37_io_out_uop_lrs2_rtype : _GEN_119 ? _slots_36_io_out_uop_lrs2_rtype : _GEN_118 ? _slots_35_io_out_uop_lrs2_rtype : _slots_34_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_120 ? _slots_37_io_out_uop_frs3_en : _GEN_119 ? _slots_36_io_out_uop_frs3_en : _GEN_118 ? _slots_35_io_out_uop_frs3_en : _slots_34_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_120 ? _slots_37_io_out_uop_fp_val : _GEN_119 ? _slots_36_io_out_uop_fp_val : _GEN_118 ? _slots_35_io_out_uop_fp_val : _slots_34_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_120 ? _slots_37_io_out_uop_fp_single : _GEN_119 ? _slots_36_io_out_uop_fp_single : _GEN_118 ? _slots_35_io_out_uop_fp_single : _slots_34_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_120 ? _slots_37_io_out_uop_xcpt_pf_if : _GEN_119 ? _slots_36_io_out_uop_xcpt_pf_if : _GEN_118 ? _slots_35_io_out_uop_xcpt_pf_if : _slots_34_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_120 ? _slots_37_io_out_uop_xcpt_ae_if : _GEN_119 ? _slots_36_io_out_uop_xcpt_ae_if : _GEN_118 ? _slots_35_io_out_uop_xcpt_ae_if : _slots_34_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_120 ? _slots_37_io_out_uop_xcpt_ma_if : _GEN_119 ? _slots_36_io_out_uop_xcpt_ma_if : _GEN_118 ? _slots_35_io_out_uop_xcpt_ma_if : _slots_34_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_120 ? _slots_37_io_out_uop_bp_debug_if : _GEN_119 ? _slots_36_io_out_uop_bp_debug_if : _GEN_118 ? _slots_35_io_out_uop_bp_debug_if : _slots_34_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_120 ? _slots_37_io_out_uop_bp_xcpt_if : _GEN_119 ? _slots_36_io_out_uop_bp_xcpt_if : _GEN_118 ? _slots_35_io_out_uop_bp_xcpt_if : _slots_34_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_120 ? _slots_37_io_out_uop_debug_fsrc : _GEN_119 ? _slots_36_io_out_uop_debug_fsrc : _GEN_118 ? _slots_35_io_out_uop_debug_fsrc : _slots_34_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_120 ? _slots_37_io_out_uop_debug_tsrc : _GEN_119 ? _slots_36_io_out_uop_debug_tsrc : _GEN_118 ? _slots_35_io_out_uop_debug_tsrc : _slots_34_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_33_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_33_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_33_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_33_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_33_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_33_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_33_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_33_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_33_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_33_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_33_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_33_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_33_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_33_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_33_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_33_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_33_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_33_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_33_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_33_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_33_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_33_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_33_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_33_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_33_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_33_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_33_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_33_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_33_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_33_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_33_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_33_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_33_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_33_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_33_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_33_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_33_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_33_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_33_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_33_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_33_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_33_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_33_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_33_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_33_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_33_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_33_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_33_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_33_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_33_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_33_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_33_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_33_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_33_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_33_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_33_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_33_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_33_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_33_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_33_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_33_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_33_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_33_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_33_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_33_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_33_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_33_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_33_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_33_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_33_io_uop_uopc),
    .io_uop_inst                    (_slots_33_io_uop_inst),
    .io_uop_debug_inst              (_slots_33_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_33_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_33_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_33_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_33_io_uop_fu_code),
    .io_uop_iw_state                (_slots_33_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_33_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_33_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_33_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_33_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_33_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_33_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_33_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_33_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_33_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_33_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_33_io_uop_pc_lob),
    .io_uop_taken                   (_slots_33_io_uop_taken),
    .io_uop_imm_packed              (_slots_33_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_33_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_33_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_33_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_33_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_33_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_33_io_uop_pdst),
    .io_uop_prs1                    (_slots_33_io_uop_prs1),
    .io_uop_prs2                    (_slots_33_io_uop_prs2),
    .io_uop_prs3                    (_slots_33_io_uop_prs3),
    .io_uop_ppred                   (_slots_33_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_33_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_33_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_33_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_33_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_33_io_uop_stale_pdst),
    .io_uop_exception               (_slots_33_io_uop_exception),
    .io_uop_exc_cause               (_slots_33_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_33_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_33_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_33_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_33_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_33_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_33_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_33_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_33_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_33_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_33_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_33_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_33_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_33_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_33_io_uop_ldst),
    .io_uop_lrs1                    (_slots_33_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_33_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_33_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_33_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_33_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_33_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_33_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_33_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_33_io_uop_fp_val),
    .io_uop_fp_single               (_slots_33_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_33_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_33_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_33_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_33_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_33_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_33_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_33_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_34 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_34_io_valid),
    .io_will_be_valid               (_slots_34_io_will_be_valid),
    .io_request                     (_slots_34_io_request),
    .io_grant                       (issue_slots_34_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_33),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_34_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_123 ? _slots_38_io_out_uop_uopc : _GEN_122 ? _slots_37_io_out_uop_uopc : _GEN_121 ? _slots_36_io_out_uop_uopc : _slots_35_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_123 ? _slots_38_io_out_uop_inst : _GEN_122 ? _slots_37_io_out_uop_inst : _GEN_121 ? _slots_36_io_out_uop_inst : _slots_35_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_123 ? _slots_38_io_out_uop_debug_inst : _GEN_122 ? _slots_37_io_out_uop_debug_inst : _GEN_121 ? _slots_36_io_out_uop_debug_inst : _slots_35_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_123 ? _slots_38_io_out_uop_is_rvc : _GEN_122 ? _slots_37_io_out_uop_is_rvc : _GEN_121 ? _slots_36_io_out_uop_is_rvc : _slots_35_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_123 ? _slots_38_io_out_uop_debug_pc : _GEN_122 ? _slots_37_io_out_uop_debug_pc : _GEN_121 ? _slots_36_io_out_uop_debug_pc : _slots_35_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_123 ? _slots_38_io_out_uop_iq_type : _GEN_122 ? _slots_37_io_out_uop_iq_type : _GEN_121 ? _slots_36_io_out_uop_iq_type : _slots_35_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_123 ? _slots_38_io_out_uop_fu_code : _GEN_122 ? _slots_37_io_out_uop_fu_code : _GEN_121 ? _slots_36_io_out_uop_fu_code : _slots_35_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_123 ? _slots_38_io_out_uop_iw_state : _GEN_122 ? _slots_37_io_out_uop_iw_state : _GEN_121 ? _slots_36_io_out_uop_iw_state : _slots_35_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_123 ? _slots_38_io_out_uop_iw_p1_poisoned : _GEN_122 ? _slots_37_io_out_uop_iw_p1_poisoned : _GEN_121 ? _slots_36_io_out_uop_iw_p1_poisoned : _slots_35_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_123 ? _slots_38_io_out_uop_iw_p2_poisoned : _GEN_122 ? _slots_37_io_out_uop_iw_p2_poisoned : _GEN_121 ? _slots_36_io_out_uop_iw_p2_poisoned : _slots_35_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_123 ? _slots_38_io_out_uop_is_br : _GEN_122 ? _slots_37_io_out_uop_is_br : _GEN_121 ? _slots_36_io_out_uop_is_br : _slots_35_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_123 ? _slots_38_io_out_uop_is_jalr : _GEN_122 ? _slots_37_io_out_uop_is_jalr : _GEN_121 ? _slots_36_io_out_uop_is_jalr : _slots_35_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_123 ? _slots_38_io_out_uop_is_jal : _GEN_122 ? _slots_37_io_out_uop_is_jal : _GEN_121 ? _slots_36_io_out_uop_is_jal : _slots_35_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_123 ? _slots_38_io_out_uop_is_sfb : _GEN_122 ? _slots_37_io_out_uop_is_sfb : _GEN_121 ? _slots_36_io_out_uop_is_sfb : _slots_35_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_123 ? _slots_38_io_out_uop_br_mask : _GEN_122 ? _slots_37_io_out_uop_br_mask : _GEN_121 ? _slots_36_io_out_uop_br_mask : _slots_35_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_123 ? _slots_38_io_out_uop_br_tag : _GEN_122 ? _slots_37_io_out_uop_br_tag : _GEN_121 ? _slots_36_io_out_uop_br_tag : _slots_35_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_123 ? _slots_38_io_out_uop_ftq_idx : _GEN_122 ? _slots_37_io_out_uop_ftq_idx : _GEN_121 ? _slots_36_io_out_uop_ftq_idx : _slots_35_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_123 ? _slots_38_io_out_uop_edge_inst : _GEN_122 ? _slots_37_io_out_uop_edge_inst : _GEN_121 ? _slots_36_io_out_uop_edge_inst : _slots_35_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_123 ? _slots_38_io_out_uop_pc_lob : _GEN_122 ? _slots_37_io_out_uop_pc_lob : _GEN_121 ? _slots_36_io_out_uop_pc_lob : _slots_35_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_123 ? _slots_38_io_out_uop_taken : _GEN_122 ? _slots_37_io_out_uop_taken : _GEN_121 ? _slots_36_io_out_uop_taken : _slots_35_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_123 ? _slots_38_io_out_uop_imm_packed : _GEN_122 ? _slots_37_io_out_uop_imm_packed : _GEN_121 ? _slots_36_io_out_uop_imm_packed : _slots_35_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_123 ? _slots_38_io_out_uop_csr_addr : _GEN_122 ? _slots_37_io_out_uop_csr_addr : _GEN_121 ? _slots_36_io_out_uop_csr_addr : _slots_35_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_123 ? _slots_38_io_out_uop_rob_idx : _GEN_122 ? _slots_37_io_out_uop_rob_idx : _GEN_121 ? _slots_36_io_out_uop_rob_idx : _slots_35_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_123 ? _slots_38_io_out_uop_ldq_idx : _GEN_122 ? _slots_37_io_out_uop_ldq_idx : _GEN_121 ? _slots_36_io_out_uop_ldq_idx : _slots_35_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_123 ? _slots_38_io_out_uop_stq_idx : _GEN_122 ? _slots_37_io_out_uop_stq_idx : _GEN_121 ? _slots_36_io_out_uop_stq_idx : _slots_35_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_123 ? _slots_38_io_out_uop_rxq_idx : _GEN_122 ? _slots_37_io_out_uop_rxq_idx : _GEN_121 ? _slots_36_io_out_uop_rxq_idx : _slots_35_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_123 ? _slots_38_io_out_uop_pdst : _GEN_122 ? _slots_37_io_out_uop_pdst : _GEN_121 ? _slots_36_io_out_uop_pdst : _slots_35_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_123 ? _slots_38_io_out_uop_prs1 : _GEN_122 ? _slots_37_io_out_uop_prs1 : _GEN_121 ? _slots_36_io_out_uop_prs1 : _slots_35_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_123 ? _slots_38_io_out_uop_prs2 : _GEN_122 ? _slots_37_io_out_uop_prs2 : _GEN_121 ? _slots_36_io_out_uop_prs2 : _slots_35_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_123 ? _slots_38_io_out_uop_prs3 : _GEN_122 ? _slots_37_io_out_uop_prs3 : _GEN_121 ? _slots_36_io_out_uop_prs3 : _slots_35_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_123 ? _slots_38_io_out_uop_ppred : _GEN_122 ? _slots_37_io_out_uop_ppred : _GEN_121 ? _slots_36_io_out_uop_ppred : _slots_35_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_123 ? _slots_38_io_out_uop_prs1_busy : _GEN_122 ? _slots_37_io_out_uop_prs1_busy : _GEN_121 ? _slots_36_io_out_uop_prs1_busy : _slots_35_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_123 ? _slots_38_io_out_uop_prs2_busy : _GEN_122 ? _slots_37_io_out_uop_prs2_busy : _GEN_121 ? _slots_36_io_out_uop_prs2_busy : _slots_35_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_123 ? _slots_38_io_out_uop_prs3_busy : _GEN_122 ? _slots_37_io_out_uop_prs3_busy : _GEN_121 ? _slots_36_io_out_uop_prs3_busy : _slots_35_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_123 ? _slots_38_io_out_uop_ppred_busy : _GEN_122 ? _slots_37_io_out_uop_ppred_busy : _GEN_121 ? _slots_36_io_out_uop_ppred_busy : _slots_35_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_123 ? _slots_38_io_out_uop_stale_pdst : _GEN_122 ? _slots_37_io_out_uop_stale_pdst : _GEN_121 ? _slots_36_io_out_uop_stale_pdst : _slots_35_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_123 ? _slots_38_io_out_uop_exception : _GEN_122 ? _slots_37_io_out_uop_exception : _GEN_121 ? _slots_36_io_out_uop_exception : _slots_35_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_123 ? _slots_38_io_out_uop_exc_cause : _GEN_122 ? _slots_37_io_out_uop_exc_cause : _GEN_121 ? _slots_36_io_out_uop_exc_cause : _slots_35_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_123 ? _slots_38_io_out_uop_bypassable : _GEN_122 ? _slots_37_io_out_uop_bypassable : _GEN_121 ? _slots_36_io_out_uop_bypassable : _slots_35_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_123 ? _slots_38_io_out_uop_mem_cmd : _GEN_122 ? _slots_37_io_out_uop_mem_cmd : _GEN_121 ? _slots_36_io_out_uop_mem_cmd : _slots_35_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_123 ? _slots_38_io_out_uop_mem_size : _GEN_122 ? _slots_37_io_out_uop_mem_size : _GEN_121 ? _slots_36_io_out_uop_mem_size : _slots_35_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_123 ? _slots_38_io_out_uop_mem_signed : _GEN_122 ? _slots_37_io_out_uop_mem_signed : _GEN_121 ? _slots_36_io_out_uop_mem_signed : _slots_35_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_123 ? _slots_38_io_out_uop_is_fence : _GEN_122 ? _slots_37_io_out_uop_is_fence : _GEN_121 ? _slots_36_io_out_uop_is_fence : _slots_35_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_123 ? _slots_38_io_out_uop_is_fencei : _GEN_122 ? _slots_37_io_out_uop_is_fencei : _GEN_121 ? _slots_36_io_out_uop_is_fencei : _slots_35_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_123 ? _slots_38_io_out_uop_is_amo : _GEN_122 ? _slots_37_io_out_uop_is_amo : _GEN_121 ? _slots_36_io_out_uop_is_amo : _slots_35_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_123 ? _slots_38_io_out_uop_uses_ldq : _GEN_122 ? _slots_37_io_out_uop_uses_ldq : _GEN_121 ? _slots_36_io_out_uop_uses_ldq : _slots_35_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_123 ? _slots_38_io_out_uop_uses_stq : _GEN_122 ? _slots_37_io_out_uop_uses_stq : _GEN_121 ? _slots_36_io_out_uop_uses_stq : _slots_35_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_123 ? _slots_38_io_out_uop_is_sys_pc2epc : _GEN_122 ? _slots_37_io_out_uop_is_sys_pc2epc : _GEN_121 ? _slots_36_io_out_uop_is_sys_pc2epc : _slots_35_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_123 ? _slots_38_io_out_uop_is_unique : _GEN_122 ? _slots_37_io_out_uop_is_unique : _GEN_121 ? _slots_36_io_out_uop_is_unique : _slots_35_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_123 ? _slots_38_io_out_uop_flush_on_commit : _GEN_122 ? _slots_37_io_out_uop_flush_on_commit : _GEN_121 ? _slots_36_io_out_uop_flush_on_commit : _slots_35_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_123 ? _slots_38_io_out_uop_ldst_is_rs1 : _GEN_122 ? _slots_37_io_out_uop_ldst_is_rs1 : _GEN_121 ? _slots_36_io_out_uop_ldst_is_rs1 : _slots_35_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_123 ? _slots_38_io_out_uop_ldst : _GEN_122 ? _slots_37_io_out_uop_ldst : _GEN_121 ? _slots_36_io_out_uop_ldst : _slots_35_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_123 ? _slots_38_io_out_uop_lrs1 : _GEN_122 ? _slots_37_io_out_uop_lrs1 : _GEN_121 ? _slots_36_io_out_uop_lrs1 : _slots_35_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_123 ? _slots_38_io_out_uop_lrs2 : _GEN_122 ? _slots_37_io_out_uop_lrs2 : _GEN_121 ? _slots_36_io_out_uop_lrs2 : _slots_35_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_123 ? _slots_38_io_out_uop_lrs3 : _GEN_122 ? _slots_37_io_out_uop_lrs3 : _GEN_121 ? _slots_36_io_out_uop_lrs3 : _slots_35_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_123 ? _slots_38_io_out_uop_ldst_val : _GEN_122 ? _slots_37_io_out_uop_ldst_val : _GEN_121 ? _slots_36_io_out_uop_ldst_val : _slots_35_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_123 ? _slots_38_io_out_uop_dst_rtype : _GEN_122 ? _slots_37_io_out_uop_dst_rtype : _GEN_121 ? _slots_36_io_out_uop_dst_rtype : _slots_35_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_123 ? _slots_38_io_out_uop_lrs1_rtype : _GEN_122 ? _slots_37_io_out_uop_lrs1_rtype : _GEN_121 ? _slots_36_io_out_uop_lrs1_rtype : _slots_35_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_123 ? _slots_38_io_out_uop_lrs2_rtype : _GEN_122 ? _slots_37_io_out_uop_lrs2_rtype : _GEN_121 ? _slots_36_io_out_uop_lrs2_rtype : _slots_35_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_123 ? _slots_38_io_out_uop_frs3_en : _GEN_122 ? _slots_37_io_out_uop_frs3_en : _GEN_121 ? _slots_36_io_out_uop_frs3_en : _slots_35_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_123 ? _slots_38_io_out_uop_fp_val : _GEN_122 ? _slots_37_io_out_uop_fp_val : _GEN_121 ? _slots_36_io_out_uop_fp_val : _slots_35_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_123 ? _slots_38_io_out_uop_fp_single : _GEN_122 ? _slots_37_io_out_uop_fp_single : _GEN_121 ? _slots_36_io_out_uop_fp_single : _slots_35_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_123 ? _slots_38_io_out_uop_xcpt_pf_if : _GEN_122 ? _slots_37_io_out_uop_xcpt_pf_if : _GEN_121 ? _slots_36_io_out_uop_xcpt_pf_if : _slots_35_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_123 ? _slots_38_io_out_uop_xcpt_ae_if : _GEN_122 ? _slots_37_io_out_uop_xcpt_ae_if : _GEN_121 ? _slots_36_io_out_uop_xcpt_ae_if : _slots_35_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_123 ? _slots_38_io_out_uop_xcpt_ma_if : _GEN_122 ? _slots_37_io_out_uop_xcpt_ma_if : _GEN_121 ? _slots_36_io_out_uop_xcpt_ma_if : _slots_35_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_123 ? _slots_38_io_out_uop_bp_debug_if : _GEN_122 ? _slots_37_io_out_uop_bp_debug_if : _GEN_121 ? _slots_36_io_out_uop_bp_debug_if : _slots_35_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_123 ? _slots_38_io_out_uop_bp_xcpt_if : _GEN_122 ? _slots_37_io_out_uop_bp_xcpt_if : _GEN_121 ? _slots_36_io_out_uop_bp_xcpt_if : _slots_35_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_123 ? _slots_38_io_out_uop_debug_fsrc : _GEN_122 ? _slots_37_io_out_uop_debug_fsrc : _GEN_121 ? _slots_36_io_out_uop_debug_fsrc : _slots_35_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_123 ? _slots_38_io_out_uop_debug_tsrc : _GEN_122 ? _slots_37_io_out_uop_debug_tsrc : _GEN_121 ? _slots_36_io_out_uop_debug_tsrc : _slots_35_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_34_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_34_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_34_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_34_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_34_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_34_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_34_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_34_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_34_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_34_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_34_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_34_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_34_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_34_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_34_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_34_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_34_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_34_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_34_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_34_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_34_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_34_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_34_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_34_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_34_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_34_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_34_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_34_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_34_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_34_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_34_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_34_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_34_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_34_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_34_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_34_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_34_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_34_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_34_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_34_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_34_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_34_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_34_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_34_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_34_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_34_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_34_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_34_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_34_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_34_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_34_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_34_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_34_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_34_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_34_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_34_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_34_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_34_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_34_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_34_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_34_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_34_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_34_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_34_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_34_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_34_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_34_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_34_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_34_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_34_io_uop_uopc),
    .io_uop_inst                    (_slots_34_io_uop_inst),
    .io_uop_debug_inst              (_slots_34_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_34_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_34_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_34_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_34_io_uop_fu_code),
    .io_uop_iw_state                (_slots_34_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_34_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_34_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_34_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_34_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_34_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_34_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_34_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_34_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_34_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_34_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_34_io_uop_pc_lob),
    .io_uop_taken                   (_slots_34_io_uop_taken),
    .io_uop_imm_packed              (_slots_34_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_34_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_34_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_34_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_34_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_34_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_34_io_uop_pdst),
    .io_uop_prs1                    (_slots_34_io_uop_prs1),
    .io_uop_prs2                    (_slots_34_io_uop_prs2),
    .io_uop_prs3                    (_slots_34_io_uop_prs3),
    .io_uop_ppred                   (_slots_34_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_34_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_34_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_34_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_34_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_34_io_uop_stale_pdst),
    .io_uop_exception               (_slots_34_io_uop_exception),
    .io_uop_exc_cause               (_slots_34_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_34_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_34_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_34_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_34_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_34_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_34_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_34_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_34_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_34_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_34_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_34_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_34_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_34_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_34_io_uop_ldst),
    .io_uop_lrs1                    (_slots_34_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_34_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_34_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_34_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_34_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_34_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_34_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_34_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_34_io_uop_fp_val),
    .io_uop_fp_single               (_slots_34_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_34_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_34_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_34_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_34_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_34_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_34_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_34_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_35 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_35_io_valid),
    .io_will_be_valid               (_slots_35_io_will_be_valid),
    .io_request                     (_slots_35_io_request),
    .io_grant                       (issue_slots_35_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_34),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_35_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_126 ? _slots_39_io_out_uop_uopc : _GEN_125 ? _slots_38_io_out_uop_uopc : _GEN_124 ? _slots_37_io_out_uop_uopc : _slots_36_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_126 ? _slots_39_io_out_uop_inst : _GEN_125 ? _slots_38_io_out_uop_inst : _GEN_124 ? _slots_37_io_out_uop_inst : _slots_36_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_126 ? _slots_39_io_out_uop_debug_inst : _GEN_125 ? _slots_38_io_out_uop_debug_inst : _GEN_124 ? _slots_37_io_out_uop_debug_inst : _slots_36_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_126 ? _slots_39_io_out_uop_is_rvc : _GEN_125 ? _slots_38_io_out_uop_is_rvc : _GEN_124 ? _slots_37_io_out_uop_is_rvc : _slots_36_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_126 ? _slots_39_io_out_uop_debug_pc : _GEN_125 ? _slots_38_io_out_uop_debug_pc : _GEN_124 ? _slots_37_io_out_uop_debug_pc : _slots_36_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_126 ? _slots_39_io_out_uop_iq_type : _GEN_125 ? _slots_38_io_out_uop_iq_type : _GEN_124 ? _slots_37_io_out_uop_iq_type : _slots_36_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_126 ? _slots_39_io_out_uop_fu_code : _GEN_125 ? _slots_38_io_out_uop_fu_code : _GEN_124 ? _slots_37_io_out_uop_fu_code : _slots_36_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_126 ? _slots_39_io_out_uop_iw_state : _GEN_125 ? _slots_38_io_out_uop_iw_state : _GEN_124 ? _slots_37_io_out_uop_iw_state : _slots_36_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_126 ? _slots_39_io_out_uop_iw_p1_poisoned : _GEN_125 ? _slots_38_io_out_uop_iw_p1_poisoned : _GEN_124 ? _slots_37_io_out_uop_iw_p1_poisoned : _slots_36_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_126 ? _slots_39_io_out_uop_iw_p2_poisoned : _GEN_125 ? _slots_38_io_out_uop_iw_p2_poisoned : _GEN_124 ? _slots_37_io_out_uop_iw_p2_poisoned : _slots_36_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_126 ? _slots_39_io_out_uop_is_br : _GEN_125 ? _slots_38_io_out_uop_is_br : _GEN_124 ? _slots_37_io_out_uop_is_br : _slots_36_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_126 ? _slots_39_io_out_uop_is_jalr : _GEN_125 ? _slots_38_io_out_uop_is_jalr : _GEN_124 ? _slots_37_io_out_uop_is_jalr : _slots_36_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_126 ? _slots_39_io_out_uop_is_jal : _GEN_125 ? _slots_38_io_out_uop_is_jal : _GEN_124 ? _slots_37_io_out_uop_is_jal : _slots_36_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_126 ? _slots_39_io_out_uop_is_sfb : _GEN_125 ? _slots_38_io_out_uop_is_sfb : _GEN_124 ? _slots_37_io_out_uop_is_sfb : _slots_36_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_126 ? _slots_39_io_out_uop_br_mask : _GEN_125 ? _slots_38_io_out_uop_br_mask : _GEN_124 ? _slots_37_io_out_uop_br_mask : _slots_36_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_126 ? _slots_39_io_out_uop_br_tag : _GEN_125 ? _slots_38_io_out_uop_br_tag : _GEN_124 ? _slots_37_io_out_uop_br_tag : _slots_36_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_126 ? _slots_39_io_out_uop_ftq_idx : _GEN_125 ? _slots_38_io_out_uop_ftq_idx : _GEN_124 ? _slots_37_io_out_uop_ftq_idx : _slots_36_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_126 ? _slots_39_io_out_uop_edge_inst : _GEN_125 ? _slots_38_io_out_uop_edge_inst : _GEN_124 ? _slots_37_io_out_uop_edge_inst : _slots_36_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_126 ? _slots_39_io_out_uop_pc_lob : _GEN_125 ? _slots_38_io_out_uop_pc_lob : _GEN_124 ? _slots_37_io_out_uop_pc_lob : _slots_36_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_126 ? _slots_39_io_out_uop_taken : _GEN_125 ? _slots_38_io_out_uop_taken : _GEN_124 ? _slots_37_io_out_uop_taken : _slots_36_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_126 ? _slots_39_io_out_uop_imm_packed : _GEN_125 ? _slots_38_io_out_uop_imm_packed : _GEN_124 ? _slots_37_io_out_uop_imm_packed : _slots_36_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_126 ? _slots_39_io_out_uop_csr_addr : _GEN_125 ? _slots_38_io_out_uop_csr_addr : _GEN_124 ? _slots_37_io_out_uop_csr_addr : _slots_36_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_126 ? _slots_39_io_out_uop_rob_idx : _GEN_125 ? _slots_38_io_out_uop_rob_idx : _GEN_124 ? _slots_37_io_out_uop_rob_idx : _slots_36_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_126 ? _slots_39_io_out_uop_ldq_idx : _GEN_125 ? _slots_38_io_out_uop_ldq_idx : _GEN_124 ? _slots_37_io_out_uop_ldq_idx : _slots_36_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_126 ? _slots_39_io_out_uop_stq_idx : _GEN_125 ? _slots_38_io_out_uop_stq_idx : _GEN_124 ? _slots_37_io_out_uop_stq_idx : _slots_36_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_126 ? _slots_39_io_out_uop_rxq_idx : _GEN_125 ? _slots_38_io_out_uop_rxq_idx : _GEN_124 ? _slots_37_io_out_uop_rxq_idx : _slots_36_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_126 ? _slots_39_io_out_uop_pdst : _GEN_125 ? _slots_38_io_out_uop_pdst : _GEN_124 ? _slots_37_io_out_uop_pdst : _slots_36_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_126 ? _slots_39_io_out_uop_prs1 : _GEN_125 ? _slots_38_io_out_uop_prs1 : _GEN_124 ? _slots_37_io_out_uop_prs1 : _slots_36_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_126 ? _slots_39_io_out_uop_prs2 : _GEN_125 ? _slots_38_io_out_uop_prs2 : _GEN_124 ? _slots_37_io_out_uop_prs2 : _slots_36_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_126 ? _slots_39_io_out_uop_prs3 : _GEN_125 ? _slots_38_io_out_uop_prs3 : _GEN_124 ? _slots_37_io_out_uop_prs3 : _slots_36_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_126 ? _slots_39_io_out_uop_ppred : _GEN_125 ? _slots_38_io_out_uop_ppred : _GEN_124 ? _slots_37_io_out_uop_ppred : _slots_36_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_126 ? _slots_39_io_out_uop_prs1_busy : _GEN_125 ? _slots_38_io_out_uop_prs1_busy : _GEN_124 ? _slots_37_io_out_uop_prs1_busy : _slots_36_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_126 ? _slots_39_io_out_uop_prs2_busy : _GEN_125 ? _slots_38_io_out_uop_prs2_busy : _GEN_124 ? _slots_37_io_out_uop_prs2_busy : _slots_36_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_126 ? _slots_39_io_out_uop_prs3_busy : _GEN_125 ? _slots_38_io_out_uop_prs3_busy : _GEN_124 ? _slots_37_io_out_uop_prs3_busy : _slots_36_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_126 ? _slots_39_io_out_uop_ppred_busy : _GEN_125 ? _slots_38_io_out_uop_ppred_busy : _GEN_124 ? _slots_37_io_out_uop_ppred_busy : _slots_36_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_126 ? _slots_39_io_out_uop_stale_pdst : _GEN_125 ? _slots_38_io_out_uop_stale_pdst : _GEN_124 ? _slots_37_io_out_uop_stale_pdst : _slots_36_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_126 ? _slots_39_io_out_uop_exception : _GEN_125 ? _slots_38_io_out_uop_exception : _GEN_124 ? _slots_37_io_out_uop_exception : _slots_36_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_126 ? _slots_39_io_out_uop_exc_cause : _GEN_125 ? _slots_38_io_out_uop_exc_cause : _GEN_124 ? _slots_37_io_out_uop_exc_cause : _slots_36_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_126 ? _slots_39_io_out_uop_bypassable : _GEN_125 ? _slots_38_io_out_uop_bypassable : _GEN_124 ? _slots_37_io_out_uop_bypassable : _slots_36_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_126 ? _slots_39_io_out_uop_mem_cmd : _GEN_125 ? _slots_38_io_out_uop_mem_cmd : _GEN_124 ? _slots_37_io_out_uop_mem_cmd : _slots_36_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_126 ? _slots_39_io_out_uop_mem_size : _GEN_125 ? _slots_38_io_out_uop_mem_size : _GEN_124 ? _slots_37_io_out_uop_mem_size : _slots_36_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_126 ? _slots_39_io_out_uop_mem_signed : _GEN_125 ? _slots_38_io_out_uop_mem_signed : _GEN_124 ? _slots_37_io_out_uop_mem_signed : _slots_36_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_126 ? _slots_39_io_out_uop_is_fence : _GEN_125 ? _slots_38_io_out_uop_is_fence : _GEN_124 ? _slots_37_io_out_uop_is_fence : _slots_36_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_126 ? _slots_39_io_out_uop_is_fencei : _GEN_125 ? _slots_38_io_out_uop_is_fencei : _GEN_124 ? _slots_37_io_out_uop_is_fencei : _slots_36_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_126 ? _slots_39_io_out_uop_is_amo : _GEN_125 ? _slots_38_io_out_uop_is_amo : _GEN_124 ? _slots_37_io_out_uop_is_amo : _slots_36_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_126 ? _slots_39_io_out_uop_uses_ldq : _GEN_125 ? _slots_38_io_out_uop_uses_ldq : _GEN_124 ? _slots_37_io_out_uop_uses_ldq : _slots_36_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_126 ? _slots_39_io_out_uop_uses_stq : _GEN_125 ? _slots_38_io_out_uop_uses_stq : _GEN_124 ? _slots_37_io_out_uop_uses_stq : _slots_36_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_126 ? _slots_39_io_out_uop_is_sys_pc2epc : _GEN_125 ? _slots_38_io_out_uop_is_sys_pc2epc : _GEN_124 ? _slots_37_io_out_uop_is_sys_pc2epc : _slots_36_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_126 ? _slots_39_io_out_uop_is_unique : _GEN_125 ? _slots_38_io_out_uop_is_unique : _GEN_124 ? _slots_37_io_out_uop_is_unique : _slots_36_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_126 ? _slots_39_io_out_uop_flush_on_commit : _GEN_125 ? _slots_38_io_out_uop_flush_on_commit : _GEN_124 ? _slots_37_io_out_uop_flush_on_commit : _slots_36_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_126 ? _slots_39_io_out_uop_ldst_is_rs1 : _GEN_125 ? _slots_38_io_out_uop_ldst_is_rs1 : _GEN_124 ? _slots_37_io_out_uop_ldst_is_rs1 : _slots_36_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_126 ? _slots_39_io_out_uop_ldst : _GEN_125 ? _slots_38_io_out_uop_ldst : _GEN_124 ? _slots_37_io_out_uop_ldst : _slots_36_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_126 ? _slots_39_io_out_uop_lrs1 : _GEN_125 ? _slots_38_io_out_uop_lrs1 : _GEN_124 ? _slots_37_io_out_uop_lrs1 : _slots_36_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_126 ? _slots_39_io_out_uop_lrs2 : _GEN_125 ? _slots_38_io_out_uop_lrs2 : _GEN_124 ? _slots_37_io_out_uop_lrs2 : _slots_36_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_126 ? _slots_39_io_out_uop_lrs3 : _GEN_125 ? _slots_38_io_out_uop_lrs3 : _GEN_124 ? _slots_37_io_out_uop_lrs3 : _slots_36_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_126 ? _slots_39_io_out_uop_ldst_val : _GEN_125 ? _slots_38_io_out_uop_ldst_val : _GEN_124 ? _slots_37_io_out_uop_ldst_val : _slots_36_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_126 ? _slots_39_io_out_uop_dst_rtype : _GEN_125 ? _slots_38_io_out_uop_dst_rtype : _GEN_124 ? _slots_37_io_out_uop_dst_rtype : _slots_36_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_126 ? _slots_39_io_out_uop_lrs1_rtype : _GEN_125 ? _slots_38_io_out_uop_lrs1_rtype : _GEN_124 ? _slots_37_io_out_uop_lrs1_rtype : _slots_36_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_126 ? _slots_39_io_out_uop_lrs2_rtype : _GEN_125 ? _slots_38_io_out_uop_lrs2_rtype : _GEN_124 ? _slots_37_io_out_uop_lrs2_rtype : _slots_36_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_126 ? _slots_39_io_out_uop_frs3_en : _GEN_125 ? _slots_38_io_out_uop_frs3_en : _GEN_124 ? _slots_37_io_out_uop_frs3_en : _slots_36_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_126 ? _slots_39_io_out_uop_fp_val : _GEN_125 ? _slots_38_io_out_uop_fp_val : _GEN_124 ? _slots_37_io_out_uop_fp_val : _slots_36_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_126 ? _slots_39_io_out_uop_fp_single : _GEN_125 ? _slots_38_io_out_uop_fp_single : _GEN_124 ? _slots_37_io_out_uop_fp_single : _slots_36_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_126 ? _slots_39_io_out_uop_xcpt_pf_if : _GEN_125 ? _slots_38_io_out_uop_xcpt_pf_if : _GEN_124 ? _slots_37_io_out_uop_xcpt_pf_if : _slots_36_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_126 ? _slots_39_io_out_uop_xcpt_ae_if : _GEN_125 ? _slots_38_io_out_uop_xcpt_ae_if : _GEN_124 ? _slots_37_io_out_uop_xcpt_ae_if : _slots_36_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_126 ? _slots_39_io_out_uop_xcpt_ma_if : _GEN_125 ? _slots_38_io_out_uop_xcpt_ma_if : _GEN_124 ? _slots_37_io_out_uop_xcpt_ma_if : _slots_36_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_126 ? _slots_39_io_out_uop_bp_debug_if : _GEN_125 ? _slots_38_io_out_uop_bp_debug_if : _GEN_124 ? _slots_37_io_out_uop_bp_debug_if : _slots_36_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_126 ? _slots_39_io_out_uop_bp_xcpt_if : _GEN_125 ? _slots_38_io_out_uop_bp_xcpt_if : _GEN_124 ? _slots_37_io_out_uop_bp_xcpt_if : _slots_36_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_126 ? _slots_39_io_out_uop_debug_fsrc : _GEN_125 ? _slots_38_io_out_uop_debug_fsrc : _GEN_124 ? _slots_37_io_out_uop_debug_fsrc : _slots_36_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_126 ? _slots_39_io_out_uop_debug_tsrc : _GEN_125 ? _slots_38_io_out_uop_debug_tsrc : _GEN_124 ? _slots_37_io_out_uop_debug_tsrc : _slots_36_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_35_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_35_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_35_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_35_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_35_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_35_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_35_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_35_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_35_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_35_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_35_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_35_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_35_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_35_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_35_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_35_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_35_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_35_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_35_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_35_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_35_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_35_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_35_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_35_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_35_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_35_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_35_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_35_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_35_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_35_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_35_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_35_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_35_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_35_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_35_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_35_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_35_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_35_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_35_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_35_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_35_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_35_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_35_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_35_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_35_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_35_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_35_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_35_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_35_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_35_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_35_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_35_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_35_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_35_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_35_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_35_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_35_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_35_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_35_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_35_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_35_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_35_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_35_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_35_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_35_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_35_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_35_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_35_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_35_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_35_io_uop_uopc),
    .io_uop_inst                    (_slots_35_io_uop_inst),
    .io_uop_debug_inst              (_slots_35_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_35_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_35_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_35_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_35_io_uop_fu_code),
    .io_uop_iw_state                (_slots_35_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_35_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_35_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_35_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_35_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_35_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_35_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_35_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_35_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_35_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_35_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_35_io_uop_pc_lob),
    .io_uop_taken                   (_slots_35_io_uop_taken),
    .io_uop_imm_packed              (_slots_35_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_35_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_35_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_35_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_35_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_35_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_35_io_uop_pdst),
    .io_uop_prs1                    (_slots_35_io_uop_prs1),
    .io_uop_prs2                    (_slots_35_io_uop_prs2),
    .io_uop_prs3                    (_slots_35_io_uop_prs3),
    .io_uop_ppred                   (_slots_35_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_35_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_35_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_35_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_35_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_35_io_uop_stale_pdst),
    .io_uop_exception               (_slots_35_io_uop_exception),
    .io_uop_exc_cause               (_slots_35_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_35_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_35_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_35_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_35_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_35_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_35_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_35_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_35_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_35_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_35_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_35_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_35_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_35_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_35_io_uop_ldst),
    .io_uop_lrs1                    (_slots_35_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_35_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_35_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_35_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_35_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_35_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_35_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_35_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_35_io_uop_fp_val),
    .io_uop_fp_single               (_slots_35_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_35_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_35_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_35_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_35_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_35_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_35_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_35_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_36 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_36_io_valid),
    .io_will_be_valid               (_slots_36_io_will_be_valid),
    .io_request                     (_slots_36_io_request),
    .io_grant                       (issue_slots_36_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_35),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_36_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_129 ? io_dis_uops_0_bits_uopc : _GEN_128 ? _slots_39_io_out_uop_uopc : _GEN_127 ? _slots_38_io_out_uop_uopc : _slots_37_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_129 ? io_dis_uops_0_bits_inst : _GEN_128 ? _slots_39_io_out_uop_inst : _GEN_127 ? _slots_38_io_out_uop_inst : _slots_37_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_129 ? io_dis_uops_0_bits_debug_inst : _GEN_128 ? _slots_39_io_out_uop_debug_inst : _GEN_127 ? _slots_38_io_out_uop_debug_inst : _slots_37_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_129 ? io_dis_uops_0_bits_is_rvc : _GEN_128 ? _slots_39_io_out_uop_is_rvc : _GEN_127 ? _slots_38_io_out_uop_is_rvc : _slots_37_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_129 ? io_dis_uops_0_bits_debug_pc : _GEN_128 ? _slots_39_io_out_uop_debug_pc : _GEN_127 ? _slots_38_io_out_uop_debug_pc : _slots_37_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_129 ? io_dis_uops_0_bits_iq_type : _GEN_128 ? _slots_39_io_out_uop_iq_type : _GEN_127 ? _slots_38_io_out_uop_iq_type : _slots_37_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_129 ? io_dis_uops_0_bits_fu_code : _GEN_128 ? _slots_39_io_out_uop_fu_code : _GEN_127 ? _slots_38_io_out_uop_fu_code : _slots_37_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_129 ? _GEN_1 : _GEN_128 ? _slots_39_io_out_uop_iw_state : _GEN_127 ? _slots_38_io_out_uop_iw_state : _slots_37_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_129 & (_GEN_128 ? _slots_39_io_out_uop_iw_p1_poisoned : _GEN_127 ? _slots_38_io_out_uop_iw_p1_poisoned : _slots_37_io_out_uop_iw_p1_poisoned)),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_129 & (_GEN_128 ? _slots_39_io_out_uop_iw_p2_poisoned : _GEN_127 ? _slots_38_io_out_uop_iw_p2_poisoned : _slots_37_io_out_uop_iw_p2_poisoned)),
    .io_in_uop_bits_is_br           (_GEN_129 ? io_dis_uops_0_bits_is_br : _GEN_128 ? _slots_39_io_out_uop_is_br : _GEN_127 ? _slots_38_io_out_uop_is_br : _slots_37_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_129 ? io_dis_uops_0_bits_is_jalr : _GEN_128 ? _slots_39_io_out_uop_is_jalr : _GEN_127 ? _slots_38_io_out_uop_is_jalr : _slots_37_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_129 ? io_dis_uops_0_bits_is_jal : _GEN_128 ? _slots_39_io_out_uop_is_jal : _GEN_127 ? _slots_38_io_out_uop_is_jal : _slots_37_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_129 ? io_dis_uops_0_bits_is_sfb : _GEN_128 ? _slots_39_io_out_uop_is_sfb : _GEN_127 ? _slots_38_io_out_uop_is_sfb : _slots_37_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_129 ? io_dis_uops_0_bits_br_mask : _GEN_128 ? _slots_39_io_out_uop_br_mask : _GEN_127 ? _slots_38_io_out_uop_br_mask : _slots_37_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_129 ? io_dis_uops_0_bits_br_tag : _GEN_128 ? _slots_39_io_out_uop_br_tag : _GEN_127 ? _slots_38_io_out_uop_br_tag : _slots_37_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_129 ? io_dis_uops_0_bits_ftq_idx : _GEN_128 ? _slots_39_io_out_uop_ftq_idx : _GEN_127 ? _slots_38_io_out_uop_ftq_idx : _slots_37_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_129 ? io_dis_uops_0_bits_edge_inst : _GEN_128 ? _slots_39_io_out_uop_edge_inst : _GEN_127 ? _slots_38_io_out_uop_edge_inst : _slots_37_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_129 ? io_dis_uops_0_bits_pc_lob : _GEN_128 ? _slots_39_io_out_uop_pc_lob : _GEN_127 ? _slots_38_io_out_uop_pc_lob : _slots_37_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_129 ? io_dis_uops_0_bits_taken : _GEN_128 ? _slots_39_io_out_uop_taken : _GEN_127 ? _slots_38_io_out_uop_taken : _slots_37_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_129 ? io_dis_uops_0_bits_imm_packed : _GEN_128 ? _slots_39_io_out_uop_imm_packed : _GEN_127 ? _slots_38_io_out_uop_imm_packed : _slots_37_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_129 ? io_dis_uops_0_bits_csr_addr : _GEN_128 ? _slots_39_io_out_uop_csr_addr : _GEN_127 ? _slots_38_io_out_uop_csr_addr : _slots_37_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_129 ? io_dis_uops_0_bits_rob_idx : _GEN_128 ? _slots_39_io_out_uop_rob_idx : _GEN_127 ? _slots_38_io_out_uop_rob_idx : _slots_37_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_129 ? io_dis_uops_0_bits_ldq_idx : _GEN_128 ? _slots_39_io_out_uop_ldq_idx : _GEN_127 ? _slots_38_io_out_uop_ldq_idx : _slots_37_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_129 ? io_dis_uops_0_bits_stq_idx : _GEN_128 ? _slots_39_io_out_uop_stq_idx : _GEN_127 ? _slots_38_io_out_uop_stq_idx : _slots_37_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_129 ? io_dis_uops_0_bits_rxq_idx : _GEN_128 ? _slots_39_io_out_uop_rxq_idx : _GEN_127 ? _slots_38_io_out_uop_rxq_idx : _slots_37_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_129 ? io_dis_uops_0_bits_pdst : _GEN_128 ? _slots_39_io_out_uop_pdst : _GEN_127 ? _slots_38_io_out_uop_pdst : _slots_37_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_129 ? io_dis_uops_0_bits_prs1 : _GEN_128 ? _slots_39_io_out_uop_prs1 : _GEN_127 ? _slots_38_io_out_uop_prs1 : _slots_37_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_129 ? io_dis_uops_0_bits_prs2 : _GEN_128 ? _slots_39_io_out_uop_prs2 : _GEN_127 ? _slots_38_io_out_uop_prs2 : _slots_37_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_129 ? io_dis_uops_0_bits_prs3 : _GEN_128 ? _slots_39_io_out_uop_prs3 : _GEN_127 ? _slots_38_io_out_uop_prs3 : _slots_37_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_129 ? 6'h0 : _GEN_128 ? _slots_39_io_out_uop_ppred : _GEN_127 ? _slots_38_io_out_uop_ppred : _slots_37_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_129 ? io_dis_uops_0_bits_prs1_busy : _GEN_128 ? _slots_39_io_out_uop_prs1_busy : _GEN_127 ? _slots_38_io_out_uop_prs1_busy : _slots_37_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_129 ? _GEN_4 : _GEN_128 ? _slots_39_io_out_uop_prs2_busy : _GEN_127 ? _slots_38_io_out_uop_prs2_busy : _slots_37_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_129 & (_GEN_128 ? _slots_39_io_out_uop_prs3_busy : _GEN_127 ? _slots_38_io_out_uop_prs3_busy : _slots_37_io_out_uop_prs3_busy)),
    .io_in_uop_bits_ppred_busy      (~_GEN_129 & (_GEN_128 ? _slots_39_io_out_uop_ppred_busy : _GEN_127 ? _slots_38_io_out_uop_ppred_busy : _slots_37_io_out_uop_ppred_busy)),
    .io_in_uop_bits_stale_pdst      (_GEN_129 ? io_dis_uops_0_bits_stale_pdst : _GEN_128 ? _slots_39_io_out_uop_stale_pdst : _GEN_127 ? _slots_38_io_out_uop_stale_pdst : _slots_37_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_129 ? io_dis_uops_0_bits_exception : _GEN_128 ? _slots_39_io_out_uop_exception : _GEN_127 ? _slots_38_io_out_uop_exception : _slots_37_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_129 ? io_dis_uops_0_bits_exc_cause : _GEN_128 ? _slots_39_io_out_uop_exc_cause : _GEN_127 ? _slots_38_io_out_uop_exc_cause : _slots_37_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_129 ? io_dis_uops_0_bits_bypassable : _GEN_128 ? _slots_39_io_out_uop_bypassable : _GEN_127 ? _slots_38_io_out_uop_bypassable : _slots_37_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_129 ? io_dis_uops_0_bits_mem_cmd : _GEN_128 ? _slots_39_io_out_uop_mem_cmd : _GEN_127 ? _slots_38_io_out_uop_mem_cmd : _slots_37_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_129 ? io_dis_uops_0_bits_mem_size : _GEN_128 ? _slots_39_io_out_uop_mem_size : _GEN_127 ? _slots_38_io_out_uop_mem_size : _slots_37_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_129 ? io_dis_uops_0_bits_mem_signed : _GEN_128 ? _slots_39_io_out_uop_mem_signed : _GEN_127 ? _slots_38_io_out_uop_mem_signed : _slots_37_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_129 ? io_dis_uops_0_bits_is_fence : _GEN_128 ? _slots_39_io_out_uop_is_fence : _GEN_127 ? _slots_38_io_out_uop_is_fence : _slots_37_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_129 ? io_dis_uops_0_bits_is_fencei : _GEN_128 ? _slots_39_io_out_uop_is_fencei : _GEN_127 ? _slots_38_io_out_uop_is_fencei : _slots_37_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_129 ? io_dis_uops_0_bits_is_amo : _GEN_128 ? _slots_39_io_out_uop_is_amo : _GEN_127 ? _slots_38_io_out_uop_is_amo : _slots_37_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_129 ? io_dis_uops_0_bits_uses_ldq : _GEN_128 ? _slots_39_io_out_uop_uses_ldq : _GEN_127 ? _slots_38_io_out_uop_uses_ldq : _slots_37_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_129 ? io_dis_uops_0_bits_uses_stq : _GEN_128 ? _slots_39_io_out_uop_uses_stq : _GEN_127 ? _slots_38_io_out_uop_uses_stq : _slots_37_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_129 ? io_dis_uops_0_bits_is_sys_pc2epc : _GEN_128 ? _slots_39_io_out_uop_is_sys_pc2epc : _GEN_127 ? _slots_38_io_out_uop_is_sys_pc2epc : _slots_37_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_129 ? io_dis_uops_0_bits_is_unique : _GEN_128 ? _slots_39_io_out_uop_is_unique : _GEN_127 ? _slots_38_io_out_uop_is_unique : _slots_37_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_129 ? io_dis_uops_0_bits_flush_on_commit : _GEN_128 ? _slots_39_io_out_uop_flush_on_commit : _GEN_127 ? _slots_38_io_out_uop_flush_on_commit : _slots_37_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_129 ? io_dis_uops_0_bits_ldst_is_rs1 : _GEN_128 ? _slots_39_io_out_uop_ldst_is_rs1 : _GEN_127 ? _slots_38_io_out_uop_ldst_is_rs1 : _slots_37_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_129 ? io_dis_uops_0_bits_ldst : _GEN_128 ? _slots_39_io_out_uop_ldst : _GEN_127 ? _slots_38_io_out_uop_ldst : _slots_37_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_129 ? io_dis_uops_0_bits_lrs1 : _GEN_128 ? _slots_39_io_out_uop_lrs1 : _GEN_127 ? _slots_38_io_out_uop_lrs1 : _slots_37_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_129 ? io_dis_uops_0_bits_lrs2 : _GEN_128 ? _slots_39_io_out_uop_lrs2 : _GEN_127 ? _slots_38_io_out_uop_lrs2 : _slots_37_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_129 ? io_dis_uops_0_bits_lrs3 : _GEN_128 ? _slots_39_io_out_uop_lrs3 : _GEN_127 ? _slots_38_io_out_uop_lrs3 : _slots_37_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_129 ? io_dis_uops_0_bits_ldst_val : _GEN_128 ? _slots_39_io_out_uop_ldst_val : _GEN_127 ? _slots_38_io_out_uop_ldst_val : _slots_37_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_129 ? io_dis_uops_0_bits_dst_rtype : _GEN_128 ? _slots_39_io_out_uop_dst_rtype : _GEN_127 ? _slots_38_io_out_uop_dst_rtype : _slots_37_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_129 ? io_dis_uops_0_bits_lrs1_rtype : _GEN_128 ? _slots_39_io_out_uop_lrs1_rtype : _GEN_127 ? _slots_38_io_out_uop_lrs1_rtype : _slots_37_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_129 ? _GEN_3 : _GEN_128 ? _slots_39_io_out_uop_lrs2_rtype : _GEN_127 ? _slots_38_io_out_uop_lrs2_rtype : _slots_37_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_129 ? io_dis_uops_0_bits_frs3_en : _GEN_128 ? _slots_39_io_out_uop_frs3_en : _GEN_127 ? _slots_38_io_out_uop_frs3_en : _slots_37_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_129 ? io_dis_uops_0_bits_fp_val : _GEN_128 ? _slots_39_io_out_uop_fp_val : _GEN_127 ? _slots_38_io_out_uop_fp_val : _slots_37_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_129 ? io_dis_uops_0_bits_fp_single : _GEN_128 ? _slots_39_io_out_uop_fp_single : _GEN_127 ? _slots_38_io_out_uop_fp_single : _slots_37_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_129 ? io_dis_uops_0_bits_xcpt_pf_if : _GEN_128 ? _slots_39_io_out_uop_xcpt_pf_if : _GEN_127 ? _slots_38_io_out_uop_xcpt_pf_if : _slots_37_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_129 ? io_dis_uops_0_bits_xcpt_ae_if : _GEN_128 ? _slots_39_io_out_uop_xcpt_ae_if : _GEN_127 ? _slots_38_io_out_uop_xcpt_ae_if : _slots_37_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_129 ? io_dis_uops_0_bits_xcpt_ma_if : _GEN_128 ? _slots_39_io_out_uop_xcpt_ma_if : _GEN_127 ? _slots_38_io_out_uop_xcpt_ma_if : _slots_37_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_129 ? io_dis_uops_0_bits_bp_debug_if : _GEN_128 ? _slots_39_io_out_uop_bp_debug_if : _GEN_127 ? _slots_38_io_out_uop_bp_debug_if : _slots_37_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_129 ? io_dis_uops_0_bits_bp_xcpt_if : _GEN_128 ? _slots_39_io_out_uop_bp_xcpt_if : _GEN_127 ? _slots_38_io_out_uop_bp_xcpt_if : _slots_37_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_129 ? io_dis_uops_0_bits_debug_fsrc : _GEN_128 ? _slots_39_io_out_uop_debug_fsrc : _GEN_127 ? _slots_38_io_out_uop_debug_fsrc : _slots_37_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_129 ? io_dis_uops_0_bits_debug_tsrc : _GEN_128 ? _slots_39_io_out_uop_debug_tsrc : _GEN_127 ? _slots_38_io_out_uop_debug_tsrc : _slots_37_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_36_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_36_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_36_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_36_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_36_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_36_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_36_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_36_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_36_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_36_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_36_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_36_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_36_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_36_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_36_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_36_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_36_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_36_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_36_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_36_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_36_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_36_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_36_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_36_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_36_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_36_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_36_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_36_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_36_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_36_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_36_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_36_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_36_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_36_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_36_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_36_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_36_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_36_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_36_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_36_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_36_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_36_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_36_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_36_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_36_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_36_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_36_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_36_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_36_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_36_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_36_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_36_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_36_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_36_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_36_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_36_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_36_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_36_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_36_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_36_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_36_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_36_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_36_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_36_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_36_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_36_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_36_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_36_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_36_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_36_io_uop_uopc),
    .io_uop_inst                    (_slots_36_io_uop_inst),
    .io_uop_debug_inst              (_slots_36_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_36_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_36_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_36_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_36_io_uop_fu_code),
    .io_uop_iw_state                (_slots_36_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_36_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_36_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_36_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_36_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_36_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_36_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_36_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_36_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_36_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_36_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_36_io_uop_pc_lob),
    .io_uop_taken                   (_slots_36_io_uop_taken),
    .io_uop_imm_packed              (_slots_36_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_36_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_36_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_36_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_36_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_36_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_36_io_uop_pdst),
    .io_uop_prs1                    (_slots_36_io_uop_prs1),
    .io_uop_prs2                    (_slots_36_io_uop_prs2),
    .io_uop_prs3                    (_slots_36_io_uop_prs3),
    .io_uop_ppred                   (_slots_36_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_36_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_36_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_36_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_36_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_36_io_uop_stale_pdst),
    .io_uop_exception               (_slots_36_io_uop_exception),
    .io_uop_exc_cause               (_slots_36_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_36_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_36_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_36_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_36_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_36_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_36_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_36_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_36_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_36_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_36_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_36_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_36_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_36_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_36_io_uop_ldst),
    .io_uop_lrs1                    (_slots_36_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_36_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_36_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_36_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_36_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_36_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_36_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_36_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_36_io_uop_fp_val),
    .io_uop_fp_single               (_slots_36_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_36_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_36_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_36_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_36_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_36_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_36_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_36_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_37 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_37_io_valid),
    .io_will_be_valid               (_slots_37_io_will_be_valid),
    .io_request                     (_slots_37_io_request),
    .io_grant                       (issue_slots_37_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_36),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_37_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_132 ? io_dis_uops_1_bits_uopc : _GEN_131 ? io_dis_uops_0_bits_uopc : _GEN_130 ? _slots_39_io_out_uop_uopc : _slots_38_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_132 ? io_dis_uops_1_bits_inst : _GEN_131 ? io_dis_uops_0_bits_inst : _GEN_130 ? _slots_39_io_out_uop_inst : _slots_38_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_132 ? io_dis_uops_1_bits_debug_inst : _GEN_131 ? io_dis_uops_0_bits_debug_inst : _GEN_130 ? _slots_39_io_out_uop_debug_inst : _slots_38_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_132 ? io_dis_uops_1_bits_is_rvc : _GEN_131 ? io_dis_uops_0_bits_is_rvc : _GEN_130 ? _slots_39_io_out_uop_is_rvc : _slots_38_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_132 ? io_dis_uops_1_bits_debug_pc : _GEN_131 ? io_dis_uops_0_bits_debug_pc : _GEN_130 ? _slots_39_io_out_uop_debug_pc : _slots_38_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_132 ? io_dis_uops_1_bits_iq_type : _GEN_131 ? io_dis_uops_0_bits_iq_type : _GEN_130 ? _slots_39_io_out_uop_iq_type : _slots_38_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_132 ? io_dis_uops_1_bits_fu_code : _GEN_131 ? io_dis_uops_0_bits_fu_code : _GEN_130 ? _slots_39_io_out_uop_fu_code : _slots_38_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_132 ? _GEN_7 : _GEN_131 ? _GEN_1 : _GEN_130 ? _slots_39_io_out_uop_iw_state : _slots_38_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_133 & (_GEN_130 ? _slots_39_io_out_uop_iw_p1_poisoned : _slots_38_io_out_uop_iw_p1_poisoned)),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_133 & (_GEN_130 ? _slots_39_io_out_uop_iw_p2_poisoned : _slots_38_io_out_uop_iw_p2_poisoned)),
    .io_in_uop_bits_is_br           (_GEN_132 ? io_dis_uops_1_bits_is_br : _GEN_131 ? io_dis_uops_0_bits_is_br : _GEN_130 ? _slots_39_io_out_uop_is_br : _slots_38_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_132 ? io_dis_uops_1_bits_is_jalr : _GEN_131 ? io_dis_uops_0_bits_is_jalr : _GEN_130 ? _slots_39_io_out_uop_is_jalr : _slots_38_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_132 ? io_dis_uops_1_bits_is_jal : _GEN_131 ? io_dis_uops_0_bits_is_jal : _GEN_130 ? _slots_39_io_out_uop_is_jal : _slots_38_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_132 ? io_dis_uops_1_bits_is_sfb : _GEN_131 ? io_dis_uops_0_bits_is_sfb : _GEN_130 ? _slots_39_io_out_uop_is_sfb : _slots_38_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_132 ? io_dis_uops_1_bits_br_mask : _GEN_131 ? io_dis_uops_0_bits_br_mask : _GEN_130 ? _slots_39_io_out_uop_br_mask : _slots_38_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_132 ? io_dis_uops_1_bits_br_tag : _GEN_131 ? io_dis_uops_0_bits_br_tag : _GEN_130 ? _slots_39_io_out_uop_br_tag : _slots_38_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_132 ? io_dis_uops_1_bits_ftq_idx : _GEN_131 ? io_dis_uops_0_bits_ftq_idx : _GEN_130 ? _slots_39_io_out_uop_ftq_idx : _slots_38_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_132 ? io_dis_uops_1_bits_edge_inst : _GEN_131 ? io_dis_uops_0_bits_edge_inst : _GEN_130 ? _slots_39_io_out_uop_edge_inst : _slots_38_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_132 ? io_dis_uops_1_bits_pc_lob : _GEN_131 ? io_dis_uops_0_bits_pc_lob : _GEN_130 ? _slots_39_io_out_uop_pc_lob : _slots_38_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_132 ? io_dis_uops_1_bits_taken : _GEN_131 ? io_dis_uops_0_bits_taken : _GEN_130 ? _slots_39_io_out_uop_taken : _slots_38_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_132 ? io_dis_uops_1_bits_imm_packed : _GEN_131 ? io_dis_uops_0_bits_imm_packed : _GEN_130 ? _slots_39_io_out_uop_imm_packed : _slots_38_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_132 ? io_dis_uops_1_bits_csr_addr : _GEN_131 ? io_dis_uops_0_bits_csr_addr : _GEN_130 ? _slots_39_io_out_uop_csr_addr : _slots_38_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_132 ? io_dis_uops_1_bits_rob_idx : _GEN_131 ? io_dis_uops_0_bits_rob_idx : _GEN_130 ? _slots_39_io_out_uop_rob_idx : _slots_38_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_132 ? io_dis_uops_1_bits_ldq_idx : _GEN_131 ? io_dis_uops_0_bits_ldq_idx : _GEN_130 ? _slots_39_io_out_uop_ldq_idx : _slots_38_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_132 ? io_dis_uops_1_bits_stq_idx : _GEN_131 ? io_dis_uops_0_bits_stq_idx : _GEN_130 ? _slots_39_io_out_uop_stq_idx : _slots_38_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_132 ? io_dis_uops_1_bits_rxq_idx : _GEN_131 ? io_dis_uops_0_bits_rxq_idx : _GEN_130 ? _slots_39_io_out_uop_rxq_idx : _slots_38_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_132 ? io_dis_uops_1_bits_pdst : _GEN_131 ? io_dis_uops_0_bits_pdst : _GEN_130 ? _slots_39_io_out_uop_pdst : _slots_38_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_132 ? io_dis_uops_1_bits_prs1 : _GEN_131 ? io_dis_uops_0_bits_prs1 : _GEN_130 ? _slots_39_io_out_uop_prs1 : _slots_38_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_132 ? io_dis_uops_1_bits_prs2 : _GEN_131 ? io_dis_uops_0_bits_prs2 : _GEN_130 ? _slots_39_io_out_uop_prs2 : _slots_38_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_132 ? io_dis_uops_1_bits_prs3 : _GEN_131 ? io_dis_uops_0_bits_prs3 : _GEN_130 ? _slots_39_io_out_uop_prs3 : _slots_38_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_133 ? 6'h0 : _GEN_130 ? _slots_39_io_out_uop_ppred : _slots_38_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_132 ? io_dis_uops_1_bits_prs1_busy : _GEN_131 ? io_dis_uops_0_bits_prs1_busy : _GEN_130 ? _slots_39_io_out_uop_prs1_busy : _slots_38_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_132 ? _GEN_10 : _GEN_131 ? _GEN_4 : _GEN_130 ? _slots_39_io_out_uop_prs2_busy : _slots_38_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_133 & (_GEN_130 ? _slots_39_io_out_uop_prs3_busy : _slots_38_io_out_uop_prs3_busy)),
    .io_in_uop_bits_ppred_busy      (~_GEN_133 & (_GEN_130 ? _slots_39_io_out_uop_ppred_busy : _slots_38_io_out_uop_ppred_busy)),
    .io_in_uop_bits_stale_pdst      (_GEN_132 ? io_dis_uops_1_bits_stale_pdst : _GEN_131 ? io_dis_uops_0_bits_stale_pdst : _GEN_130 ? _slots_39_io_out_uop_stale_pdst : _slots_38_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_132 ? io_dis_uops_1_bits_exception : _GEN_131 ? io_dis_uops_0_bits_exception : _GEN_130 ? _slots_39_io_out_uop_exception : _slots_38_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_132 ? io_dis_uops_1_bits_exc_cause : _GEN_131 ? io_dis_uops_0_bits_exc_cause : _GEN_130 ? _slots_39_io_out_uop_exc_cause : _slots_38_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_132 ? io_dis_uops_1_bits_bypassable : _GEN_131 ? io_dis_uops_0_bits_bypassable : _GEN_130 ? _slots_39_io_out_uop_bypassable : _slots_38_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_132 ? io_dis_uops_1_bits_mem_cmd : _GEN_131 ? io_dis_uops_0_bits_mem_cmd : _GEN_130 ? _slots_39_io_out_uop_mem_cmd : _slots_38_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_132 ? io_dis_uops_1_bits_mem_size : _GEN_131 ? io_dis_uops_0_bits_mem_size : _GEN_130 ? _slots_39_io_out_uop_mem_size : _slots_38_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_132 ? io_dis_uops_1_bits_mem_signed : _GEN_131 ? io_dis_uops_0_bits_mem_signed : _GEN_130 ? _slots_39_io_out_uop_mem_signed : _slots_38_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_132 ? io_dis_uops_1_bits_is_fence : _GEN_131 ? io_dis_uops_0_bits_is_fence : _GEN_130 ? _slots_39_io_out_uop_is_fence : _slots_38_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_132 ? io_dis_uops_1_bits_is_fencei : _GEN_131 ? io_dis_uops_0_bits_is_fencei : _GEN_130 ? _slots_39_io_out_uop_is_fencei : _slots_38_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_132 ? io_dis_uops_1_bits_is_amo : _GEN_131 ? io_dis_uops_0_bits_is_amo : _GEN_130 ? _slots_39_io_out_uop_is_amo : _slots_38_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_132 ? io_dis_uops_1_bits_uses_ldq : _GEN_131 ? io_dis_uops_0_bits_uses_ldq : _GEN_130 ? _slots_39_io_out_uop_uses_ldq : _slots_38_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_132 ? io_dis_uops_1_bits_uses_stq : _GEN_131 ? io_dis_uops_0_bits_uses_stq : _GEN_130 ? _slots_39_io_out_uop_uses_stq : _slots_38_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_132 ? io_dis_uops_1_bits_is_sys_pc2epc : _GEN_131 ? io_dis_uops_0_bits_is_sys_pc2epc : _GEN_130 ? _slots_39_io_out_uop_is_sys_pc2epc : _slots_38_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_132 ? io_dis_uops_1_bits_is_unique : _GEN_131 ? io_dis_uops_0_bits_is_unique : _GEN_130 ? _slots_39_io_out_uop_is_unique : _slots_38_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_132 ? io_dis_uops_1_bits_flush_on_commit : _GEN_131 ? io_dis_uops_0_bits_flush_on_commit : _GEN_130 ? _slots_39_io_out_uop_flush_on_commit : _slots_38_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_132 ? io_dis_uops_1_bits_ldst_is_rs1 : _GEN_131 ? io_dis_uops_0_bits_ldst_is_rs1 : _GEN_130 ? _slots_39_io_out_uop_ldst_is_rs1 : _slots_38_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_132 ? io_dis_uops_1_bits_ldst : _GEN_131 ? io_dis_uops_0_bits_ldst : _GEN_130 ? _slots_39_io_out_uop_ldst : _slots_38_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_132 ? io_dis_uops_1_bits_lrs1 : _GEN_131 ? io_dis_uops_0_bits_lrs1 : _GEN_130 ? _slots_39_io_out_uop_lrs1 : _slots_38_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_132 ? io_dis_uops_1_bits_lrs2 : _GEN_131 ? io_dis_uops_0_bits_lrs2 : _GEN_130 ? _slots_39_io_out_uop_lrs2 : _slots_38_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_132 ? io_dis_uops_1_bits_lrs3 : _GEN_131 ? io_dis_uops_0_bits_lrs3 : _GEN_130 ? _slots_39_io_out_uop_lrs3 : _slots_38_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_132 ? io_dis_uops_1_bits_ldst_val : _GEN_131 ? io_dis_uops_0_bits_ldst_val : _GEN_130 ? _slots_39_io_out_uop_ldst_val : _slots_38_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_132 ? io_dis_uops_1_bits_dst_rtype : _GEN_131 ? io_dis_uops_0_bits_dst_rtype : _GEN_130 ? _slots_39_io_out_uop_dst_rtype : _slots_38_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_132 ? io_dis_uops_1_bits_lrs1_rtype : _GEN_131 ? io_dis_uops_0_bits_lrs1_rtype : _GEN_130 ? _slots_39_io_out_uop_lrs1_rtype : _slots_38_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_132 ? _GEN_9 : _GEN_131 ? _GEN_3 : _GEN_130 ? _slots_39_io_out_uop_lrs2_rtype : _slots_38_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_132 ? io_dis_uops_1_bits_frs3_en : _GEN_131 ? io_dis_uops_0_bits_frs3_en : _GEN_130 ? _slots_39_io_out_uop_frs3_en : _slots_38_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_132 ? io_dis_uops_1_bits_fp_val : _GEN_131 ? io_dis_uops_0_bits_fp_val : _GEN_130 ? _slots_39_io_out_uop_fp_val : _slots_38_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_132 ? io_dis_uops_1_bits_fp_single : _GEN_131 ? io_dis_uops_0_bits_fp_single : _GEN_130 ? _slots_39_io_out_uop_fp_single : _slots_38_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_132 ? io_dis_uops_1_bits_xcpt_pf_if : _GEN_131 ? io_dis_uops_0_bits_xcpt_pf_if : _GEN_130 ? _slots_39_io_out_uop_xcpt_pf_if : _slots_38_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_132 ? io_dis_uops_1_bits_xcpt_ae_if : _GEN_131 ? io_dis_uops_0_bits_xcpt_ae_if : _GEN_130 ? _slots_39_io_out_uop_xcpt_ae_if : _slots_38_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_132 ? io_dis_uops_1_bits_xcpt_ma_if : _GEN_131 ? io_dis_uops_0_bits_xcpt_ma_if : _GEN_130 ? _slots_39_io_out_uop_xcpt_ma_if : _slots_38_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_132 ? io_dis_uops_1_bits_bp_debug_if : _GEN_131 ? io_dis_uops_0_bits_bp_debug_if : _GEN_130 ? _slots_39_io_out_uop_bp_debug_if : _slots_38_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_132 ? io_dis_uops_1_bits_bp_xcpt_if : _GEN_131 ? io_dis_uops_0_bits_bp_xcpt_if : _GEN_130 ? _slots_39_io_out_uop_bp_xcpt_if : _slots_38_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_132 ? io_dis_uops_1_bits_debug_fsrc : _GEN_131 ? io_dis_uops_0_bits_debug_fsrc : _GEN_130 ? _slots_39_io_out_uop_debug_fsrc : _slots_38_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_132 ? io_dis_uops_1_bits_debug_tsrc : _GEN_131 ? io_dis_uops_0_bits_debug_tsrc : _GEN_130 ? _slots_39_io_out_uop_debug_tsrc : _slots_38_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_37_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_37_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_37_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_37_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_37_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_37_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_37_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_37_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_37_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_37_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_37_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_37_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_37_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_37_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_37_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_37_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_37_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_37_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_37_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_37_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_37_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_37_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_37_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_37_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_37_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_37_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_37_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_37_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_37_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_37_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_37_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_37_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_37_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_37_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_37_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_37_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_37_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_37_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_37_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_37_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_37_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_37_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_37_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_37_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_37_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_37_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_37_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_37_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_37_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_37_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_37_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_37_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_37_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_37_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_37_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_37_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_37_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_37_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_37_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_37_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_37_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_37_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_37_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_37_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_37_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_37_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_37_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_37_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_37_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_37_io_uop_uopc),
    .io_uop_inst                    (_slots_37_io_uop_inst),
    .io_uop_debug_inst              (_slots_37_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_37_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_37_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_37_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_37_io_uop_fu_code),
    .io_uop_iw_state                (_slots_37_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_37_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_37_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_37_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_37_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_37_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_37_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_37_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_37_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_37_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_37_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_37_io_uop_pc_lob),
    .io_uop_taken                   (_slots_37_io_uop_taken),
    .io_uop_imm_packed              (_slots_37_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_37_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_37_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_37_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_37_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_37_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_37_io_uop_pdst),
    .io_uop_prs1                    (_slots_37_io_uop_prs1),
    .io_uop_prs2                    (_slots_37_io_uop_prs2),
    .io_uop_prs3                    (_slots_37_io_uop_prs3),
    .io_uop_ppred                   (_slots_37_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_37_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_37_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_37_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_37_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_37_io_uop_stale_pdst),
    .io_uop_exception               (_slots_37_io_uop_exception),
    .io_uop_exc_cause               (_slots_37_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_37_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_37_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_37_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_37_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_37_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_37_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_37_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_37_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_37_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_37_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_37_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_37_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_37_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_37_io_uop_ldst),
    .io_uop_lrs1                    (_slots_37_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_37_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_37_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_37_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_37_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_37_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_37_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_37_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_37_io_uop_fp_val),
    .io_uop_fp_single               (_slots_37_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_37_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_37_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_37_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_37_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_37_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_37_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_37_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_38 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_38_io_valid),
    .io_will_be_valid               (_slots_38_io_will_be_valid),
    .io_request                     (_slots_38_io_request),
    .io_grant                       (issue_slots_38_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_37),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_38_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_136 ? io_dis_uops_2_bits_uopc : _GEN_135 ? io_dis_uops_1_bits_uopc : _GEN_134 ? io_dis_uops_0_bits_uopc : _slots_39_io_out_uop_uopc),
    .io_in_uop_bits_inst            (_GEN_136 ? io_dis_uops_2_bits_inst : _GEN_135 ? io_dis_uops_1_bits_inst : _GEN_134 ? io_dis_uops_0_bits_inst : _slots_39_io_out_uop_inst),
    .io_in_uop_bits_debug_inst      (_GEN_136 ? io_dis_uops_2_bits_debug_inst : _GEN_135 ? io_dis_uops_1_bits_debug_inst : _GEN_134 ? io_dis_uops_0_bits_debug_inst : _slots_39_io_out_uop_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_136 ? io_dis_uops_2_bits_is_rvc : _GEN_135 ? io_dis_uops_1_bits_is_rvc : _GEN_134 ? io_dis_uops_0_bits_is_rvc : _slots_39_io_out_uop_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_136 ? io_dis_uops_2_bits_debug_pc : _GEN_135 ? io_dis_uops_1_bits_debug_pc : _GEN_134 ? io_dis_uops_0_bits_debug_pc : _slots_39_io_out_uop_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_136 ? io_dis_uops_2_bits_iq_type : _GEN_135 ? io_dis_uops_1_bits_iq_type : _GEN_134 ? io_dis_uops_0_bits_iq_type : _slots_39_io_out_uop_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_136 ? io_dis_uops_2_bits_fu_code : _GEN_135 ? io_dis_uops_1_bits_fu_code : _GEN_134 ? io_dis_uops_0_bits_fu_code : _slots_39_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_136 ? (_GEN_12 ? 2'h2 : 2'h1) : _GEN_135 ? _GEN_7 : _GEN_134 ? _GEN_1 : _slots_39_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_137 & _slots_39_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_137 & _slots_39_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_136 ? io_dis_uops_2_bits_is_br : _GEN_135 ? io_dis_uops_1_bits_is_br : _GEN_134 ? io_dis_uops_0_bits_is_br : _slots_39_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_136 ? io_dis_uops_2_bits_is_jalr : _GEN_135 ? io_dis_uops_1_bits_is_jalr : _GEN_134 ? io_dis_uops_0_bits_is_jalr : _slots_39_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_136 ? io_dis_uops_2_bits_is_jal : _GEN_135 ? io_dis_uops_1_bits_is_jal : _GEN_134 ? io_dis_uops_0_bits_is_jal : _slots_39_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_136 ? io_dis_uops_2_bits_is_sfb : _GEN_135 ? io_dis_uops_1_bits_is_sfb : _GEN_134 ? io_dis_uops_0_bits_is_sfb : _slots_39_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_136 ? io_dis_uops_2_bits_br_mask : _GEN_135 ? io_dis_uops_1_bits_br_mask : _GEN_134 ? io_dis_uops_0_bits_br_mask : _slots_39_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_136 ? io_dis_uops_2_bits_br_tag : _GEN_135 ? io_dis_uops_1_bits_br_tag : _GEN_134 ? io_dis_uops_0_bits_br_tag : _slots_39_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_136 ? io_dis_uops_2_bits_ftq_idx : _GEN_135 ? io_dis_uops_1_bits_ftq_idx : _GEN_134 ? io_dis_uops_0_bits_ftq_idx : _slots_39_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_136 ? io_dis_uops_2_bits_edge_inst : _GEN_135 ? io_dis_uops_1_bits_edge_inst : _GEN_134 ? io_dis_uops_0_bits_edge_inst : _slots_39_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_136 ? io_dis_uops_2_bits_pc_lob : _GEN_135 ? io_dis_uops_1_bits_pc_lob : _GEN_134 ? io_dis_uops_0_bits_pc_lob : _slots_39_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_136 ? io_dis_uops_2_bits_taken : _GEN_135 ? io_dis_uops_1_bits_taken : _GEN_134 ? io_dis_uops_0_bits_taken : _slots_39_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_136 ? io_dis_uops_2_bits_imm_packed : _GEN_135 ? io_dis_uops_1_bits_imm_packed : _GEN_134 ? io_dis_uops_0_bits_imm_packed : _slots_39_io_out_uop_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_136 ? io_dis_uops_2_bits_csr_addr : _GEN_135 ? io_dis_uops_1_bits_csr_addr : _GEN_134 ? io_dis_uops_0_bits_csr_addr : _slots_39_io_out_uop_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_136 ? io_dis_uops_2_bits_rob_idx : _GEN_135 ? io_dis_uops_1_bits_rob_idx : _GEN_134 ? io_dis_uops_0_bits_rob_idx : _slots_39_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_136 ? io_dis_uops_2_bits_ldq_idx : _GEN_135 ? io_dis_uops_1_bits_ldq_idx : _GEN_134 ? io_dis_uops_0_bits_ldq_idx : _slots_39_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_136 ? io_dis_uops_2_bits_stq_idx : _GEN_135 ? io_dis_uops_1_bits_stq_idx : _GEN_134 ? io_dis_uops_0_bits_stq_idx : _slots_39_io_out_uop_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_136 ? io_dis_uops_2_bits_rxq_idx : _GEN_135 ? io_dis_uops_1_bits_rxq_idx : _GEN_134 ? io_dis_uops_0_bits_rxq_idx : _slots_39_io_out_uop_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_136 ? io_dis_uops_2_bits_pdst : _GEN_135 ? io_dis_uops_1_bits_pdst : _GEN_134 ? io_dis_uops_0_bits_pdst : _slots_39_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_136 ? io_dis_uops_2_bits_prs1 : _GEN_135 ? io_dis_uops_1_bits_prs1 : _GEN_134 ? io_dis_uops_0_bits_prs1 : _slots_39_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_136 ? io_dis_uops_2_bits_prs2 : _GEN_135 ? io_dis_uops_1_bits_prs2 : _GEN_134 ? io_dis_uops_0_bits_prs2 : _slots_39_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_136 ? io_dis_uops_2_bits_prs3 : _GEN_135 ? io_dis_uops_1_bits_prs3 : _GEN_134 ? io_dis_uops_0_bits_prs3 : _slots_39_io_out_uop_prs3),
    .io_in_uop_bits_ppred           (_GEN_137 ? 6'h0 : _slots_39_io_out_uop_ppred),
    .io_in_uop_bits_prs1_busy       (_GEN_136 ? io_dis_uops_2_bits_prs1_busy : _GEN_135 ? io_dis_uops_1_bits_prs1_busy : _GEN_134 ? io_dis_uops_0_bits_prs1_busy : _slots_39_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_136 ? _GEN_15 : _GEN_135 ? _GEN_10 : _GEN_134 ? _GEN_4 : _slots_39_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_137 & _slots_39_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (~_GEN_137 & _slots_39_io_out_uop_ppred_busy),
    .io_in_uop_bits_stale_pdst      (_GEN_136 ? io_dis_uops_2_bits_stale_pdst : _GEN_135 ? io_dis_uops_1_bits_stale_pdst : _GEN_134 ? io_dis_uops_0_bits_stale_pdst : _slots_39_io_out_uop_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_136 ? io_dis_uops_2_bits_exception : _GEN_135 ? io_dis_uops_1_bits_exception : _GEN_134 ? io_dis_uops_0_bits_exception : _slots_39_io_out_uop_exception),
    .io_in_uop_bits_exc_cause       (_GEN_136 ? io_dis_uops_2_bits_exc_cause : _GEN_135 ? io_dis_uops_1_bits_exc_cause : _GEN_134 ? io_dis_uops_0_bits_exc_cause : _slots_39_io_out_uop_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_136 ? io_dis_uops_2_bits_bypassable : _GEN_135 ? io_dis_uops_1_bits_bypassable : _GEN_134 ? io_dis_uops_0_bits_bypassable : _slots_39_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_136 ? io_dis_uops_2_bits_mem_cmd : _GEN_135 ? io_dis_uops_1_bits_mem_cmd : _GEN_134 ? io_dis_uops_0_bits_mem_cmd : _slots_39_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_136 ? io_dis_uops_2_bits_mem_size : _GEN_135 ? io_dis_uops_1_bits_mem_size : _GEN_134 ? io_dis_uops_0_bits_mem_size : _slots_39_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_136 ? io_dis_uops_2_bits_mem_signed : _GEN_135 ? io_dis_uops_1_bits_mem_signed : _GEN_134 ? io_dis_uops_0_bits_mem_signed : _slots_39_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_136 ? io_dis_uops_2_bits_is_fence : _GEN_135 ? io_dis_uops_1_bits_is_fence : _GEN_134 ? io_dis_uops_0_bits_is_fence : _slots_39_io_out_uop_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_136 ? io_dis_uops_2_bits_is_fencei : _GEN_135 ? io_dis_uops_1_bits_is_fencei : _GEN_134 ? io_dis_uops_0_bits_is_fencei : _slots_39_io_out_uop_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_136 ? io_dis_uops_2_bits_is_amo : _GEN_135 ? io_dis_uops_1_bits_is_amo : _GEN_134 ? io_dis_uops_0_bits_is_amo : _slots_39_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_136 ? io_dis_uops_2_bits_uses_ldq : _GEN_135 ? io_dis_uops_1_bits_uses_ldq : _GEN_134 ? io_dis_uops_0_bits_uses_ldq : _slots_39_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_136 ? io_dis_uops_2_bits_uses_stq : _GEN_135 ? io_dis_uops_1_bits_uses_stq : _GEN_134 ? io_dis_uops_0_bits_uses_stq : _slots_39_io_out_uop_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_136 ? io_dis_uops_2_bits_is_sys_pc2epc : _GEN_135 ? io_dis_uops_1_bits_is_sys_pc2epc : _GEN_134 ? io_dis_uops_0_bits_is_sys_pc2epc : _slots_39_io_out_uop_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_136 ? io_dis_uops_2_bits_is_unique : _GEN_135 ? io_dis_uops_1_bits_is_unique : _GEN_134 ? io_dis_uops_0_bits_is_unique : _slots_39_io_out_uop_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_136 ? io_dis_uops_2_bits_flush_on_commit : _GEN_135 ? io_dis_uops_1_bits_flush_on_commit : _GEN_134 ? io_dis_uops_0_bits_flush_on_commit : _slots_39_io_out_uop_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_136 ? io_dis_uops_2_bits_ldst_is_rs1 : _GEN_135 ? io_dis_uops_1_bits_ldst_is_rs1 : _GEN_134 ? io_dis_uops_0_bits_ldst_is_rs1 : _slots_39_io_out_uop_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_136 ? io_dis_uops_2_bits_ldst : _GEN_135 ? io_dis_uops_1_bits_ldst : _GEN_134 ? io_dis_uops_0_bits_ldst : _slots_39_io_out_uop_ldst),
    .io_in_uop_bits_lrs1            (_GEN_136 ? io_dis_uops_2_bits_lrs1 : _GEN_135 ? io_dis_uops_1_bits_lrs1 : _GEN_134 ? io_dis_uops_0_bits_lrs1 : _slots_39_io_out_uop_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_136 ? io_dis_uops_2_bits_lrs2 : _GEN_135 ? io_dis_uops_1_bits_lrs2 : _GEN_134 ? io_dis_uops_0_bits_lrs2 : _slots_39_io_out_uop_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_136 ? io_dis_uops_2_bits_lrs3 : _GEN_135 ? io_dis_uops_1_bits_lrs3 : _GEN_134 ? io_dis_uops_0_bits_lrs3 : _slots_39_io_out_uop_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_136 ? io_dis_uops_2_bits_ldst_val : _GEN_135 ? io_dis_uops_1_bits_ldst_val : _GEN_134 ? io_dis_uops_0_bits_ldst_val : _slots_39_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_136 ? io_dis_uops_2_bits_dst_rtype : _GEN_135 ? io_dis_uops_1_bits_dst_rtype : _GEN_134 ? io_dis_uops_0_bits_dst_rtype : _slots_39_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_136 ? io_dis_uops_2_bits_lrs1_rtype : _GEN_135 ? io_dis_uops_1_bits_lrs1_rtype : _GEN_134 ? io_dis_uops_0_bits_lrs1_rtype : _slots_39_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_136 ? _GEN_14 : _GEN_135 ? _GEN_9 : _GEN_134 ? _GEN_3 : _slots_39_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_frs3_en         (_GEN_136 ? io_dis_uops_2_bits_frs3_en : _GEN_135 ? io_dis_uops_1_bits_frs3_en : _GEN_134 ? io_dis_uops_0_bits_frs3_en : _slots_39_io_out_uop_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_136 ? io_dis_uops_2_bits_fp_val : _GEN_135 ? io_dis_uops_1_bits_fp_val : _GEN_134 ? io_dis_uops_0_bits_fp_val : _slots_39_io_out_uop_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_136 ? io_dis_uops_2_bits_fp_single : _GEN_135 ? io_dis_uops_1_bits_fp_single : _GEN_134 ? io_dis_uops_0_bits_fp_single : _slots_39_io_out_uop_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_136 ? io_dis_uops_2_bits_xcpt_pf_if : _GEN_135 ? io_dis_uops_1_bits_xcpt_pf_if : _GEN_134 ? io_dis_uops_0_bits_xcpt_pf_if : _slots_39_io_out_uop_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_136 ? io_dis_uops_2_bits_xcpt_ae_if : _GEN_135 ? io_dis_uops_1_bits_xcpt_ae_if : _GEN_134 ? io_dis_uops_0_bits_xcpt_ae_if : _slots_39_io_out_uop_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_136 ? io_dis_uops_2_bits_xcpt_ma_if : _GEN_135 ? io_dis_uops_1_bits_xcpt_ma_if : _GEN_134 ? io_dis_uops_0_bits_xcpt_ma_if : _slots_39_io_out_uop_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_136 ? io_dis_uops_2_bits_bp_debug_if : _GEN_135 ? io_dis_uops_1_bits_bp_debug_if : _GEN_134 ? io_dis_uops_0_bits_bp_debug_if : _slots_39_io_out_uop_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_136 ? io_dis_uops_2_bits_bp_xcpt_if : _GEN_135 ? io_dis_uops_1_bits_bp_xcpt_if : _GEN_134 ? io_dis_uops_0_bits_bp_xcpt_if : _slots_39_io_out_uop_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_136 ? io_dis_uops_2_bits_debug_fsrc : _GEN_135 ? io_dis_uops_1_bits_debug_fsrc : _GEN_134 ? io_dis_uops_0_bits_debug_fsrc : _slots_39_io_out_uop_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_136 ? io_dis_uops_2_bits_debug_tsrc : _GEN_135 ? io_dis_uops_1_bits_debug_tsrc : _GEN_134 ? io_dis_uops_0_bits_debug_tsrc : _slots_39_io_out_uop_debug_tsrc),
    .io_out_uop_uopc                (_slots_38_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_38_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_38_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_38_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_38_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_38_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_38_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_38_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_38_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_38_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_38_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_38_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_38_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_38_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_38_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_38_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_38_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_38_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_38_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_38_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_38_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_38_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_38_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_38_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_38_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_38_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_38_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_38_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_38_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_38_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_38_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_38_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_38_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_38_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_38_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_38_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_38_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_38_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_38_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_38_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_38_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_38_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_38_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_38_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_38_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_38_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_38_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_38_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_38_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_38_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_38_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_38_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_38_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_38_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_38_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_38_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_38_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_38_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_38_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_38_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_38_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_38_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_38_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_38_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_38_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_38_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_38_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_38_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_38_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_38_io_uop_uopc),
    .io_uop_inst                    (_slots_38_io_uop_inst),
    .io_uop_debug_inst              (_slots_38_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_38_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_38_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_38_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_38_io_uop_fu_code),
    .io_uop_iw_state                (_slots_38_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_38_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_38_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_38_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_38_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_38_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_38_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_38_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_38_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_38_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_38_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_38_io_uop_pc_lob),
    .io_uop_taken                   (_slots_38_io_uop_taken),
    .io_uop_imm_packed              (_slots_38_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_38_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_38_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_38_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_38_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_38_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_38_io_uop_pdst),
    .io_uop_prs1                    (_slots_38_io_uop_prs1),
    .io_uop_prs2                    (_slots_38_io_uop_prs2),
    .io_uop_prs3                    (_slots_38_io_uop_prs3),
    .io_uop_ppred                   (_slots_38_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_38_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_38_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_38_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_38_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_38_io_uop_stale_pdst),
    .io_uop_exception               (_slots_38_io_uop_exception),
    .io_uop_exc_cause               (_slots_38_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_38_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_38_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_38_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_38_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_38_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_38_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_38_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_38_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_38_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_38_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_38_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_38_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_38_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_38_io_uop_ldst),
    .io_uop_lrs1                    (_slots_38_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_38_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_38_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_38_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_38_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_38_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_38_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_38_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_38_io_uop_fp_val),
    .io_uop_fp_single               (_slots_38_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_38_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_38_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_38_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_38_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_38_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_38_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_38_io_uop_debug_tsrc)
  );
  IssueSlot_32 slots_39 (
    .clock                          (clock),
    .reset                          (reset),
    .io_valid                       (_slots_39_io_valid),
    .io_will_be_valid               (_slots_39_io_will_be_valid),
    .io_request                     (_slots_39_io_request),
    .io_grant                       (issue_slots_39_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|next_38),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_39_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_140 ? io_dis_uops_3_bits_uopc : _GEN_139 ? io_dis_uops_2_bits_uopc : _GEN_138 ? io_dis_uops_1_bits_uopc : io_dis_uops_0_bits_uopc),
    .io_in_uop_bits_inst            (_GEN_140 ? io_dis_uops_3_bits_inst : _GEN_139 ? io_dis_uops_2_bits_inst : _GEN_138 ? io_dis_uops_1_bits_inst : io_dis_uops_0_bits_inst),
    .io_in_uop_bits_debug_inst      (_GEN_140 ? io_dis_uops_3_bits_debug_inst : _GEN_139 ? io_dis_uops_2_bits_debug_inst : _GEN_138 ? io_dis_uops_1_bits_debug_inst : io_dis_uops_0_bits_debug_inst),
    .io_in_uop_bits_is_rvc          (_GEN_140 ? io_dis_uops_3_bits_is_rvc : _GEN_139 ? io_dis_uops_2_bits_is_rvc : _GEN_138 ? io_dis_uops_1_bits_is_rvc : io_dis_uops_0_bits_is_rvc),
    .io_in_uop_bits_debug_pc        (_GEN_140 ? io_dis_uops_3_bits_debug_pc : _GEN_139 ? io_dis_uops_2_bits_debug_pc : _GEN_138 ? io_dis_uops_1_bits_debug_pc : io_dis_uops_0_bits_debug_pc),
    .io_in_uop_bits_iq_type         (_GEN_140 ? io_dis_uops_3_bits_iq_type : _GEN_139 ? io_dis_uops_2_bits_iq_type : _GEN_138 ? io_dis_uops_1_bits_iq_type : io_dis_uops_0_bits_iq_type),
    .io_in_uop_bits_fu_code         (_GEN_140 ? io_dis_uops_3_bits_fu_code : _GEN_139 ? io_dis_uops_2_bits_fu_code : _GEN_138 ? io_dis_uops_1_bits_fu_code : io_dis_uops_0_bits_fu_code),
    .io_in_uop_bits_iw_state        ((_GEN_140 ? _GEN_17 : _GEN_139 ? _GEN_12 : _GEN_138 ? _GEN_6 : _GEN_0) ? 2'h2 : 2'h1),
    .io_in_uop_bits_iw_p1_poisoned  (1'h0),
    .io_in_uop_bits_iw_p2_poisoned  (1'h0),
    .io_in_uop_bits_is_br           (_GEN_140 ? io_dis_uops_3_bits_is_br : _GEN_139 ? io_dis_uops_2_bits_is_br : _GEN_138 ? io_dis_uops_1_bits_is_br : io_dis_uops_0_bits_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_140 ? io_dis_uops_3_bits_is_jalr : _GEN_139 ? io_dis_uops_2_bits_is_jalr : _GEN_138 ? io_dis_uops_1_bits_is_jalr : io_dis_uops_0_bits_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_140 ? io_dis_uops_3_bits_is_jal : _GEN_139 ? io_dis_uops_2_bits_is_jal : _GEN_138 ? io_dis_uops_1_bits_is_jal : io_dis_uops_0_bits_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_140 ? io_dis_uops_3_bits_is_sfb : _GEN_139 ? io_dis_uops_2_bits_is_sfb : _GEN_138 ? io_dis_uops_1_bits_is_sfb : io_dis_uops_0_bits_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_140 ? io_dis_uops_3_bits_br_mask : _GEN_139 ? io_dis_uops_2_bits_br_mask : _GEN_138 ? io_dis_uops_1_bits_br_mask : io_dis_uops_0_bits_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_140 ? io_dis_uops_3_bits_br_tag : _GEN_139 ? io_dis_uops_2_bits_br_tag : _GEN_138 ? io_dis_uops_1_bits_br_tag : io_dis_uops_0_bits_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_140 ? io_dis_uops_3_bits_ftq_idx : _GEN_139 ? io_dis_uops_2_bits_ftq_idx : _GEN_138 ? io_dis_uops_1_bits_ftq_idx : io_dis_uops_0_bits_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_140 ? io_dis_uops_3_bits_edge_inst : _GEN_139 ? io_dis_uops_2_bits_edge_inst : _GEN_138 ? io_dis_uops_1_bits_edge_inst : io_dis_uops_0_bits_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_140 ? io_dis_uops_3_bits_pc_lob : _GEN_139 ? io_dis_uops_2_bits_pc_lob : _GEN_138 ? io_dis_uops_1_bits_pc_lob : io_dis_uops_0_bits_pc_lob),
    .io_in_uop_bits_taken           (_GEN_140 ? io_dis_uops_3_bits_taken : _GEN_139 ? io_dis_uops_2_bits_taken : _GEN_138 ? io_dis_uops_1_bits_taken : io_dis_uops_0_bits_taken),
    .io_in_uop_bits_imm_packed      (_GEN_140 ? io_dis_uops_3_bits_imm_packed : _GEN_139 ? io_dis_uops_2_bits_imm_packed : _GEN_138 ? io_dis_uops_1_bits_imm_packed : io_dis_uops_0_bits_imm_packed),
    .io_in_uop_bits_csr_addr        (_GEN_140 ? io_dis_uops_3_bits_csr_addr : _GEN_139 ? io_dis_uops_2_bits_csr_addr : _GEN_138 ? io_dis_uops_1_bits_csr_addr : io_dis_uops_0_bits_csr_addr),
    .io_in_uop_bits_rob_idx         (_GEN_140 ? io_dis_uops_3_bits_rob_idx : _GEN_139 ? io_dis_uops_2_bits_rob_idx : _GEN_138 ? io_dis_uops_1_bits_rob_idx : io_dis_uops_0_bits_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_140 ? io_dis_uops_3_bits_ldq_idx : _GEN_139 ? io_dis_uops_2_bits_ldq_idx : _GEN_138 ? io_dis_uops_1_bits_ldq_idx : io_dis_uops_0_bits_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_140 ? io_dis_uops_3_bits_stq_idx : _GEN_139 ? io_dis_uops_2_bits_stq_idx : _GEN_138 ? io_dis_uops_1_bits_stq_idx : io_dis_uops_0_bits_stq_idx),
    .io_in_uop_bits_rxq_idx         (_GEN_140 ? io_dis_uops_3_bits_rxq_idx : _GEN_139 ? io_dis_uops_2_bits_rxq_idx : _GEN_138 ? io_dis_uops_1_bits_rxq_idx : io_dis_uops_0_bits_rxq_idx),
    .io_in_uop_bits_pdst            (_GEN_140 ? io_dis_uops_3_bits_pdst : _GEN_139 ? io_dis_uops_2_bits_pdst : _GEN_138 ? io_dis_uops_1_bits_pdst : io_dis_uops_0_bits_pdst),
    .io_in_uop_bits_prs1            (_GEN_140 ? io_dis_uops_3_bits_prs1 : _GEN_139 ? io_dis_uops_2_bits_prs1 : _GEN_138 ? io_dis_uops_1_bits_prs1 : io_dis_uops_0_bits_prs1),
    .io_in_uop_bits_prs2            (_GEN_140 ? io_dis_uops_3_bits_prs2 : _GEN_139 ? io_dis_uops_2_bits_prs2 : _GEN_138 ? io_dis_uops_1_bits_prs2 : io_dis_uops_0_bits_prs2),
    .io_in_uop_bits_prs3            (_GEN_140 ? io_dis_uops_3_bits_prs3 : _GEN_139 ? io_dis_uops_2_bits_prs3 : _GEN_138 ? io_dis_uops_1_bits_prs3 : io_dis_uops_0_bits_prs3),
    .io_in_uop_bits_ppred           (6'h0),
    .io_in_uop_bits_prs1_busy       (_GEN_140 ? io_dis_uops_3_bits_prs1_busy : _GEN_139 ? io_dis_uops_2_bits_prs1_busy : _GEN_138 ? io_dis_uops_1_bits_prs1_busy : io_dis_uops_0_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_140 ? _GEN_18 & io_dis_uops_3_bits_prs2_busy : _GEN_139 ? _GEN_15 : _GEN_138 ? _GEN_10 : _GEN_4),
    .io_in_uop_bits_prs3_busy       (1'h0),
    .io_in_uop_bits_ppred_busy      (1'h0),
    .io_in_uop_bits_stale_pdst      (_GEN_140 ? io_dis_uops_3_bits_stale_pdst : _GEN_139 ? io_dis_uops_2_bits_stale_pdst : _GEN_138 ? io_dis_uops_1_bits_stale_pdst : io_dis_uops_0_bits_stale_pdst),
    .io_in_uop_bits_exception       (_GEN_140 ? io_dis_uops_3_bits_exception : _GEN_139 ? io_dis_uops_2_bits_exception : _GEN_138 ? io_dis_uops_1_bits_exception : io_dis_uops_0_bits_exception),
    .io_in_uop_bits_exc_cause       (_GEN_140 ? io_dis_uops_3_bits_exc_cause : _GEN_139 ? io_dis_uops_2_bits_exc_cause : _GEN_138 ? io_dis_uops_1_bits_exc_cause : io_dis_uops_0_bits_exc_cause),
    .io_in_uop_bits_bypassable      (_GEN_140 ? io_dis_uops_3_bits_bypassable : _GEN_139 ? io_dis_uops_2_bits_bypassable : _GEN_138 ? io_dis_uops_1_bits_bypassable : io_dis_uops_0_bits_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_140 ? io_dis_uops_3_bits_mem_cmd : _GEN_139 ? io_dis_uops_2_bits_mem_cmd : _GEN_138 ? io_dis_uops_1_bits_mem_cmd : io_dis_uops_0_bits_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_140 ? io_dis_uops_3_bits_mem_size : _GEN_139 ? io_dis_uops_2_bits_mem_size : _GEN_138 ? io_dis_uops_1_bits_mem_size : io_dis_uops_0_bits_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_140 ? io_dis_uops_3_bits_mem_signed : _GEN_139 ? io_dis_uops_2_bits_mem_signed : _GEN_138 ? io_dis_uops_1_bits_mem_signed : io_dis_uops_0_bits_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_140 ? io_dis_uops_3_bits_is_fence : _GEN_139 ? io_dis_uops_2_bits_is_fence : _GEN_138 ? io_dis_uops_1_bits_is_fence : io_dis_uops_0_bits_is_fence),
    .io_in_uop_bits_is_fencei       (_GEN_140 ? io_dis_uops_3_bits_is_fencei : _GEN_139 ? io_dis_uops_2_bits_is_fencei : _GEN_138 ? io_dis_uops_1_bits_is_fencei : io_dis_uops_0_bits_is_fencei),
    .io_in_uop_bits_is_amo          (_GEN_140 ? io_dis_uops_3_bits_is_amo : _GEN_139 ? io_dis_uops_2_bits_is_amo : _GEN_138 ? io_dis_uops_1_bits_is_amo : io_dis_uops_0_bits_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_140 ? io_dis_uops_3_bits_uses_ldq : _GEN_139 ? io_dis_uops_2_bits_uses_ldq : _GEN_138 ? io_dis_uops_1_bits_uses_ldq : io_dis_uops_0_bits_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_140 ? io_dis_uops_3_bits_uses_stq : _GEN_139 ? io_dis_uops_2_bits_uses_stq : _GEN_138 ? io_dis_uops_1_bits_uses_stq : io_dis_uops_0_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc   (_GEN_140 ? io_dis_uops_3_bits_is_sys_pc2epc : _GEN_139 ? io_dis_uops_2_bits_is_sys_pc2epc : _GEN_138 ? io_dis_uops_1_bits_is_sys_pc2epc : io_dis_uops_0_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique       (_GEN_140 ? io_dis_uops_3_bits_is_unique : _GEN_139 ? io_dis_uops_2_bits_is_unique : _GEN_138 ? io_dis_uops_1_bits_is_unique : io_dis_uops_0_bits_is_unique),
    .io_in_uop_bits_flush_on_commit (_GEN_140 ? io_dis_uops_3_bits_flush_on_commit : _GEN_139 ? io_dis_uops_2_bits_flush_on_commit : _GEN_138 ? io_dis_uops_1_bits_flush_on_commit : io_dis_uops_0_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1     (_GEN_140 ? io_dis_uops_3_bits_ldst_is_rs1 : _GEN_139 ? io_dis_uops_2_bits_ldst_is_rs1 : _GEN_138 ? io_dis_uops_1_bits_ldst_is_rs1 : io_dis_uops_0_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst            (_GEN_140 ? io_dis_uops_3_bits_ldst : _GEN_139 ? io_dis_uops_2_bits_ldst : _GEN_138 ? io_dis_uops_1_bits_ldst : io_dis_uops_0_bits_ldst),
    .io_in_uop_bits_lrs1            (_GEN_140 ? io_dis_uops_3_bits_lrs1 : _GEN_139 ? io_dis_uops_2_bits_lrs1 : _GEN_138 ? io_dis_uops_1_bits_lrs1 : io_dis_uops_0_bits_lrs1),
    .io_in_uop_bits_lrs2            (_GEN_140 ? io_dis_uops_3_bits_lrs2 : _GEN_139 ? io_dis_uops_2_bits_lrs2 : _GEN_138 ? io_dis_uops_1_bits_lrs2 : io_dis_uops_0_bits_lrs2),
    .io_in_uop_bits_lrs3            (_GEN_140 ? io_dis_uops_3_bits_lrs3 : _GEN_139 ? io_dis_uops_2_bits_lrs3 : _GEN_138 ? io_dis_uops_1_bits_lrs3 : io_dis_uops_0_bits_lrs3),
    .io_in_uop_bits_ldst_val        (_GEN_140 ? io_dis_uops_3_bits_ldst_val : _GEN_139 ? io_dis_uops_2_bits_ldst_val : _GEN_138 ? io_dis_uops_1_bits_ldst_val : io_dis_uops_0_bits_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_140 ? io_dis_uops_3_bits_dst_rtype : _GEN_139 ? io_dis_uops_2_bits_dst_rtype : _GEN_138 ? io_dis_uops_1_bits_dst_rtype : io_dis_uops_0_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_140 ? io_dis_uops_3_bits_lrs1_rtype : _GEN_139 ? io_dis_uops_2_bits_lrs1_rtype : _GEN_138 ? io_dis_uops_1_bits_lrs1_rtype : io_dis_uops_0_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_140 ? (_GEN_18 ? io_dis_uops_3_bits_lrs2_rtype : 2'h2) : _GEN_139 ? _GEN_14 : _GEN_138 ? _GEN_9 : _GEN_3),
    .io_in_uop_bits_frs3_en         (_GEN_140 ? io_dis_uops_3_bits_frs3_en : _GEN_139 ? io_dis_uops_2_bits_frs3_en : _GEN_138 ? io_dis_uops_1_bits_frs3_en : io_dis_uops_0_bits_frs3_en),
    .io_in_uop_bits_fp_val          (_GEN_140 ? io_dis_uops_3_bits_fp_val : _GEN_139 ? io_dis_uops_2_bits_fp_val : _GEN_138 ? io_dis_uops_1_bits_fp_val : io_dis_uops_0_bits_fp_val),
    .io_in_uop_bits_fp_single       (_GEN_140 ? io_dis_uops_3_bits_fp_single : _GEN_139 ? io_dis_uops_2_bits_fp_single : _GEN_138 ? io_dis_uops_1_bits_fp_single : io_dis_uops_0_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if      (_GEN_140 ? io_dis_uops_3_bits_xcpt_pf_if : _GEN_139 ? io_dis_uops_2_bits_xcpt_pf_if : _GEN_138 ? io_dis_uops_1_bits_xcpt_pf_if : io_dis_uops_0_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if      (_GEN_140 ? io_dis_uops_3_bits_xcpt_ae_if : _GEN_139 ? io_dis_uops_2_bits_xcpt_ae_if : _GEN_138 ? io_dis_uops_1_bits_xcpt_ae_if : io_dis_uops_0_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if      (_GEN_140 ? io_dis_uops_3_bits_xcpt_ma_if : _GEN_139 ? io_dis_uops_2_bits_xcpt_ma_if : _GEN_138 ? io_dis_uops_1_bits_xcpt_ma_if : io_dis_uops_0_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if     (_GEN_140 ? io_dis_uops_3_bits_bp_debug_if : _GEN_139 ? io_dis_uops_2_bits_bp_debug_if : _GEN_138 ? io_dis_uops_1_bits_bp_debug_if : io_dis_uops_0_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if      (_GEN_140 ? io_dis_uops_3_bits_bp_xcpt_if : _GEN_139 ? io_dis_uops_2_bits_bp_xcpt_if : _GEN_138 ? io_dis_uops_1_bits_bp_xcpt_if : io_dis_uops_0_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc      (_GEN_140 ? io_dis_uops_3_bits_debug_fsrc : _GEN_139 ? io_dis_uops_2_bits_debug_fsrc : _GEN_138 ? io_dis_uops_1_bits_debug_fsrc : io_dis_uops_0_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc      (_GEN_140 ? io_dis_uops_3_bits_debug_tsrc : _GEN_139 ? io_dis_uops_2_bits_debug_tsrc : _GEN_138 ? io_dis_uops_1_bits_debug_tsrc : io_dis_uops_0_bits_debug_tsrc),
    .io_out_uop_uopc                (_slots_39_io_out_uop_uopc),
    .io_out_uop_inst                (_slots_39_io_out_uop_inst),
    .io_out_uop_debug_inst          (_slots_39_io_out_uop_debug_inst),
    .io_out_uop_is_rvc              (_slots_39_io_out_uop_is_rvc),
    .io_out_uop_debug_pc            (_slots_39_io_out_uop_debug_pc),
    .io_out_uop_iq_type             (_slots_39_io_out_uop_iq_type),
    .io_out_uop_fu_code             (_slots_39_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_39_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_39_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_39_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_39_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_39_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_39_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_39_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_39_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_39_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_39_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_39_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_39_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_39_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_39_io_out_uop_imm_packed),
    .io_out_uop_csr_addr            (_slots_39_io_out_uop_csr_addr),
    .io_out_uop_rob_idx             (_slots_39_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_39_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_39_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx             (_slots_39_io_out_uop_rxq_idx),
    .io_out_uop_pdst                (_slots_39_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_39_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_39_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_39_io_out_uop_prs3),
    .io_out_uop_ppred               (_slots_39_io_out_uop_ppred),
    .io_out_uop_prs1_busy           (_slots_39_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_39_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_39_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_39_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst          (_slots_39_io_out_uop_stale_pdst),
    .io_out_uop_exception           (_slots_39_io_out_uop_exception),
    .io_out_uop_exc_cause           (_slots_39_io_out_uop_exc_cause),
    .io_out_uop_bypassable          (_slots_39_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_39_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_39_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_39_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_39_io_out_uop_is_fence),
    .io_out_uop_is_fencei           (_slots_39_io_out_uop_is_fencei),
    .io_out_uop_is_amo              (_slots_39_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_39_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_39_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc       (_slots_39_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique           (_slots_39_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit     (_slots_39_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1         (_slots_39_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst                (_slots_39_io_out_uop_ldst),
    .io_out_uop_lrs1                (_slots_39_io_out_uop_lrs1),
    .io_out_uop_lrs2                (_slots_39_io_out_uop_lrs2),
    .io_out_uop_lrs3                (_slots_39_io_out_uop_lrs3),
    .io_out_uop_ldst_val            (_slots_39_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_39_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_39_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_39_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en             (_slots_39_io_out_uop_frs3_en),
    .io_out_uop_fp_val              (_slots_39_io_out_uop_fp_val),
    .io_out_uop_fp_single           (_slots_39_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if          (_slots_39_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if          (_slots_39_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if          (_slots_39_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if         (_slots_39_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if          (_slots_39_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc          (_slots_39_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc          (_slots_39_io_out_uop_debug_tsrc),
    .io_uop_uopc                    (_slots_39_io_uop_uopc),
    .io_uop_inst                    (_slots_39_io_uop_inst),
    .io_uop_debug_inst              (_slots_39_io_uop_debug_inst),
    .io_uop_is_rvc                  (_slots_39_io_uop_is_rvc),
    .io_uop_debug_pc                (_slots_39_io_uop_debug_pc),
    .io_uop_iq_type                 (_slots_39_io_uop_iq_type),
    .io_uop_fu_code                 (_slots_39_io_uop_fu_code),
    .io_uop_iw_state                (_slots_39_io_uop_iw_state),
    .io_uop_iw_p1_poisoned          (_slots_39_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_39_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_39_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_39_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_39_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_39_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_39_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_39_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_39_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_39_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_39_io_uop_pc_lob),
    .io_uop_taken                   (_slots_39_io_uop_taken),
    .io_uop_imm_packed              (_slots_39_io_uop_imm_packed),
    .io_uop_csr_addr                (_slots_39_io_uop_csr_addr),
    .io_uop_rob_idx                 (_slots_39_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_39_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_39_io_uop_stq_idx),
    .io_uop_rxq_idx                 (_slots_39_io_uop_rxq_idx),
    .io_uop_pdst                    (_slots_39_io_uop_pdst),
    .io_uop_prs1                    (_slots_39_io_uop_prs1),
    .io_uop_prs2                    (_slots_39_io_uop_prs2),
    .io_uop_prs3                    (_slots_39_io_uop_prs3),
    .io_uop_ppred                   (_slots_39_io_uop_ppred),
    .io_uop_prs1_busy               (_slots_39_io_uop_prs1_busy),
    .io_uop_prs2_busy               (_slots_39_io_uop_prs2_busy),
    .io_uop_prs3_busy               (_slots_39_io_uop_prs3_busy),
    .io_uop_ppred_busy              (_slots_39_io_uop_ppred_busy),
    .io_uop_stale_pdst              (_slots_39_io_uop_stale_pdst),
    .io_uop_exception               (_slots_39_io_uop_exception),
    .io_uop_exc_cause               (_slots_39_io_uop_exc_cause),
    .io_uop_bypassable              (_slots_39_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_39_io_uop_mem_cmd),
    .io_uop_mem_size                (_slots_39_io_uop_mem_size),
    .io_uop_mem_signed              (_slots_39_io_uop_mem_signed),
    .io_uop_is_fence                (_slots_39_io_uop_is_fence),
    .io_uop_is_fencei               (_slots_39_io_uop_is_fencei),
    .io_uop_is_amo                  (_slots_39_io_uop_is_amo),
    .io_uop_uses_ldq                (_slots_39_io_uop_uses_ldq),
    .io_uop_uses_stq                (_slots_39_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc           (_slots_39_io_uop_is_sys_pc2epc),
    .io_uop_is_unique               (_slots_39_io_uop_is_unique),
    .io_uop_flush_on_commit         (_slots_39_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1             (_slots_39_io_uop_ldst_is_rs1),
    .io_uop_ldst                    (_slots_39_io_uop_ldst),
    .io_uop_lrs1                    (_slots_39_io_uop_lrs1),
    .io_uop_lrs2                    (_slots_39_io_uop_lrs2),
    .io_uop_lrs3                    (_slots_39_io_uop_lrs3),
    .io_uop_ldst_val                (_slots_39_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_39_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_39_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_39_io_uop_lrs2_rtype),
    .io_uop_frs3_en                 (_slots_39_io_uop_frs3_en),
    .io_uop_fp_val                  (_slots_39_io_uop_fp_val),
    .io_uop_fp_single               (_slots_39_io_uop_fp_single),
    .io_uop_xcpt_pf_if              (_slots_39_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if              (_slots_39_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if              (_slots_39_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if             (_slots_39_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if              (_slots_39_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc              (_slots_39_io_uop_debug_fsrc),
    .io_uop_debug_tsrc              (_slots_39_io_uop_debug_tsrc)
  );
  assign io_dis_uops_0_ready = io_dis_uops_0_ready_REG;
  assign io_dis_uops_1_ready = io_dis_uops_1_ready_REG;
  assign io_dis_uops_2_ready = io_dis_uops_2_ready_REG;
  assign io_dis_uops_3_ready = io_dis_uops_3_ready_REG;
  assign io_iss_valids_0 = _GEN_677 | _GEN_666 | _GEN_652 | _GEN_638 | _GEN_624 | _GEN_610 | _GEN_596 | _GEN_582 | _GEN_568 | _GEN_554 | _GEN_540 | _GEN_526 | _GEN_512 | _GEN_498 | _GEN_484 | _GEN_470 | _GEN_456 | _GEN_442 | _GEN_428 | _GEN_414 | _GEN_400 | _GEN_386 | _GEN_372 | _GEN_358 | _GEN_344 | _GEN_330 | _GEN_316 | _GEN_302 | _GEN_288 | _GEN_274 | _GEN_260 | _GEN_246 | _GEN_232 | _GEN_218 | _GEN_204 | _GEN_190 | _GEN_176 | _GEN_162 | _GEN_148 | _GEN_141;
  assign io_iss_valids_1 = _GEN_679 | _GEN_669 | _GEN_656 | _GEN_642 | _GEN_628 | _GEN_614 | _GEN_600 | _GEN_586 | _GEN_572 | _GEN_558 | _GEN_544 | _GEN_530 | _GEN_516 | _GEN_502 | _GEN_488 | _GEN_474 | _GEN_460 | _GEN_446 | _GEN_432 | _GEN_418 | _GEN_404 | _GEN_390 | _GEN_376 | _GEN_362 | _GEN_348 | _GEN_334 | _GEN_320 | _GEN_306 | _GEN_292 | _GEN_278 | _GEN_264 | _GEN_250 | _GEN_236 | _GEN_222 | _GEN_208 | _GEN_194 | _GEN_180 | _GEN_166 | _GEN_152 | _GEN_143;
  assign io_iss_valids_2 = _GEN_681 | _GEN_673 | _GEN_660 | _GEN_646 | _GEN_632 | _GEN_618 | _GEN_604 | _GEN_590 | _GEN_576 | _GEN_562 | _GEN_548 | _GEN_534 | _GEN_520 | _GEN_506 | _GEN_492 | _GEN_478 | _GEN_464 | _GEN_450 | _GEN_436 | _GEN_422 | _GEN_408 | _GEN_394 | _GEN_380 | _GEN_366 | _GEN_352 | _GEN_338 | _GEN_324 | _GEN_310 | _GEN_296 | _GEN_282 | _GEN_268 | _GEN_254 | _GEN_240 | _GEN_226 | _GEN_212 | _GEN_198 | _GEN_184 | _GEN_170 | _GEN_156 | _GEN_145;
  assign io_iss_valids_3 = _GEN_682 | _GEN_676 | _GEN_663 | _GEN_649 | _GEN_635 | _GEN_621 | _GEN_607 | _GEN_593 | _GEN_579 | _GEN_565 | _GEN_551 | _GEN_537 | _GEN_523 | _GEN_509 | _GEN_495 | _GEN_481 | _GEN_467 | _GEN_453 | _GEN_439 | _GEN_425 | _GEN_411 | _GEN_397 | _GEN_383 | _GEN_369 | _GEN_355 | _GEN_341 | _GEN_327 | _GEN_313 | _GEN_299 | _GEN_285 | _GEN_271 | _GEN_257 | _GEN_243 | _GEN_229 | _GEN_215 | _GEN_201 | _GEN_187 | _GEN_173 | _GEN_159 | _GEN_146;
  assign io_iss_uops_0_uopc = _GEN_677 ? _slots_39_io_uop_uopc : _GEN_666 ? _slots_38_io_uop_uopc : _GEN_652 ? _slots_37_io_uop_uopc : _GEN_638 ? _slots_36_io_uop_uopc : _GEN_624 ? _slots_35_io_uop_uopc : _GEN_610 ? _slots_34_io_uop_uopc : _GEN_596 ? _slots_33_io_uop_uopc : _GEN_582 ? _slots_32_io_uop_uopc : _GEN_568 ? _slots_31_io_uop_uopc : _GEN_554 ? _slots_30_io_uop_uopc : _GEN_540 ? _slots_29_io_uop_uopc : _GEN_526 ? _slots_28_io_uop_uopc : _GEN_512 ? _slots_27_io_uop_uopc : _GEN_498 ? _slots_26_io_uop_uopc : _GEN_484 ? _slots_25_io_uop_uopc : _GEN_470 ? _slots_24_io_uop_uopc : _GEN_456 ? _slots_23_io_uop_uopc : _GEN_442 ? _slots_22_io_uop_uopc : _GEN_428 ? _slots_21_io_uop_uopc : _GEN_414 ? _slots_20_io_uop_uopc : _GEN_400 ? _slots_19_io_uop_uopc : _GEN_386 ? _slots_18_io_uop_uopc : _GEN_372 ? _slots_17_io_uop_uopc : _GEN_358 ? _slots_16_io_uop_uopc : _GEN_344 ? _slots_15_io_uop_uopc : _GEN_330 ? _slots_14_io_uop_uopc : _GEN_316 ? _slots_13_io_uop_uopc : _GEN_302 ? _slots_12_io_uop_uopc : _GEN_288 ? _slots_11_io_uop_uopc : _GEN_274 ? _slots_10_io_uop_uopc : _GEN_260 ? _slots_9_io_uop_uopc : _GEN_246 ? _slots_8_io_uop_uopc : _GEN_232 ? _slots_7_io_uop_uopc : _GEN_218 ? _slots_6_io_uop_uopc : _GEN_204 ? _slots_5_io_uop_uopc : _GEN_190 ? _slots_4_io_uop_uopc : _GEN_176 ? _slots_3_io_uop_uopc : _GEN_162 ? _slots_2_io_uop_uopc : _GEN_148 ? _slots_1_io_uop_uopc : _GEN_141 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_0_inst = _GEN_677 ? _slots_39_io_uop_inst : _GEN_666 ? _slots_38_io_uop_inst : _GEN_652 ? _slots_37_io_uop_inst : _GEN_638 ? _slots_36_io_uop_inst : _GEN_624 ? _slots_35_io_uop_inst : _GEN_610 ? _slots_34_io_uop_inst : _GEN_596 ? _slots_33_io_uop_inst : _GEN_582 ? _slots_32_io_uop_inst : _GEN_568 ? _slots_31_io_uop_inst : _GEN_554 ? _slots_30_io_uop_inst : _GEN_540 ? _slots_29_io_uop_inst : _GEN_526 ? _slots_28_io_uop_inst : _GEN_512 ? _slots_27_io_uop_inst : _GEN_498 ? _slots_26_io_uop_inst : _GEN_484 ? _slots_25_io_uop_inst : _GEN_470 ? _slots_24_io_uop_inst : _GEN_456 ? _slots_23_io_uop_inst : _GEN_442 ? _slots_22_io_uop_inst : _GEN_428 ? _slots_21_io_uop_inst : _GEN_414 ? _slots_20_io_uop_inst : _GEN_400 ? _slots_19_io_uop_inst : _GEN_386 ? _slots_18_io_uop_inst : _GEN_372 ? _slots_17_io_uop_inst : _GEN_358 ? _slots_16_io_uop_inst : _GEN_344 ? _slots_15_io_uop_inst : _GEN_330 ? _slots_14_io_uop_inst : _GEN_316 ? _slots_13_io_uop_inst : _GEN_302 ? _slots_12_io_uop_inst : _GEN_288 ? _slots_11_io_uop_inst : _GEN_274 ? _slots_10_io_uop_inst : _GEN_260 ? _slots_9_io_uop_inst : _GEN_246 ? _slots_8_io_uop_inst : _GEN_232 ? _slots_7_io_uop_inst : _GEN_218 ? _slots_6_io_uop_inst : _GEN_204 ? _slots_5_io_uop_inst : _GEN_190 ? _slots_4_io_uop_inst : _GEN_176 ? _slots_3_io_uop_inst : _GEN_162 ? _slots_2_io_uop_inst : _GEN_148 ? _slots_1_io_uop_inst : _GEN_141 ? _slots_0_io_uop_inst : 32'h0;
  assign io_iss_uops_0_debug_inst = _GEN_677 ? _slots_39_io_uop_debug_inst : _GEN_666 ? _slots_38_io_uop_debug_inst : _GEN_652 ? _slots_37_io_uop_debug_inst : _GEN_638 ? _slots_36_io_uop_debug_inst : _GEN_624 ? _slots_35_io_uop_debug_inst : _GEN_610 ? _slots_34_io_uop_debug_inst : _GEN_596 ? _slots_33_io_uop_debug_inst : _GEN_582 ? _slots_32_io_uop_debug_inst : _GEN_568 ? _slots_31_io_uop_debug_inst : _GEN_554 ? _slots_30_io_uop_debug_inst : _GEN_540 ? _slots_29_io_uop_debug_inst : _GEN_526 ? _slots_28_io_uop_debug_inst : _GEN_512 ? _slots_27_io_uop_debug_inst : _GEN_498 ? _slots_26_io_uop_debug_inst : _GEN_484 ? _slots_25_io_uop_debug_inst : _GEN_470 ? _slots_24_io_uop_debug_inst : _GEN_456 ? _slots_23_io_uop_debug_inst : _GEN_442 ? _slots_22_io_uop_debug_inst : _GEN_428 ? _slots_21_io_uop_debug_inst : _GEN_414 ? _slots_20_io_uop_debug_inst : _GEN_400 ? _slots_19_io_uop_debug_inst : _GEN_386 ? _slots_18_io_uop_debug_inst : _GEN_372 ? _slots_17_io_uop_debug_inst : _GEN_358 ? _slots_16_io_uop_debug_inst : _GEN_344 ? _slots_15_io_uop_debug_inst : _GEN_330 ? _slots_14_io_uop_debug_inst : _GEN_316 ? _slots_13_io_uop_debug_inst : _GEN_302 ? _slots_12_io_uop_debug_inst : _GEN_288 ? _slots_11_io_uop_debug_inst : _GEN_274 ? _slots_10_io_uop_debug_inst : _GEN_260 ? _slots_9_io_uop_debug_inst : _GEN_246 ? _slots_8_io_uop_debug_inst : _GEN_232 ? _slots_7_io_uop_debug_inst : _GEN_218 ? _slots_6_io_uop_debug_inst : _GEN_204 ? _slots_5_io_uop_debug_inst : _GEN_190 ? _slots_4_io_uop_debug_inst : _GEN_176 ? _slots_3_io_uop_debug_inst : _GEN_162 ? _slots_2_io_uop_debug_inst : _GEN_148 ? _slots_1_io_uop_debug_inst : _GEN_141 ? _slots_0_io_uop_debug_inst : 32'h0;
  assign io_iss_uops_0_is_rvc = _GEN_677 ? _slots_39_io_uop_is_rvc : _GEN_666 ? _slots_38_io_uop_is_rvc : _GEN_652 ? _slots_37_io_uop_is_rvc : _GEN_638 ? _slots_36_io_uop_is_rvc : _GEN_624 ? _slots_35_io_uop_is_rvc : _GEN_610 ? _slots_34_io_uop_is_rvc : _GEN_596 ? _slots_33_io_uop_is_rvc : _GEN_582 ? _slots_32_io_uop_is_rvc : _GEN_568 ? _slots_31_io_uop_is_rvc : _GEN_554 ? _slots_30_io_uop_is_rvc : _GEN_540 ? _slots_29_io_uop_is_rvc : _GEN_526 ? _slots_28_io_uop_is_rvc : _GEN_512 ? _slots_27_io_uop_is_rvc : _GEN_498 ? _slots_26_io_uop_is_rvc : _GEN_484 ? _slots_25_io_uop_is_rvc : _GEN_470 ? _slots_24_io_uop_is_rvc : _GEN_456 ? _slots_23_io_uop_is_rvc : _GEN_442 ? _slots_22_io_uop_is_rvc : _GEN_428 ? _slots_21_io_uop_is_rvc : _GEN_414 ? _slots_20_io_uop_is_rvc : _GEN_400 ? _slots_19_io_uop_is_rvc : _GEN_386 ? _slots_18_io_uop_is_rvc : _GEN_372 ? _slots_17_io_uop_is_rvc : _GEN_358 ? _slots_16_io_uop_is_rvc : _GEN_344 ? _slots_15_io_uop_is_rvc : _GEN_330 ? _slots_14_io_uop_is_rvc : _GEN_316 ? _slots_13_io_uop_is_rvc : _GEN_302 ? _slots_12_io_uop_is_rvc : _GEN_288 ? _slots_11_io_uop_is_rvc : _GEN_274 ? _slots_10_io_uop_is_rvc : _GEN_260 ? _slots_9_io_uop_is_rvc : _GEN_246 ? _slots_8_io_uop_is_rvc : _GEN_232 ? _slots_7_io_uop_is_rvc : _GEN_218 ? _slots_6_io_uop_is_rvc : _GEN_204 ? _slots_5_io_uop_is_rvc : _GEN_190 ? _slots_4_io_uop_is_rvc : _GEN_176 ? _slots_3_io_uop_is_rvc : _GEN_162 ? _slots_2_io_uop_is_rvc : _GEN_148 ? _slots_1_io_uop_is_rvc : _GEN_141 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_0_debug_pc = _GEN_677 ? _slots_39_io_uop_debug_pc : _GEN_666 ? _slots_38_io_uop_debug_pc : _GEN_652 ? _slots_37_io_uop_debug_pc : _GEN_638 ? _slots_36_io_uop_debug_pc : _GEN_624 ? _slots_35_io_uop_debug_pc : _GEN_610 ? _slots_34_io_uop_debug_pc : _GEN_596 ? _slots_33_io_uop_debug_pc : _GEN_582 ? _slots_32_io_uop_debug_pc : _GEN_568 ? _slots_31_io_uop_debug_pc : _GEN_554 ? _slots_30_io_uop_debug_pc : _GEN_540 ? _slots_29_io_uop_debug_pc : _GEN_526 ? _slots_28_io_uop_debug_pc : _GEN_512 ? _slots_27_io_uop_debug_pc : _GEN_498 ? _slots_26_io_uop_debug_pc : _GEN_484 ? _slots_25_io_uop_debug_pc : _GEN_470 ? _slots_24_io_uop_debug_pc : _GEN_456 ? _slots_23_io_uop_debug_pc : _GEN_442 ? _slots_22_io_uop_debug_pc : _GEN_428 ? _slots_21_io_uop_debug_pc : _GEN_414 ? _slots_20_io_uop_debug_pc : _GEN_400 ? _slots_19_io_uop_debug_pc : _GEN_386 ? _slots_18_io_uop_debug_pc : _GEN_372 ? _slots_17_io_uop_debug_pc : _GEN_358 ? _slots_16_io_uop_debug_pc : _GEN_344 ? _slots_15_io_uop_debug_pc : _GEN_330 ? _slots_14_io_uop_debug_pc : _GEN_316 ? _slots_13_io_uop_debug_pc : _GEN_302 ? _slots_12_io_uop_debug_pc : _GEN_288 ? _slots_11_io_uop_debug_pc : _GEN_274 ? _slots_10_io_uop_debug_pc : _GEN_260 ? _slots_9_io_uop_debug_pc : _GEN_246 ? _slots_8_io_uop_debug_pc : _GEN_232 ? _slots_7_io_uop_debug_pc : _GEN_218 ? _slots_6_io_uop_debug_pc : _GEN_204 ? _slots_5_io_uop_debug_pc : _GEN_190 ? _slots_4_io_uop_debug_pc : _GEN_176 ? _slots_3_io_uop_debug_pc : _GEN_162 ? _slots_2_io_uop_debug_pc : _GEN_148 ? _slots_1_io_uop_debug_pc : _GEN_141 ? _slots_0_io_uop_debug_pc : 40'h0;
  assign io_iss_uops_0_iq_type = _GEN_677 ? _slots_39_io_uop_iq_type : _GEN_666 ? _slots_38_io_uop_iq_type : _GEN_652 ? _slots_37_io_uop_iq_type : _GEN_638 ? _slots_36_io_uop_iq_type : _GEN_624 ? _slots_35_io_uop_iq_type : _GEN_610 ? _slots_34_io_uop_iq_type : _GEN_596 ? _slots_33_io_uop_iq_type : _GEN_582 ? _slots_32_io_uop_iq_type : _GEN_568 ? _slots_31_io_uop_iq_type : _GEN_554 ? _slots_30_io_uop_iq_type : _GEN_540 ? _slots_29_io_uop_iq_type : _GEN_526 ? _slots_28_io_uop_iq_type : _GEN_512 ? _slots_27_io_uop_iq_type : _GEN_498 ? _slots_26_io_uop_iq_type : _GEN_484 ? _slots_25_io_uop_iq_type : _GEN_470 ? _slots_24_io_uop_iq_type : _GEN_456 ? _slots_23_io_uop_iq_type : _GEN_442 ? _slots_22_io_uop_iq_type : _GEN_428 ? _slots_21_io_uop_iq_type : _GEN_414 ? _slots_20_io_uop_iq_type : _GEN_400 ? _slots_19_io_uop_iq_type : _GEN_386 ? _slots_18_io_uop_iq_type : _GEN_372 ? _slots_17_io_uop_iq_type : _GEN_358 ? _slots_16_io_uop_iq_type : _GEN_344 ? _slots_15_io_uop_iq_type : _GEN_330 ? _slots_14_io_uop_iq_type : _GEN_316 ? _slots_13_io_uop_iq_type : _GEN_302 ? _slots_12_io_uop_iq_type : _GEN_288 ? _slots_11_io_uop_iq_type : _GEN_274 ? _slots_10_io_uop_iq_type : _GEN_260 ? _slots_9_io_uop_iq_type : _GEN_246 ? _slots_8_io_uop_iq_type : _GEN_232 ? _slots_7_io_uop_iq_type : _GEN_218 ? _slots_6_io_uop_iq_type : _GEN_204 ? _slots_5_io_uop_iq_type : _GEN_190 ? _slots_4_io_uop_iq_type : _GEN_176 ? _slots_3_io_uop_iq_type : _GEN_162 ? _slots_2_io_uop_iq_type : _GEN_148 ? _slots_1_io_uop_iq_type : _GEN_141 ? _slots_0_io_uop_iq_type : 3'h0;
  assign io_iss_uops_0_fu_code = _GEN_677 ? _slots_39_io_uop_fu_code : _GEN_666 ? _slots_38_io_uop_fu_code : _GEN_652 ? _slots_37_io_uop_fu_code : _GEN_638 ? _slots_36_io_uop_fu_code : _GEN_624 ? _slots_35_io_uop_fu_code : _GEN_610 ? _slots_34_io_uop_fu_code : _GEN_596 ? _slots_33_io_uop_fu_code : _GEN_582 ? _slots_32_io_uop_fu_code : _GEN_568 ? _slots_31_io_uop_fu_code : _GEN_554 ? _slots_30_io_uop_fu_code : _GEN_540 ? _slots_29_io_uop_fu_code : _GEN_526 ? _slots_28_io_uop_fu_code : _GEN_512 ? _slots_27_io_uop_fu_code : _GEN_498 ? _slots_26_io_uop_fu_code : _GEN_484 ? _slots_25_io_uop_fu_code : _GEN_470 ? _slots_24_io_uop_fu_code : _GEN_456 ? _slots_23_io_uop_fu_code : _GEN_442 ? _slots_22_io_uop_fu_code : _GEN_428 ? _slots_21_io_uop_fu_code : _GEN_414 ? _slots_20_io_uop_fu_code : _GEN_400 ? _slots_19_io_uop_fu_code : _GEN_386 ? _slots_18_io_uop_fu_code : _GEN_372 ? _slots_17_io_uop_fu_code : _GEN_358 ? _slots_16_io_uop_fu_code : _GEN_344 ? _slots_15_io_uop_fu_code : _GEN_330 ? _slots_14_io_uop_fu_code : _GEN_316 ? _slots_13_io_uop_fu_code : _GEN_302 ? _slots_12_io_uop_fu_code : _GEN_288 ? _slots_11_io_uop_fu_code : _GEN_274 ? _slots_10_io_uop_fu_code : _GEN_260 ? _slots_9_io_uop_fu_code : _GEN_246 ? _slots_8_io_uop_fu_code : _GEN_232 ? _slots_7_io_uop_fu_code : _GEN_218 ? _slots_6_io_uop_fu_code : _GEN_204 ? _slots_5_io_uop_fu_code : _GEN_190 ? _slots_4_io_uop_fu_code : _GEN_176 ? _slots_3_io_uop_fu_code : _GEN_162 ? _slots_2_io_uop_fu_code : _GEN_148 ? _slots_1_io_uop_fu_code : _GEN_141 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_0_iw_state = _GEN_677 ? _slots_39_io_uop_iw_state : _GEN_666 ? _slots_38_io_uop_iw_state : _GEN_652 ? _slots_37_io_uop_iw_state : _GEN_638 ? _slots_36_io_uop_iw_state : _GEN_624 ? _slots_35_io_uop_iw_state : _GEN_610 ? _slots_34_io_uop_iw_state : _GEN_596 ? _slots_33_io_uop_iw_state : _GEN_582 ? _slots_32_io_uop_iw_state : _GEN_568 ? _slots_31_io_uop_iw_state : _GEN_554 ? _slots_30_io_uop_iw_state : _GEN_540 ? _slots_29_io_uop_iw_state : _GEN_526 ? _slots_28_io_uop_iw_state : _GEN_512 ? _slots_27_io_uop_iw_state : _GEN_498 ? _slots_26_io_uop_iw_state : _GEN_484 ? _slots_25_io_uop_iw_state : _GEN_470 ? _slots_24_io_uop_iw_state : _GEN_456 ? _slots_23_io_uop_iw_state : _GEN_442 ? _slots_22_io_uop_iw_state : _GEN_428 ? _slots_21_io_uop_iw_state : _GEN_414 ? _slots_20_io_uop_iw_state : _GEN_400 ? _slots_19_io_uop_iw_state : _GEN_386 ? _slots_18_io_uop_iw_state : _GEN_372 ? _slots_17_io_uop_iw_state : _GEN_358 ? _slots_16_io_uop_iw_state : _GEN_344 ? _slots_15_io_uop_iw_state : _GEN_330 ? _slots_14_io_uop_iw_state : _GEN_316 ? _slots_13_io_uop_iw_state : _GEN_302 ? _slots_12_io_uop_iw_state : _GEN_288 ? _slots_11_io_uop_iw_state : _GEN_274 ? _slots_10_io_uop_iw_state : _GEN_260 ? _slots_9_io_uop_iw_state : _GEN_246 ? _slots_8_io_uop_iw_state : _GEN_232 ? _slots_7_io_uop_iw_state : _GEN_218 ? _slots_6_io_uop_iw_state : _GEN_204 ? _slots_5_io_uop_iw_state : _GEN_190 ? _slots_4_io_uop_iw_state : _GEN_176 ? _slots_3_io_uop_iw_state : _GEN_162 ? _slots_2_io_uop_iw_state : _GEN_148 ? _slots_1_io_uop_iw_state : _GEN_141 ? _slots_0_io_uop_iw_state : 2'h0;
  assign io_iss_uops_0_iw_p1_poisoned = _GEN_677 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_666 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_652 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_638 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_624 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_610 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_596 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_582 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_568 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_554 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_540 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_526 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_512 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_498 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_484 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_470 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_456 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_442 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_428 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_414 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_400 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_386 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_372 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_358 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_344 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_330 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_316 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_302 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_288 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_274 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_260 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_246 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_232 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_218 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_204 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_190 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_176 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_162 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_148 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_141 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_0_iw_p2_poisoned = _GEN_677 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_666 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_652 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_638 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_624 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_610 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_596 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_582 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_568 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_554 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_540 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_526 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_512 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_498 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_484 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_470 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_456 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_442 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_428 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_414 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_400 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_386 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_372 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_358 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_344 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_330 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_316 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_302 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_288 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_274 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_260 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_246 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_232 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_218 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_204 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_190 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_176 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_162 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_148 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_141 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_0_is_br = _GEN_677 ? _slots_39_io_uop_is_br : _GEN_666 ? _slots_38_io_uop_is_br : _GEN_652 ? _slots_37_io_uop_is_br : _GEN_638 ? _slots_36_io_uop_is_br : _GEN_624 ? _slots_35_io_uop_is_br : _GEN_610 ? _slots_34_io_uop_is_br : _GEN_596 ? _slots_33_io_uop_is_br : _GEN_582 ? _slots_32_io_uop_is_br : _GEN_568 ? _slots_31_io_uop_is_br : _GEN_554 ? _slots_30_io_uop_is_br : _GEN_540 ? _slots_29_io_uop_is_br : _GEN_526 ? _slots_28_io_uop_is_br : _GEN_512 ? _slots_27_io_uop_is_br : _GEN_498 ? _slots_26_io_uop_is_br : _GEN_484 ? _slots_25_io_uop_is_br : _GEN_470 ? _slots_24_io_uop_is_br : _GEN_456 ? _slots_23_io_uop_is_br : _GEN_442 ? _slots_22_io_uop_is_br : _GEN_428 ? _slots_21_io_uop_is_br : _GEN_414 ? _slots_20_io_uop_is_br : _GEN_400 ? _slots_19_io_uop_is_br : _GEN_386 ? _slots_18_io_uop_is_br : _GEN_372 ? _slots_17_io_uop_is_br : _GEN_358 ? _slots_16_io_uop_is_br : _GEN_344 ? _slots_15_io_uop_is_br : _GEN_330 ? _slots_14_io_uop_is_br : _GEN_316 ? _slots_13_io_uop_is_br : _GEN_302 ? _slots_12_io_uop_is_br : _GEN_288 ? _slots_11_io_uop_is_br : _GEN_274 ? _slots_10_io_uop_is_br : _GEN_260 ? _slots_9_io_uop_is_br : _GEN_246 ? _slots_8_io_uop_is_br : _GEN_232 ? _slots_7_io_uop_is_br : _GEN_218 ? _slots_6_io_uop_is_br : _GEN_204 ? _slots_5_io_uop_is_br : _GEN_190 ? _slots_4_io_uop_is_br : _GEN_176 ? _slots_3_io_uop_is_br : _GEN_162 ? _slots_2_io_uop_is_br : _GEN_148 ? _slots_1_io_uop_is_br : _GEN_141 & _slots_0_io_uop_is_br;
  assign io_iss_uops_0_is_jalr = _GEN_677 ? _slots_39_io_uop_is_jalr : _GEN_666 ? _slots_38_io_uop_is_jalr : _GEN_652 ? _slots_37_io_uop_is_jalr : _GEN_638 ? _slots_36_io_uop_is_jalr : _GEN_624 ? _slots_35_io_uop_is_jalr : _GEN_610 ? _slots_34_io_uop_is_jalr : _GEN_596 ? _slots_33_io_uop_is_jalr : _GEN_582 ? _slots_32_io_uop_is_jalr : _GEN_568 ? _slots_31_io_uop_is_jalr : _GEN_554 ? _slots_30_io_uop_is_jalr : _GEN_540 ? _slots_29_io_uop_is_jalr : _GEN_526 ? _slots_28_io_uop_is_jalr : _GEN_512 ? _slots_27_io_uop_is_jalr : _GEN_498 ? _slots_26_io_uop_is_jalr : _GEN_484 ? _slots_25_io_uop_is_jalr : _GEN_470 ? _slots_24_io_uop_is_jalr : _GEN_456 ? _slots_23_io_uop_is_jalr : _GEN_442 ? _slots_22_io_uop_is_jalr : _GEN_428 ? _slots_21_io_uop_is_jalr : _GEN_414 ? _slots_20_io_uop_is_jalr : _GEN_400 ? _slots_19_io_uop_is_jalr : _GEN_386 ? _slots_18_io_uop_is_jalr : _GEN_372 ? _slots_17_io_uop_is_jalr : _GEN_358 ? _slots_16_io_uop_is_jalr : _GEN_344 ? _slots_15_io_uop_is_jalr : _GEN_330 ? _slots_14_io_uop_is_jalr : _GEN_316 ? _slots_13_io_uop_is_jalr : _GEN_302 ? _slots_12_io_uop_is_jalr : _GEN_288 ? _slots_11_io_uop_is_jalr : _GEN_274 ? _slots_10_io_uop_is_jalr : _GEN_260 ? _slots_9_io_uop_is_jalr : _GEN_246 ? _slots_8_io_uop_is_jalr : _GEN_232 ? _slots_7_io_uop_is_jalr : _GEN_218 ? _slots_6_io_uop_is_jalr : _GEN_204 ? _slots_5_io_uop_is_jalr : _GEN_190 ? _slots_4_io_uop_is_jalr : _GEN_176 ? _slots_3_io_uop_is_jalr : _GEN_162 ? _slots_2_io_uop_is_jalr : _GEN_148 ? _slots_1_io_uop_is_jalr : _GEN_141 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_0_is_jal = _GEN_677 ? _slots_39_io_uop_is_jal : _GEN_666 ? _slots_38_io_uop_is_jal : _GEN_652 ? _slots_37_io_uop_is_jal : _GEN_638 ? _slots_36_io_uop_is_jal : _GEN_624 ? _slots_35_io_uop_is_jal : _GEN_610 ? _slots_34_io_uop_is_jal : _GEN_596 ? _slots_33_io_uop_is_jal : _GEN_582 ? _slots_32_io_uop_is_jal : _GEN_568 ? _slots_31_io_uop_is_jal : _GEN_554 ? _slots_30_io_uop_is_jal : _GEN_540 ? _slots_29_io_uop_is_jal : _GEN_526 ? _slots_28_io_uop_is_jal : _GEN_512 ? _slots_27_io_uop_is_jal : _GEN_498 ? _slots_26_io_uop_is_jal : _GEN_484 ? _slots_25_io_uop_is_jal : _GEN_470 ? _slots_24_io_uop_is_jal : _GEN_456 ? _slots_23_io_uop_is_jal : _GEN_442 ? _slots_22_io_uop_is_jal : _GEN_428 ? _slots_21_io_uop_is_jal : _GEN_414 ? _slots_20_io_uop_is_jal : _GEN_400 ? _slots_19_io_uop_is_jal : _GEN_386 ? _slots_18_io_uop_is_jal : _GEN_372 ? _slots_17_io_uop_is_jal : _GEN_358 ? _slots_16_io_uop_is_jal : _GEN_344 ? _slots_15_io_uop_is_jal : _GEN_330 ? _slots_14_io_uop_is_jal : _GEN_316 ? _slots_13_io_uop_is_jal : _GEN_302 ? _slots_12_io_uop_is_jal : _GEN_288 ? _slots_11_io_uop_is_jal : _GEN_274 ? _slots_10_io_uop_is_jal : _GEN_260 ? _slots_9_io_uop_is_jal : _GEN_246 ? _slots_8_io_uop_is_jal : _GEN_232 ? _slots_7_io_uop_is_jal : _GEN_218 ? _slots_6_io_uop_is_jal : _GEN_204 ? _slots_5_io_uop_is_jal : _GEN_190 ? _slots_4_io_uop_is_jal : _GEN_176 ? _slots_3_io_uop_is_jal : _GEN_162 ? _slots_2_io_uop_is_jal : _GEN_148 ? _slots_1_io_uop_is_jal : _GEN_141 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_0_is_sfb = _GEN_677 ? _slots_39_io_uop_is_sfb : _GEN_666 ? _slots_38_io_uop_is_sfb : _GEN_652 ? _slots_37_io_uop_is_sfb : _GEN_638 ? _slots_36_io_uop_is_sfb : _GEN_624 ? _slots_35_io_uop_is_sfb : _GEN_610 ? _slots_34_io_uop_is_sfb : _GEN_596 ? _slots_33_io_uop_is_sfb : _GEN_582 ? _slots_32_io_uop_is_sfb : _GEN_568 ? _slots_31_io_uop_is_sfb : _GEN_554 ? _slots_30_io_uop_is_sfb : _GEN_540 ? _slots_29_io_uop_is_sfb : _GEN_526 ? _slots_28_io_uop_is_sfb : _GEN_512 ? _slots_27_io_uop_is_sfb : _GEN_498 ? _slots_26_io_uop_is_sfb : _GEN_484 ? _slots_25_io_uop_is_sfb : _GEN_470 ? _slots_24_io_uop_is_sfb : _GEN_456 ? _slots_23_io_uop_is_sfb : _GEN_442 ? _slots_22_io_uop_is_sfb : _GEN_428 ? _slots_21_io_uop_is_sfb : _GEN_414 ? _slots_20_io_uop_is_sfb : _GEN_400 ? _slots_19_io_uop_is_sfb : _GEN_386 ? _slots_18_io_uop_is_sfb : _GEN_372 ? _slots_17_io_uop_is_sfb : _GEN_358 ? _slots_16_io_uop_is_sfb : _GEN_344 ? _slots_15_io_uop_is_sfb : _GEN_330 ? _slots_14_io_uop_is_sfb : _GEN_316 ? _slots_13_io_uop_is_sfb : _GEN_302 ? _slots_12_io_uop_is_sfb : _GEN_288 ? _slots_11_io_uop_is_sfb : _GEN_274 ? _slots_10_io_uop_is_sfb : _GEN_260 ? _slots_9_io_uop_is_sfb : _GEN_246 ? _slots_8_io_uop_is_sfb : _GEN_232 ? _slots_7_io_uop_is_sfb : _GEN_218 ? _slots_6_io_uop_is_sfb : _GEN_204 ? _slots_5_io_uop_is_sfb : _GEN_190 ? _slots_4_io_uop_is_sfb : _GEN_176 ? _slots_3_io_uop_is_sfb : _GEN_162 ? _slots_2_io_uop_is_sfb : _GEN_148 ? _slots_1_io_uop_is_sfb : _GEN_141 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_0_br_mask = _GEN_677 ? _slots_39_io_uop_br_mask : _GEN_666 ? _slots_38_io_uop_br_mask : _GEN_652 ? _slots_37_io_uop_br_mask : _GEN_638 ? _slots_36_io_uop_br_mask : _GEN_624 ? _slots_35_io_uop_br_mask : _GEN_610 ? _slots_34_io_uop_br_mask : _GEN_596 ? _slots_33_io_uop_br_mask : _GEN_582 ? _slots_32_io_uop_br_mask : _GEN_568 ? _slots_31_io_uop_br_mask : _GEN_554 ? _slots_30_io_uop_br_mask : _GEN_540 ? _slots_29_io_uop_br_mask : _GEN_526 ? _slots_28_io_uop_br_mask : _GEN_512 ? _slots_27_io_uop_br_mask : _GEN_498 ? _slots_26_io_uop_br_mask : _GEN_484 ? _slots_25_io_uop_br_mask : _GEN_470 ? _slots_24_io_uop_br_mask : _GEN_456 ? _slots_23_io_uop_br_mask : _GEN_442 ? _slots_22_io_uop_br_mask : _GEN_428 ? _slots_21_io_uop_br_mask : _GEN_414 ? _slots_20_io_uop_br_mask : _GEN_400 ? _slots_19_io_uop_br_mask : _GEN_386 ? _slots_18_io_uop_br_mask : _GEN_372 ? _slots_17_io_uop_br_mask : _GEN_358 ? _slots_16_io_uop_br_mask : _GEN_344 ? _slots_15_io_uop_br_mask : _GEN_330 ? _slots_14_io_uop_br_mask : _GEN_316 ? _slots_13_io_uop_br_mask : _GEN_302 ? _slots_12_io_uop_br_mask : _GEN_288 ? _slots_11_io_uop_br_mask : _GEN_274 ? _slots_10_io_uop_br_mask : _GEN_260 ? _slots_9_io_uop_br_mask : _GEN_246 ? _slots_8_io_uop_br_mask : _GEN_232 ? _slots_7_io_uop_br_mask : _GEN_218 ? _slots_6_io_uop_br_mask : _GEN_204 ? _slots_5_io_uop_br_mask : _GEN_190 ? _slots_4_io_uop_br_mask : _GEN_176 ? _slots_3_io_uop_br_mask : _GEN_162 ? _slots_2_io_uop_br_mask : _GEN_148 ? _slots_1_io_uop_br_mask : _GEN_141 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_0_br_tag = _GEN_677 ? _slots_39_io_uop_br_tag : _GEN_666 ? _slots_38_io_uop_br_tag : _GEN_652 ? _slots_37_io_uop_br_tag : _GEN_638 ? _slots_36_io_uop_br_tag : _GEN_624 ? _slots_35_io_uop_br_tag : _GEN_610 ? _slots_34_io_uop_br_tag : _GEN_596 ? _slots_33_io_uop_br_tag : _GEN_582 ? _slots_32_io_uop_br_tag : _GEN_568 ? _slots_31_io_uop_br_tag : _GEN_554 ? _slots_30_io_uop_br_tag : _GEN_540 ? _slots_29_io_uop_br_tag : _GEN_526 ? _slots_28_io_uop_br_tag : _GEN_512 ? _slots_27_io_uop_br_tag : _GEN_498 ? _slots_26_io_uop_br_tag : _GEN_484 ? _slots_25_io_uop_br_tag : _GEN_470 ? _slots_24_io_uop_br_tag : _GEN_456 ? _slots_23_io_uop_br_tag : _GEN_442 ? _slots_22_io_uop_br_tag : _GEN_428 ? _slots_21_io_uop_br_tag : _GEN_414 ? _slots_20_io_uop_br_tag : _GEN_400 ? _slots_19_io_uop_br_tag : _GEN_386 ? _slots_18_io_uop_br_tag : _GEN_372 ? _slots_17_io_uop_br_tag : _GEN_358 ? _slots_16_io_uop_br_tag : _GEN_344 ? _slots_15_io_uop_br_tag : _GEN_330 ? _slots_14_io_uop_br_tag : _GEN_316 ? _slots_13_io_uop_br_tag : _GEN_302 ? _slots_12_io_uop_br_tag : _GEN_288 ? _slots_11_io_uop_br_tag : _GEN_274 ? _slots_10_io_uop_br_tag : _GEN_260 ? _slots_9_io_uop_br_tag : _GEN_246 ? _slots_8_io_uop_br_tag : _GEN_232 ? _slots_7_io_uop_br_tag : _GEN_218 ? _slots_6_io_uop_br_tag : _GEN_204 ? _slots_5_io_uop_br_tag : _GEN_190 ? _slots_4_io_uop_br_tag : _GEN_176 ? _slots_3_io_uop_br_tag : _GEN_162 ? _slots_2_io_uop_br_tag : _GEN_148 ? _slots_1_io_uop_br_tag : _GEN_141 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_0_ftq_idx = _GEN_677 ? _slots_39_io_uop_ftq_idx : _GEN_666 ? _slots_38_io_uop_ftq_idx : _GEN_652 ? _slots_37_io_uop_ftq_idx : _GEN_638 ? _slots_36_io_uop_ftq_idx : _GEN_624 ? _slots_35_io_uop_ftq_idx : _GEN_610 ? _slots_34_io_uop_ftq_idx : _GEN_596 ? _slots_33_io_uop_ftq_idx : _GEN_582 ? _slots_32_io_uop_ftq_idx : _GEN_568 ? _slots_31_io_uop_ftq_idx : _GEN_554 ? _slots_30_io_uop_ftq_idx : _GEN_540 ? _slots_29_io_uop_ftq_idx : _GEN_526 ? _slots_28_io_uop_ftq_idx : _GEN_512 ? _slots_27_io_uop_ftq_idx : _GEN_498 ? _slots_26_io_uop_ftq_idx : _GEN_484 ? _slots_25_io_uop_ftq_idx : _GEN_470 ? _slots_24_io_uop_ftq_idx : _GEN_456 ? _slots_23_io_uop_ftq_idx : _GEN_442 ? _slots_22_io_uop_ftq_idx : _GEN_428 ? _slots_21_io_uop_ftq_idx : _GEN_414 ? _slots_20_io_uop_ftq_idx : _GEN_400 ? _slots_19_io_uop_ftq_idx : _GEN_386 ? _slots_18_io_uop_ftq_idx : _GEN_372 ? _slots_17_io_uop_ftq_idx : _GEN_358 ? _slots_16_io_uop_ftq_idx : _GEN_344 ? _slots_15_io_uop_ftq_idx : _GEN_330 ? _slots_14_io_uop_ftq_idx : _GEN_316 ? _slots_13_io_uop_ftq_idx : _GEN_302 ? _slots_12_io_uop_ftq_idx : _GEN_288 ? _slots_11_io_uop_ftq_idx : _GEN_274 ? _slots_10_io_uop_ftq_idx : _GEN_260 ? _slots_9_io_uop_ftq_idx : _GEN_246 ? _slots_8_io_uop_ftq_idx : _GEN_232 ? _slots_7_io_uop_ftq_idx : _GEN_218 ? _slots_6_io_uop_ftq_idx : _GEN_204 ? _slots_5_io_uop_ftq_idx : _GEN_190 ? _slots_4_io_uop_ftq_idx : _GEN_176 ? _slots_3_io_uop_ftq_idx : _GEN_162 ? _slots_2_io_uop_ftq_idx : _GEN_148 ? _slots_1_io_uop_ftq_idx : _GEN_141 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_0_edge_inst = _GEN_677 ? _slots_39_io_uop_edge_inst : _GEN_666 ? _slots_38_io_uop_edge_inst : _GEN_652 ? _slots_37_io_uop_edge_inst : _GEN_638 ? _slots_36_io_uop_edge_inst : _GEN_624 ? _slots_35_io_uop_edge_inst : _GEN_610 ? _slots_34_io_uop_edge_inst : _GEN_596 ? _slots_33_io_uop_edge_inst : _GEN_582 ? _slots_32_io_uop_edge_inst : _GEN_568 ? _slots_31_io_uop_edge_inst : _GEN_554 ? _slots_30_io_uop_edge_inst : _GEN_540 ? _slots_29_io_uop_edge_inst : _GEN_526 ? _slots_28_io_uop_edge_inst : _GEN_512 ? _slots_27_io_uop_edge_inst : _GEN_498 ? _slots_26_io_uop_edge_inst : _GEN_484 ? _slots_25_io_uop_edge_inst : _GEN_470 ? _slots_24_io_uop_edge_inst : _GEN_456 ? _slots_23_io_uop_edge_inst : _GEN_442 ? _slots_22_io_uop_edge_inst : _GEN_428 ? _slots_21_io_uop_edge_inst : _GEN_414 ? _slots_20_io_uop_edge_inst : _GEN_400 ? _slots_19_io_uop_edge_inst : _GEN_386 ? _slots_18_io_uop_edge_inst : _GEN_372 ? _slots_17_io_uop_edge_inst : _GEN_358 ? _slots_16_io_uop_edge_inst : _GEN_344 ? _slots_15_io_uop_edge_inst : _GEN_330 ? _slots_14_io_uop_edge_inst : _GEN_316 ? _slots_13_io_uop_edge_inst : _GEN_302 ? _slots_12_io_uop_edge_inst : _GEN_288 ? _slots_11_io_uop_edge_inst : _GEN_274 ? _slots_10_io_uop_edge_inst : _GEN_260 ? _slots_9_io_uop_edge_inst : _GEN_246 ? _slots_8_io_uop_edge_inst : _GEN_232 ? _slots_7_io_uop_edge_inst : _GEN_218 ? _slots_6_io_uop_edge_inst : _GEN_204 ? _slots_5_io_uop_edge_inst : _GEN_190 ? _slots_4_io_uop_edge_inst : _GEN_176 ? _slots_3_io_uop_edge_inst : _GEN_162 ? _slots_2_io_uop_edge_inst : _GEN_148 ? _slots_1_io_uop_edge_inst : _GEN_141 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_0_pc_lob = _GEN_677 ? _slots_39_io_uop_pc_lob : _GEN_666 ? _slots_38_io_uop_pc_lob : _GEN_652 ? _slots_37_io_uop_pc_lob : _GEN_638 ? _slots_36_io_uop_pc_lob : _GEN_624 ? _slots_35_io_uop_pc_lob : _GEN_610 ? _slots_34_io_uop_pc_lob : _GEN_596 ? _slots_33_io_uop_pc_lob : _GEN_582 ? _slots_32_io_uop_pc_lob : _GEN_568 ? _slots_31_io_uop_pc_lob : _GEN_554 ? _slots_30_io_uop_pc_lob : _GEN_540 ? _slots_29_io_uop_pc_lob : _GEN_526 ? _slots_28_io_uop_pc_lob : _GEN_512 ? _slots_27_io_uop_pc_lob : _GEN_498 ? _slots_26_io_uop_pc_lob : _GEN_484 ? _slots_25_io_uop_pc_lob : _GEN_470 ? _slots_24_io_uop_pc_lob : _GEN_456 ? _slots_23_io_uop_pc_lob : _GEN_442 ? _slots_22_io_uop_pc_lob : _GEN_428 ? _slots_21_io_uop_pc_lob : _GEN_414 ? _slots_20_io_uop_pc_lob : _GEN_400 ? _slots_19_io_uop_pc_lob : _GEN_386 ? _slots_18_io_uop_pc_lob : _GEN_372 ? _slots_17_io_uop_pc_lob : _GEN_358 ? _slots_16_io_uop_pc_lob : _GEN_344 ? _slots_15_io_uop_pc_lob : _GEN_330 ? _slots_14_io_uop_pc_lob : _GEN_316 ? _slots_13_io_uop_pc_lob : _GEN_302 ? _slots_12_io_uop_pc_lob : _GEN_288 ? _slots_11_io_uop_pc_lob : _GEN_274 ? _slots_10_io_uop_pc_lob : _GEN_260 ? _slots_9_io_uop_pc_lob : _GEN_246 ? _slots_8_io_uop_pc_lob : _GEN_232 ? _slots_7_io_uop_pc_lob : _GEN_218 ? _slots_6_io_uop_pc_lob : _GEN_204 ? _slots_5_io_uop_pc_lob : _GEN_190 ? _slots_4_io_uop_pc_lob : _GEN_176 ? _slots_3_io_uop_pc_lob : _GEN_162 ? _slots_2_io_uop_pc_lob : _GEN_148 ? _slots_1_io_uop_pc_lob : _GEN_141 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_0_taken = _GEN_677 ? _slots_39_io_uop_taken : _GEN_666 ? _slots_38_io_uop_taken : _GEN_652 ? _slots_37_io_uop_taken : _GEN_638 ? _slots_36_io_uop_taken : _GEN_624 ? _slots_35_io_uop_taken : _GEN_610 ? _slots_34_io_uop_taken : _GEN_596 ? _slots_33_io_uop_taken : _GEN_582 ? _slots_32_io_uop_taken : _GEN_568 ? _slots_31_io_uop_taken : _GEN_554 ? _slots_30_io_uop_taken : _GEN_540 ? _slots_29_io_uop_taken : _GEN_526 ? _slots_28_io_uop_taken : _GEN_512 ? _slots_27_io_uop_taken : _GEN_498 ? _slots_26_io_uop_taken : _GEN_484 ? _slots_25_io_uop_taken : _GEN_470 ? _slots_24_io_uop_taken : _GEN_456 ? _slots_23_io_uop_taken : _GEN_442 ? _slots_22_io_uop_taken : _GEN_428 ? _slots_21_io_uop_taken : _GEN_414 ? _slots_20_io_uop_taken : _GEN_400 ? _slots_19_io_uop_taken : _GEN_386 ? _slots_18_io_uop_taken : _GEN_372 ? _slots_17_io_uop_taken : _GEN_358 ? _slots_16_io_uop_taken : _GEN_344 ? _slots_15_io_uop_taken : _GEN_330 ? _slots_14_io_uop_taken : _GEN_316 ? _slots_13_io_uop_taken : _GEN_302 ? _slots_12_io_uop_taken : _GEN_288 ? _slots_11_io_uop_taken : _GEN_274 ? _slots_10_io_uop_taken : _GEN_260 ? _slots_9_io_uop_taken : _GEN_246 ? _slots_8_io_uop_taken : _GEN_232 ? _slots_7_io_uop_taken : _GEN_218 ? _slots_6_io_uop_taken : _GEN_204 ? _slots_5_io_uop_taken : _GEN_190 ? _slots_4_io_uop_taken : _GEN_176 ? _slots_3_io_uop_taken : _GEN_162 ? _slots_2_io_uop_taken : _GEN_148 ? _slots_1_io_uop_taken : _GEN_141 & _slots_0_io_uop_taken;
  assign io_iss_uops_0_imm_packed = _GEN_677 ? _slots_39_io_uop_imm_packed : _GEN_666 ? _slots_38_io_uop_imm_packed : _GEN_652 ? _slots_37_io_uop_imm_packed : _GEN_638 ? _slots_36_io_uop_imm_packed : _GEN_624 ? _slots_35_io_uop_imm_packed : _GEN_610 ? _slots_34_io_uop_imm_packed : _GEN_596 ? _slots_33_io_uop_imm_packed : _GEN_582 ? _slots_32_io_uop_imm_packed : _GEN_568 ? _slots_31_io_uop_imm_packed : _GEN_554 ? _slots_30_io_uop_imm_packed : _GEN_540 ? _slots_29_io_uop_imm_packed : _GEN_526 ? _slots_28_io_uop_imm_packed : _GEN_512 ? _slots_27_io_uop_imm_packed : _GEN_498 ? _slots_26_io_uop_imm_packed : _GEN_484 ? _slots_25_io_uop_imm_packed : _GEN_470 ? _slots_24_io_uop_imm_packed : _GEN_456 ? _slots_23_io_uop_imm_packed : _GEN_442 ? _slots_22_io_uop_imm_packed : _GEN_428 ? _slots_21_io_uop_imm_packed : _GEN_414 ? _slots_20_io_uop_imm_packed : _GEN_400 ? _slots_19_io_uop_imm_packed : _GEN_386 ? _slots_18_io_uop_imm_packed : _GEN_372 ? _slots_17_io_uop_imm_packed : _GEN_358 ? _slots_16_io_uop_imm_packed : _GEN_344 ? _slots_15_io_uop_imm_packed : _GEN_330 ? _slots_14_io_uop_imm_packed : _GEN_316 ? _slots_13_io_uop_imm_packed : _GEN_302 ? _slots_12_io_uop_imm_packed : _GEN_288 ? _slots_11_io_uop_imm_packed : _GEN_274 ? _slots_10_io_uop_imm_packed : _GEN_260 ? _slots_9_io_uop_imm_packed : _GEN_246 ? _slots_8_io_uop_imm_packed : _GEN_232 ? _slots_7_io_uop_imm_packed : _GEN_218 ? _slots_6_io_uop_imm_packed : _GEN_204 ? _slots_5_io_uop_imm_packed : _GEN_190 ? _slots_4_io_uop_imm_packed : _GEN_176 ? _slots_3_io_uop_imm_packed : _GEN_162 ? _slots_2_io_uop_imm_packed : _GEN_148 ? _slots_1_io_uop_imm_packed : _GEN_141 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_0_csr_addr = _GEN_677 ? _slots_39_io_uop_csr_addr : _GEN_666 ? _slots_38_io_uop_csr_addr : _GEN_652 ? _slots_37_io_uop_csr_addr : _GEN_638 ? _slots_36_io_uop_csr_addr : _GEN_624 ? _slots_35_io_uop_csr_addr : _GEN_610 ? _slots_34_io_uop_csr_addr : _GEN_596 ? _slots_33_io_uop_csr_addr : _GEN_582 ? _slots_32_io_uop_csr_addr : _GEN_568 ? _slots_31_io_uop_csr_addr : _GEN_554 ? _slots_30_io_uop_csr_addr : _GEN_540 ? _slots_29_io_uop_csr_addr : _GEN_526 ? _slots_28_io_uop_csr_addr : _GEN_512 ? _slots_27_io_uop_csr_addr : _GEN_498 ? _slots_26_io_uop_csr_addr : _GEN_484 ? _slots_25_io_uop_csr_addr : _GEN_470 ? _slots_24_io_uop_csr_addr : _GEN_456 ? _slots_23_io_uop_csr_addr : _GEN_442 ? _slots_22_io_uop_csr_addr : _GEN_428 ? _slots_21_io_uop_csr_addr : _GEN_414 ? _slots_20_io_uop_csr_addr : _GEN_400 ? _slots_19_io_uop_csr_addr : _GEN_386 ? _slots_18_io_uop_csr_addr : _GEN_372 ? _slots_17_io_uop_csr_addr : _GEN_358 ? _slots_16_io_uop_csr_addr : _GEN_344 ? _slots_15_io_uop_csr_addr : _GEN_330 ? _slots_14_io_uop_csr_addr : _GEN_316 ? _slots_13_io_uop_csr_addr : _GEN_302 ? _slots_12_io_uop_csr_addr : _GEN_288 ? _slots_11_io_uop_csr_addr : _GEN_274 ? _slots_10_io_uop_csr_addr : _GEN_260 ? _slots_9_io_uop_csr_addr : _GEN_246 ? _slots_8_io_uop_csr_addr : _GEN_232 ? _slots_7_io_uop_csr_addr : _GEN_218 ? _slots_6_io_uop_csr_addr : _GEN_204 ? _slots_5_io_uop_csr_addr : _GEN_190 ? _slots_4_io_uop_csr_addr : _GEN_176 ? _slots_3_io_uop_csr_addr : _GEN_162 ? _slots_2_io_uop_csr_addr : _GEN_148 ? _slots_1_io_uop_csr_addr : _GEN_141 ? _slots_0_io_uop_csr_addr : 12'h0;
  assign io_iss_uops_0_rob_idx = _GEN_677 ? _slots_39_io_uop_rob_idx : _GEN_666 ? _slots_38_io_uop_rob_idx : _GEN_652 ? _slots_37_io_uop_rob_idx : _GEN_638 ? _slots_36_io_uop_rob_idx : _GEN_624 ? _slots_35_io_uop_rob_idx : _GEN_610 ? _slots_34_io_uop_rob_idx : _GEN_596 ? _slots_33_io_uop_rob_idx : _GEN_582 ? _slots_32_io_uop_rob_idx : _GEN_568 ? _slots_31_io_uop_rob_idx : _GEN_554 ? _slots_30_io_uop_rob_idx : _GEN_540 ? _slots_29_io_uop_rob_idx : _GEN_526 ? _slots_28_io_uop_rob_idx : _GEN_512 ? _slots_27_io_uop_rob_idx : _GEN_498 ? _slots_26_io_uop_rob_idx : _GEN_484 ? _slots_25_io_uop_rob_idx : _GEN_470 ? _slots_24_io_uop_rob_idx : _GEN_456 ? _slots_23_io_uop_rob_idx : _GEN_442 ? _slots_22_io_uop_rob_idx : _GEN_428 ? _slots_21_io_uop_rob_idx : _GEN_414 ? _slots_20_io_uop_rob_idx : _GEN_400 ? _slots_19_io_uop_rob_idx : _GEN_386 ? _slots_18_io_uop_rob_idx : _GEN_372 ? _slots_17_io_uop_rob_idx : _GEN_358 ? _slots_16_io_uop_rob_idx : _GEN_344 ? _slots_15_io_uop_rob_idx : _GEN_330 ? _slots_14_io_uop_rob_idx : _GEN_316 ? _slots_13_io_uop_rob_idx : _GEN_302 ? _slots_12_io_uop_rob_idx : _GEN_288 ? _slots_11_io_uop_rob_idx : _GEN_274 ? _slots_10_io_uop_rob_idx : _GEN_260 ? _slots_9_io_uop_rob_idx : _GEN_246 ? _slots_8_io_uop_rob_idx : _GEN_232 ? _slots_7_io_uop_rob_idx : _GEN_218 ? _slots_6_io_uop_rob_idx : _GEN_204 ? _slots_5_io_uop_rob_idx : _GEN_190 ? _slots_4_io_uop_rob_idx : _GEN_176 ? _slots_3_io_uop_rob_idx : _GEN_162 ? _slots_2_io_uop_rob_idx : _GEN_148 ? _slots_1_io_uop_rob_idx : _GEN_141 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_0_ldq_idx = _GEN_677 ? _slots_39_io_uop_ldq_idx : _GEN_666 ? _slots_38_io_uop_ldq_idx : _GEN_652 ? _slots_37_io_uop_ldq_idx : _GEN_638 ? _slots_36_io_uop_ldq_idx : _GEN_624 ? _slots_35_io_uop_ldq_idx : _GEN_610 ? _slots_34_io_uop_ldq_idx : _GEN_596 ? _slots_33_io_uop_ldq_idx : _GEN_582 ? _slots_32_io_uop_ldq_idx : _GEN_568 ? _slots_31_io_uop_ldq_idx : _GEN_554 ? _slots_30_io_uop_ldq_idx : _GEN_540 ? _slots_29_io_uop_ldq_idx : _GEN_526 ? _slots_28_io_uop_ldq_idx : _GEN_512 ? _slots_27_io_uop_ldq_idx : _GEN_498 ? _slots_26_io_uop_ldq_idx : _GEN_484 ? _slots_25_io_uop_ldq_idx : _GEN_470 ? _slots_24_io_uop_ldq_idx : _GEN_456 ? _slots_23_io_uop_ldq_idx : _GEN_442 ? _slots_22_io_uop_ldq_idx : _GEN_428 ? _slots_21_io_uop_ldq_idx : _GEN_414 ? _slots_20_io_uop_ldq_idx : _GEN_400 ? _slots_19_io_uop_ldq_idx : _GEN_386 ? _slots_18_io_uop_ldq_idx : _GEN_372 ? _slots_17_io_uop_ldq_idx : _GEN_358 ? _slots_16_io_uop_ldq_idx : _GEN_344 ? _slots_15_io_uop_ldq_idx : _GEN_330 ? _slots_14_io_uop_ldq_idx : _GEN_316 ? _slots_13_io_uop_ldq_idx : _GEN_302 ? _slots_12_io_uop_ldq_idx : _GEN_288 ? _slots_11_io_uop_ldq_idx : _GEN_274 ? _slots_10_io_uop_ldq_idx : _GEN_260 ? _slots_9_io_uop_ldq_idx : _GEN_246 ? _slots_8_io_uop_ldq_idx : _GEN_232 ? _slots_7_io_uop_ldq_idx : _GEN_218 ? _slots_6_io_uop_ldq_idx : _GEN_204 ? _slots_5_io_uop_ldq_idx : _GEN_190 ? _slots_4_io_uop_ldq_idx : _GEN_176 ? _slots_3_io_uop_ldq_idx : _GEN_162 ? _slots_2_io_uop_ldq_idx : _GEN_148 ? _slots_1_io_uop_ldq_idx : _GEN_141 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_0_stq_idx = _GEN_677 ? _slots_39_io_uop_stq_idx : _GEN_666 ? _slots_38_io_uop_stq_idx : _GEN_652 ? _slots_37_io_uop_stq_idx : _GEN_638 ? _slots_36_io_uop_stq_idx : _GEN_624 ? _slots_35_io_uop_stq_idx : _GEN_610 ? _slots_34_io_uop_stq_idx : _GEN_596 ? _slots_33_io_uop_stq_idx : _GEN_582 ? _slots_32_io_uop_stq_idx : _GEN_568 ? _slots_31_io_uop_stq_idx : _GEN_554 ? _slots_30_io_uop_stq_idx : _GEN_540 ? _slots_29_io_uop_stq_idx : _GEN_526 ? _slots_28_io_uop_stq_idx : _GEN_512 ? _slots_27_io_uop_stq_idx : _GEN_498 ? _slots_26_io_uop_stq_idx : _GEN_484 ? _slots_25_io_uop_stq_idx : _GEN_470 ? _slots_24_io_uop_stq_idx : _GEN_456 ? _slots_23_io_uop_stq_idx : _GEN_442 ? _slots_22_io_uop_stq_idx : _GEN_428 ? _slots_21_io_uop_stq_idx : _GEN_414 ? _slots_20_io_uop_stq_idx : _GEN_400 ? _slots_19_io_uop_stq_idx : _GEN_386 ? _slots_18_io_uop_stq_idx : _GEN_372 ? _slots_17_io_uop_stq_idx : _GEN_358 ? _slots_16_io_uop_stq_idx : _GEN_344 ? _slots_15_io_uop_stq_idx : _GEN_330 ? _slots_14_io_uop_stq_idx : _GEN_316 ? _slots_13_io_uop_stq_idx : _GEN_302 ? _slots_12_io_uop_stq_idx : _GEN_288 ? _slots_11_io_uop_stq_idx : _GEN_274 ? _slots_10_io_uop_stq_idx : _GEN_260 ? _slots_9_io_uop_stq_idx : _GEN_246 ? _slots_8_io_uop_stq_idx : _GEN_232 ? _slots_7_io_uop_stq_idx : _GEN_218 ? _slots_6_io_uop_stq_idx : _GEN_204 ? _slots_5_io_uop_stq_idx : _GEN_190 ? _slots_4_io_uop_stq_idx : _GEN_176 ? _slots_3_io_uop_stq_idx : _GEN_162 ? _slots_2_io_uop_stq_idx : _GEN_148 ? _slots_1_io_uop_stq_idx : _GEN_141 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_0_rxq_idx = _GEN_677 ? _slots_39_io_uop_rxq_idx : _GEN_666 ? _slots_38_io_uop_rxq_idx : _GEN_652 ? _slots_37_io_uop_rxq_idx : _GEN_638 ? _slots_36_io_uop_rxq_idx : _GEN_624 ? _slots_35_io_uop_rxq_idx : _GEN_610 ? _slots_34_io_uop_rxq_idx : _GEN_596 ? _slots_33_io_uop_rxq_idx : _GEN_582 ? _slots_32_io_uop_rxq_idx : _GEN_568 ? _slots_31_io_uop_rxq_idx : _GEN_554 ? _slots_30_io_uop_rxq_idx : _GEN_540 ? _slots_29_io_uop_rxq_idx : _GEN_526 ? _slots_28_io_uop_rxq_idx : _GEN_512 ? _slots_27_io_uop_rxq_idx : _GEN_498 ? _slots_26_io_uop_rxq_idx : _GEN_484 ? _slots_25_io_uop_rxq_idx : _GEN_470 ? _slots_24_io_uop_rxq_idx : _GEN_456 ? _slots_23_io_uop_rxq_idx : _GEN_442 ? _slots_22_io_uop_rxq_idx : _GEN_428 ? _slots_21_io_uop_rxq_idx : _GEN_414 ? _slots_20_io_uop_rxq_idx : _GEN_400 ? _slots_19_io_uop_rxq_idx : _GEN_386 ? _slots_18_io_uop_rxq_idx : _GEN_372 ? _slots_17_io_uop_rxq_idx : _GEN_358 ? _slots_16_io_uop_rxq_idx : _GEN_344 ? _slots_15_io_uop_rxq_idx : _GEN_330 ? _slots_14_io_uop_rxq_idx : _GEN_316 ? _slots_13_io_uop_rxq_idx : _GEN_302 ? _slots_12_io_uop_rxq_idx : _GEN_288 ? _slots_11_io_uop_rxq_idx : _GEN_274 ? _slots_10_io_uop_rxq_idx : _GEN_260 ? _slots_9_io_uop_rxq_idx : _GEN_246 ? _slots_8_io_uop_rxq_idx : _GEN_232 ? _slots_7_io_uop_rxq_idx : _GEN_218 ? _slots_6_io_uop_rxq_idx : _GEN_204 ? _slots_5_io_uop_rxq_idx : _GEN_190 ? _slots_4_io_uop_rxq_idx : _GEN_176 ? _slots_3_io_uop_rxq_idx : _GEN_162 ? _slots_2_io_uop_rxq_idx : _GEN_148 ? _slots_1_io_uop_rxq_idx : _GEN_141 ? _slots_0_io_uop_rxq_idx : 2'h0;
  assign io_iss_uops_0_pdst = _GEN_677 ? _slots_39_io_uop_pdst : _GEN_666 ? _slots_38_io_uop_pdst : _GEN_652 ? _slots_37_io_uop_pdst : _GEN_638 ? _slots_36_io_uop_pdst : _GEN_624 ? _slots_35_io_uop_pdst : _GEN_610 ? _slots_34_io_uop_pdst : _GEN_596 ? _slots_33_io_uop_pdst : _GEN_582 ? _slots_32_io_uop_pdst : _GEN_568 ? _slots_31_io_uop_pdst : _GEN_554 ? _slots_30_io_uop_pdst : _GEN_540 ? _slots_29_io_uop_pdst : _GEN_526 ? _slots_28_io_uop_pdst : _GEN_512 ? _slots_27_io_uop_pdst : _GEN_498 ? _slots_26_io_uop_pdst : _GEN_484 ? _slots_25_io_uop_pdst : _GEN_470 ? _slots_24_io_uop_pdst : _GEN_456 ? _slots_23_io_uop_pdst : _GEN_442 ? _slots_22_io_uop_pdst : _GEN_428 ? _slots_21_io_uop_pdst : _GEN_414 ? _slots_20_io_uop_pdst : _GEN_400 ? _slots_19_io_uop_pdst : _GEN_386 ? _slots_18_io_uop_pdst : _GEN_372 ? _slots_17_io_uop_pdst : _GEN_358 ? _slots_16_io_uop_pdst : _GEN_344 ? _slots_15_io_uop_pdst : _GEN_330 ? _slots_14_io_uop_pdst : _GEN_316 ? _slots_13_io_uop_pdst : _GEN_302 ? _slots_12_io_uop_pdst : _GEN_288 ? _slots_11_io_uop_pdst : _GEN_274 ? _slots_10_io_uop_pdst : _GEN_260 ? _slots_9_io_uop_pdst : _GEN_246 ? _slots_8_io_uop_pdst : _GEN_232 ? _slots_7_io_uop_pdst : _GEN_218 ? _slots_6_io_uop_pdst : _GEN_204 ? _slots_5_io_uop_pdst : _GEN_190 ? _slots_4_io_uop_pdst : _GEN_176 ? _slots_3_io_uop_pdst : _GEN_162 ? _slots_2_io_uop_pdst : _GEN_148 ? _slots_1_io_uop_pdst : _GEN_141 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_0_prs1 = _GEN_677 ? _slots_39_io_uop_prs1 : _GEN_666 ? _slots_38_io_uop_prs1 : _GEN_652 ? _slots_37_io_uop_prs1 : _GEN_638 ? _slots_36_io_uop_prs1 : _GEN_624 ? _slots_35_io_uop_prs1 : _GEN_610 ? _slots_34_io_uop_prs1 : _GEN_596 ? _slots_33_io_uop_prs1 : _GEN_582 ? _slots_32_io_uop_prs1 : _GEN_568 ? _slots_31_io_uop_prs1 : _GEN_554 ? _slots_30_io_uop_prs1 : _GEN_540 ? _slots_29_io_uop_prs1 : _GEN_526 ? _slots_28_io_uop_prs1 : _GEN_512 ? _slots_27_io_uop_prs1 : _GEN_498 ? _slots_26_io_uop_prs1 : _GEN_484 ? _slots_25_io_uop_prs1 : _GEN_470 ? _slots_24_io_uop_prs1 : _GEN_456 ? _slots_23_io_uop_prs1 : _GEN_442 ? _slots_22_io_uop_prs1 : _GEN_428 ? _slots_21_io_uop_prs1 : _GEN_414 ? _slots_20_io_uop_prs1 : _GEN_400 ? _slots_19_io_uop_prs1 : _GEN_386 ? _slots_18_io_uop_prs1 : _GEN_372 ? _slots_17_io_uop_prs1 : _GEN_358 ? _slots_16_io_uop_prs1 : _GEN_344 ? _slots_15_io_uop_prs1 : _GEN_330 ? _slots_14_io_uop_prs1 : _GEN_316 ? _slots_13_io_uop_prs1 : _GEN_302 ? _slots_12_io_uop_prs1 : _GEN_288 ? _slots_11_io_uop_prs1 : _GEN_274 ? _slots_10_io_uop_prs1 : _GEN_260 ? _slots_9_io_uop_prs1 : _GEN_246 ? _slots_8_io_uop_prs1 : _GEN_232 ? _slots_7_io_uop_prs1 : _GEN_218 ? _slots_6_io_uop_prs1 : _GEN_204 ? _slots_5_io_uop_prs1 : _GEN_190 ? _slots_4_io_uop_prs1 : _GEN_176 ? _slots_3_io_uop_prs1 : _GEN_162 ? _slots_2_io_uop_prs1 : _GEN_148 ? _slots_1_io_uop_prs1 : _GEN_141 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_0_prs2 = _GEN_677 ? _slots_39_io_uop_prs2 : _GEN_666 ? _slots_38_io_uop_prs2 : _GEN_652 ? _slots_37_io_uop_prs2 : _GEN_638 ? _slots_36_io_uop_prs2 : _GEN_624 ? _slots_35_io_uop_prs2 : _GEN_610 ? _slots_34_io_uop_prs2 : _GEN_596 ? _slots_33_io_uop_prs2 : _GEN_582 ? _slots_32_io_uop_prs2 : _GEN_568 ? _slots_31_io_uop_prs2 : _GEN_554 ? _slots_30_io_uop_prs2 : _GEN_540 ? _slots_29_io_uop_prs2 : _GEN_526 ? _slots_28_io_uop_prs2 : _GEN_512 ? _slots_27_io_uop_prs2 : _GEN_498 ? _slots_26_io_uop_prs2 : _GEN_484 ? _slots_25_io_uop_prs2 : _GEN_470 ? _slots_24_io_uop_prs2 : _GEN_456 ? _slots_23_io_uop_prs2 : _GEN_442 ? _slots_22_io_uop_prs2 : _GEN_428 ? _slots_21_io_uop_prs2 : _GEN_414 ? _slots_20_io_uop_prs2 : _GEN_400 ? _slots_19_io_uop_prs2 : _GEN_386 ? _slots_18_io_uop_prs2 : _GEN_372 ? _slots_17_io_uop_prs2 : _GEN_358 ? _slots_16_io_uop_prs2 : _GEN_344 ? _slots_15_io_uop_prs2 : _GEN_330 ? _slots_14_io_uop_prs2 : _GEN_316 ? _slots_13_io_uop_prs2 : _GEN_302 ? _slots_12_io_uop_prs2 : _GEN_288 ? _slots_11_io_uop_prs2 : _GEN_274 ? _slots_10_io_uop_prs2 : _GEN_260 ? _slots_9_io_uop_prs2 : _GEN_246 ? _slots_8_io_uop_prs2 : _GEN_232 ? _slots_7_io_uop_prs2 : _GEN_218 ? _slots_6_io_uop_prs2 : _GEN_204 ? _slots_5_io_uop_prs2 : _GEN_190 ? _slots_4_io_uop_prs2 : _GEN_176 ? _slots_3_io_uop_prs2 : _GEN_162 ? _slots_2_io_uop_prs2 : _GEN_148 ? _slots_1_io_uop_prs2 : _GEN_141 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_0_prs3 = _GEN_677 ? _slots_39_io_uop_prs3 : _GEN_666 ? _slots_38_io_uop_prs3 : _GEN_652 ? _slots_37_io_uop_prs3 : _GEN_638 ? _slots_36_io_uop_prs3 : _GEN_624 ? _slots_35_io_uop_prs3 : _GEN_610 ? _slots_34_io_uop_prs3 : _GEN_596 ? _slots_33_io_uop_prs3 : _GEN_582 ? _slots_32_io_uop_prs3 : _GEN_568 ? _slots_31_io_uop_prs3 : _GEN_554 ? _slots_30_io_uop_prs3 : _GEN_540 ? _slots_29_io_uop_prs3 : _GEN_526 ? _slots_28_io_uop_prs3 : _GEN_512 ? _slots_27_io_uop_prs3 : _GEN_498 ? _slots_26_io_uop_prs3 : _GEN_484 ? _slots_25_io_uop_prs3 : _GEN_470 ? _slots_24_io_uop_prs3 : _GEN_456 ? _slots_23_io_uop_prs3 : _GEN_442 ? _slots_22_io_uop_prs3 : _GEN_428 ? _slots_21_io_uop_prs3 : _GEN_414 ? _slots_20_io_uop_prs3 : _GEN_400 ? _slots_19_io_uop_prs3 : _GEN_386 ? _slots_18_io_uop_prs3 : _GEN_372 ? _slots_17_io_uop_prs3 : _GEN_358 ? _slots_16_io_uop_prs3 : _GEN_344 ? _slots_15_io_uop_prs3 : _GEN_330 ? _slots_14_io_uop_prs3 : _GEN_316 ? _slots_13_io_uop_prs3 : _GEN_302 ? _slots_12_io_uop_prs3 : _GEN_288 ? _slots_11_io_uop_prs3 : _GEN_274 ? _slots_10_io_uop_prs3 : _GEN_260 ? _slots_9_io_uop_prs3 : _GEN_246 ? _slots_8_io_uop_prs3 : _GEN_232 ? _slots_7_io_uop_prs3 : _GEN_218 ? _slots_6_io_uop_prs3 : _GEN_204 ? _slots_5_io_uop_prs3 : _GEN_190 ? _slots_4_io_uop_prs3 : _GEN_176 ? _slots_3_io_uop_prs3 : _GEN_162 ? _slots_2_io_uop_prs3 : _GEN_148 ? _slots_1_io_uop_prs3 : _GEN_141 ? _slots_0_io_uop_prs3 : 7'h0;
  assign io_iss_uops_0_ppred = _GEN_677 ? _slots_39_io_uop_ppred : _GEN_666 ? _slots_38_io_uop_ppred : _GEN_652 ? _slots_37_io_uop_ppred : _GEN_638 ? _slots_36_io_uop_ppred : _GEN_624 ? _slots_35_io_uop_ppred : _GEN_610 ? _slots_34_io_uop_ppred : _GEN_596 ? _slots_33_io_uop_ppred : _GEN_582 ? _slots_32_io_uop_ppred : _GEN_568 ? _slots_31_io_uop_ppred : _GEN_554 ? _slots_30_io_uop_ppred : _GEN_540 ? _slots_29_io_uop_ppred : _GEN_526 ? _slots_28_io_uop_ppred : _GEN_512 ? _slots_27_io_uop_ppred : _GEN_498 ? _slots_26_io_uop_ppred : _GEN_484 ? _slots_25_io_uop_ppred : _GEN_470 ? _slots_24_io_uop_ppred : _GEN_456 ? _slots_23_io_uop_ppred : _GEN_442 ? _slots_22_io_uop_ppred : _GEN_428 ? _slots_21_io_uop_ppred : _GEN_414 ? _slots_20_io_uop_ppred : _GEN_400 ? _slots_19_io_uop_ppred : _GEN_386 ? _slots_18_io_uop_ppred : _GEN_372 ? _slots_17_io_uop_ppred : _GEN_358 ? _slots_16_io_uop_ppred : _GEN_344 ? _slots_15_io_uop_ppred : _GEN_330 ? _slots_14_io_uop_ppred : _GEN_316 ? _slots_13_io_uop_ppred : _GEN_302 ? _slots_12_io_uop_ppred : _GEN_288 ? _slots_11_io_uop_ppred : _GEN_274 ? _slots_10_io_uop_ppred : _GEN_260 ? _slots_9_io_uop_ppred : _GEN_246 ? _slots_8_io_uop_ppred : _GEN_232 ? _slots_7_io_uop_ppred : _GEN_218 ? _slots_6_io_uop_ppred : _GEN_204 ? _slots_5_io_uop_ppred : _GEN_190 ? _slots_4_io_uop_ppred : _GEN_176 ? _slots_3_io_uop_ppred : _GEN_162 ? _slots_2_io_uop_ppred : _GEN_148 ? _slots_1_io_uop_ppred : _GEN_141 ? _slots_0_io_uop_ppred : 6'h0;
  assign io_iss_uops_0_prs1_busy = _GEN_677 ? _slots_39_io_uop_prs1_busy : _GEN_666 ? _slots_38_io_uop_prs1_busy : _GEN_652 ? _slots_37_io_uop_prs1_busy : _GEN_638 ? _slots_36_io_uop_prs1_busy : _GEN_624 ? _slots_35_io_uop_prs1_busy : _GEN_610 ? _slots_34_io_uop_prs1_busy : _GEN_596 ? _slots_33_io_uop_prs1_busy : _GEN_582 ? _slots_32_io_uop_prs1_busy : _GEN_568 ? _slots_31_io_uop_prs1_busy : _GEN_554 ? _slots_30_io_uop_prs1_busy : _GEN_540 ? _slots_29_io_uop_prs1_busy : _GEN_526 ? _slots_28_io_uop_prs1_busy : _GEN_512 ? _slots_27_io_uop_prs1_busy : _GEN_498 ? _slots_26_io_uop_prs1_busy : _GEN_484 ? _slots_25_io_uop_prs1_busy : _GEN_470 ? _slots_24_io_uop_prs1_busy : _GEN_456 ? _slots_23_io_uop_prs1_busy : _GEN_442 ? _slots_22_io_uop_prs1_busy : _GEN_428 ? _slots_21_io_uop_prs1_busy : _GEN_414 ? _slots_20_io_uop_prs1_busy : _GEN_400 ? _slots_19_io_uop_prs1_busy : _GEN_386 ? _slots_18_io_uop_prs1_busy : _GEN_372 ? _slots_17_io_uop_prs1_busy : _GEN_358 ? _slots_16_io_uop_prs1_busy : _GEN_344 ? _slots_15_io_uop_prs1_busy : _GEN_330 ? _slots_14_io_uop_prs1_busy : _GEN_316 ? _slots_13_io_uop_prs1_busy : _GEN_302 ? _slots_12_io_uop_prs1_busy : _GEN_288 ? _slots_11_io_uop_prs1_busy : _GEN_274 ? _slots_10_io_uop_prs1_busy : _GEN_260 ? _slots_9_io_uop_prs1_busy : _GEN_246 ? _slots_8_io_uop_prs1_busy : _GEN_232 ? _slots_7_io_uop_prs1_busy : _GEN_218 ? _slots_6_io_uop_prs1_busy : _GEN_204 ? _slots_5_io_uop_prs1_busy : _GEN_190 ? _slots_4_io_uop_prs1_busy : _GEN_176 ? _slots_3_io_uop_prs1_busy : _GEN_162 ? _slots_2_io_uop_prs1_busy : _GEN_148 ? _slots_1_io_uop_prs1_busy : _GEN_141 & _slots_0_io_uop_prs1_busy;
  assign io_iss_uops_0_prs2_busy = _GEN_677 ? _slots_39_io_uop_prs2_busy : _GEN_666 ? _slots_38_io_uop_prs2_busy : _GEN_652 ? _slots_37_io_uop_prs2_busy : _GEN_638 ? _slots_36_io_uop_prs2_busy : _GEN_624 ? _slots_35_io_uop_prs2_busy : _GEN_610 ? _slots_34_io_uop_prs2_busy : _GEN_596 ? _slots_33_io_uop_prs2_busy : _GEN_582 ? _slots_32_io_uop_prs2_busy : _GEN_568 ? _slots_31_io_uop_prs2_busy : _GEN_554 ? _slots_30_io_uop_prs2_busy : _GEN_540 ? _slots_29_io_uop_prs2_busy : _GEN_526 ? _slots_28_io_uop_prs2_busy : _GEN_512 ? _slots_27_io_uop_prs2_busy : _GEN_498 ? _slots_26_io_uop_prs2_busy : _GEN_484 ? _slots_25_io_uop_prs2_busy : _GEN_470 ? _slots_24_io_uop_prs2_busy : _GEN_456 ? _slots_23_io_uop_prs2_busy : _GEN_442 ? _slots_22_io_uop_prs2_busy : _GEN_428 ? _slots_21_io_uop_prs2_busy : _GEN_414 ? _slots_20_io_uop_prs2_busy : _GEN_400 ? _slots_19_io_uop_prs2_busy : _GEN_386 ? _slots_18_io_uop_prs2_busy : _GEN_372 ? _slots_17_io_uop_prs2_busy : _GEN_358 ? _slots_16_io_uop_prs2_busy : _GEN_344 ? _slots_15_io_uop_prs2_busy : _GEN_330 ? _slots_14_io_uop_prs2_busy : _GEN_316 ? _slots_13_io_uop_prs2_busy : _GEN_302 ? _slots_12_io_uop_prs2_busy : _GEN_288 ? _slots_11_io_uop_prs2_busy : _GEN_274 ? _slots_10_io_uop_prs2_busy : _GEN_260 ? _slots_9_io_uop_prs2_busy : _GEN_246 ? _slots_8_io_uop_prs2_busy : _GEN_232 ? _slots_7_io_uop_prs2_busy : _GEN_218 ? _slots_6_io_uop_prs2_busy : _GEN_204 ? _slots_5_io_uop_prs2_busy : _GEN_190 ? _slots_4_io_uop_prs2_busy : _GEN_176 ? _slots_3_io_uop_prs2_busy : _GEN_162 ? _slots_2_io_uop_prs2_busy : _GEN_148 ? _slots_1_io_uop_prs2_busy : _GEN_141 & _slots_0_io_uop_prs2_busy;
  assign io_iss_uops_0_prs3_busy = _GEN_677 ? _slots_39_io_uop_prs3_busy : _GEN_666 ? _slots_38_io_uop_prs3_busy : _GEN_652 ? _slots_37_io_uop_prs3_busy : _GEN_638 ? _slots_36_io_uop_prs3_busy : _GEN_624 ? _slots_35_io_uop_prs3_busy : _GEN_610 ? _slots_34_io_uop_prs3_busy : _GEN_596 ? _slots_33_io_uop_prs3_busy : _GEN_582 ? _slots_32_io_uop_prs3_busy : _GEN_568 ? _slots_31_io_uop_prs3_busy : _GEN_554 ? _slots_30_io_uop_prs3_busy : _GEN_540 ? _slots_29_io_uop_prs3_busy : _GEN_526 ? _slots_28_io_uop_prs3_busy : _GEN_512 ? _slots_27_io_uop_prs3_busy : _GEN_498 ? _slots_26_io_uop_prs3_busy : _GEN_484 ? _slots_25_io_uop_prs3_busy : _GEN_470 ? _slots_24_io_uop_prs3_busy : _GEN_456 ? _slots_23_io_uop_prs3_busy : _GEN_442 ? _slots_22_io_uop_prs3_busy : _GEN_428 ? _slots_21_io_uop_prs3_busy : _GEN_414 ? _slots_20_io_uop_prs3_busy : _GEN_400 ? _slots_19_io_uop_prs3_busy : _GEN_386 ? _slots_18_io_uop_prs3_busy : _GEN_372 ? _slots_17_io_uop_prs3_busy : _GEN_358 ? _slots_16_io_uop_prs3_busy : _GEN_344 ? _slots_15_io_uop_prs3_busy : _GEN_330 ? _slots_14_io_uop_prs3_busy : _GEN_316 ? _slots_13_io_uop_prs3_busy : _GEN_302 ? _slots_12_io_uop_prs3_busy : _GEN_288 ? _slots_11_io_uop_prs3_busy : _GEN_274 ? _slots_10_io_uop_prs3_busy : _GEN_260 ? _slots_9_io_uop_prs3_busy : _GEN_246 ? _slots_8_io_uop_prs3_busy : _GEN_232 ? _slots_7_io_uop_prs3_busy : _GEN_218 ? _slots_6_io_uop_prs3_busy : _GEN_204 ? _slots_5_io_uop_prs3_busy : _GEN_190 ? _slots_4_io_uop_prs3_busy : _GEN_176 ? _slots_3_io_uop_prs3_busy : _GEN_162 ? _slots_2_io_uop_prs3_busy : _GEN_148 ? _slots_1_io_uop_prs3_busy : _GEN_141 & _slots_0_io_uop_prs3_busy;
  assign io_iss_uops_0_ppred_busy = _GEN_677 ? _slots_39_io_uop_ppred_busy : _GEN_666 ? _slots_38_io_uop_ppred_busy : _GEN_652 ? _slots_37_io_uop_ppred_busy : _GEN_638 ? _slots_36_io_uop_ppred_busy : _GEN_624 ? _slots_35_io_uop_ppred_busy : _GEN_610 ? _slots_34_io_uop_ppred_busy : _GEN_596 ? _slots_33_io_uop_ppred_busy : _GEN_582 ? _slots_32_io_uop_ppred_busy : _GEN_568 ? _slots_31_io_uop_ppred_busy : _GEN_554 ? _slots_30_io_uop_ppred_busy : _GEN_540 ? _slots_29_io_uop_ppred_busy : _GEN_526 ? _slots_28_io_uop_ppred_busy : _GEN_512 ? _slots_27_io_uop_ppred_busy : _GEN_498 ? _slots_26_io_uop_ppred_busy : _GEN_484 ? _slots_25_io_uop_ppred_busy : _GEN_470 ? _slots_24_io_uop_ppred_busy : _GEN_456 ? _slots_23_io_uop_ppred_busy : _GEN_442 ? _slots_22_io_uop_ppred_busy : _GEN_428 ? _slots_21_io_uop_ppred_busy : _GEN_414 ? _slots_20_io_uop_ppred_busy : _GEN_400 ? _slots_19_io_uop_ppred_busy : _GEN_386 ? _slots_18_io_uop_ppred_busy : _GEN_372 ? _slots_17_io_uop_ppred_busy : _GEN_358 ? _slots_16_io_uop_ppred_busy : _GEN_344 ? _slots_15_io_uop_ppred_busy : _GEN_330 ? _slots_14_io_uop_ppred_busy : _GEN_316 ? _slots_13_io_uop_ppred_busy : _GEN_302 ? _slots_12_io_uop_ppred_busy : _GEN_288 ? _slots_11_io_uop_ppred_busy : _GEN_274 ? _slots_10_io_uop_ppred_busy : _GEN_260 ? _slots_9_io_uop_ppred_busy : _GEN_246 ? _slots_8_io_uop_ppred_busy : _GEN_232 ? _slots_7_io_uop_ppred_busy : _GEN_218 ? _slots_6_io_uop_ppred_busy : _GEN_204 ? _slots_5_io_uop_ppred_busy : _GEN_190 ? _slots_4_io_uop_ppred_busy : _GEN_176 ? _slots_3_io_uop_ppred_busy : _GEN_162 ? _slots_2_io_uop_ppred_busy : _GEN_148 ? _slots_1_io_uop_ppred_busy : _GEN_141 & _slots_0_io_uop_ppred_busy;
  assign io_iss_uops_0_stale_pdst = _GEN_677 ? _slots_39_io_uop_stale_pdst : _GEN_666 ? _slots_38_io_uop_stale_pdst : _GEN_652 ? _slots_37_io_uop_stale_pdst : _GEN_638 ? _slots_36_io_uop_stale_pdst : _GEN_624 ? _slots_35_io_uop_stale_pdst : _GEN_610 ? _slots_34_io_uop_stale_pdst : _GEN_596 ? _slots_33_io_uop_stale_pdst : _GEN_582 ? _slots_32_io_uop_stale_pdst : _GEN_568 ? _slots_31_io_uop_stale_pdst : _GEN_554 ? _slots_30_io_uop_stale_pdst : _GEN_540 ? _slots_29_io_uop_stale_pdst : _GEN_526 ? _slots_28_io_uop_stale_pdst : _GEN_512 ? _slots_27_io_uop_stale_pdst : _GEN_498 ? _slots_26_io_uop_stale_pdst : _GEN_484 ? _slots_25_io_uop_stale_pdst : _GEN_470 ? _slots_24_io_uop_stale_pdst : _GEN_456 ? _slots_23_io_uop_stale_pdst : _GEN_442 ? _slots_22_io_uop_stale_pdst : _GEN_428 ? _slots_21_io_uop_stale_pdst : _GEN_414 ? _slots_20_io_uop_stale_pdst : _GEN_400 ? _slots_19_io_uop_stale_pdst : _GEN_386 ? _slots_18_io_uop_stale_pdst : _GEN_372 ? _slots_17_io_uop_stale_pdst : _GEN_358 ? _slots_16_io_uop_stale_pdst : _GEN_344 ? _slots_15_io_uop_stale_pdst : _GEN_330 ? _slots_14_io_uop_stale_pdst : _GEN_316 ? _slots_13_io_uop_stale_pdst : _GEN_302 ? _slots_12_io_uop_stale_pdst : _GEN_288 ? _slots_11_io_uop_stale_pdst : _GEN_274 ? _slots_10_io_uop_stale_pdst : _GEN_260 ? _slots_9_io_uop_stale_pdst : _GEN_246 ? _slots_8_io_uop_stale_pdst : _GEN_232 ? _slots_7_io_uop_stale_pdst : _GEN_218 ? _slots_6_io_uop_stale_pdst : _GEN_204 ? _slots_5_io_uop_stale_pdst : _GEN_190 ? _slots_4_io_uop_stale_pdst : _GEN_176 ? _slots_3_io_uop_stale_pdst : _GEN_162 ? _slots_2_io_uop_stale_pdst : _GEN_148 ? _slots_1_io_uop_stale_pdst : _GEN_141 ? _slots_0_io_uop_stale_pdst : 7'h0;
  assign io_iss_uops_0_exception = _GEN_677 ? _slots_39_io_uop_exception : _GEN_666 ? _slots_38_io_uop_exception : _GEN_652 ? _slots_37_io_uop_exception : _GEN_638 ? _slots_36_io_uop_exception : _GEN_624 ? _slots_35_io_uop_exception : _GEN_610 ? _slots_34_io_uop_exception : _GEN_596 ? _slots_33_io_uop_exception : _GEN_582 ? _slots_32_io_uop_exception : _GEN_568 ? _slots_31_io_uop_exception : _GEN_554 ? _slots_30_io_uop_exception : _GEN_540 ? _slots_29_io_uop_exception : _GEN_526 ? _slots_28_io_uop_exception : _GEN_512 ? _slots_27_io_uop_exception : _GEN_498 ? _slots_26_io_uop_exception : _GEN_484 ? _slots_25_io_uop_exception : _GEN_470 ? _slots_24_io_uop_exception : _GEN_456 ? _slots_23_io_uop_exception : _GEN_442 ? _slots_22_io_uop_exception : _GEN_428 ? _slots_21_io_uop_exception : _GEN_414 ? _slots_20_io_uop_exception : _GEN_400 ? _slots_19_io_uop_exception : _GEN_386 ? _slots_18_io_uop_exception : _GEN_372 ? _slots_17_io_uop_exception : _GEN_358 ? _slots_16_io_uop_exception : _GEN_344 ? _slots_15_io_uop_exception : _GEN_330 ? _slots_14_io_uop_exception : _GEN_316 ? _slots_13_io_uop_exception : _GEN_302 ? _slots_12_io_uop_exception : _GEN_288 ? _slots_11_io_uop_exception : _GEN_274 ? _slots_10_io_uop_exception : _GEN_260 ? _slots_9_io_uop_exception : _GEN_246 ? _slots_8_io_uop_exception : _GEN_232 ? _slots_7_io_uop_exception : _GEN_218 ? _slots_6_io_uop_exception : _GEN_204 ? _slots_5_io_uop_exception : _GEN_190 ? _slots_4_io_uop_exception : _GEN_176 ? _slots_3_io_uop_exception : _GEN_162 ? _slots_2_io_uop_exception : _GEN_148 ? _slots_1_io_uop_exception : _GEN_141 & _slots_0_io_uop_exception;
  assign io_iss_uops_0_exc_cause = _GEN_677 ? _slots_39_io_uop_exc_cause : _GEN_666 ? _slots_38_io_uop_exc_cause : _GEN_652 ? _slots_37_io_uop_exc_cause : _GEN_638 ? _slots_36_io_uop_exc_cause : _GEN_624 ? _slots_35_io_uop_exc_cause : _GEN_610 ? _slots_34_io_uop_exc_cause : _GEN_596 ? _slots_33_io_uop_exc_cause : _GEN_582 ? _slots_32_io_uop_exc_cause : _GEN_568 ? _slots_31_io_uop_exc_cause : _GEN_554 ? _slots_30_io_uop_exc_cause : _GEN_540 ? _slots_29_io_uop_exc_cause : _GEN_526 ? _slots_28_io_uop_exc_cause : _GEN_512 ? _slots_27_io_uop_exc_cause : _GEN_498 ? _slots_26_io_uop_exc_cause : _GEN_484 ? _slots_25_io_uop_exc_cause : _GEN_470 ? _slots_24_io_uop_exc_cause : _GEN_456 ? _slots_23_io_uop_exc_cause : _GEN_442 ? _slots_22_io_uop_exc_cause : _GEN_428 ? _slots_21_io_uop_exc_cause : _GEN_414 ? _slots_20_io_uop_exc_cause : _GEN_400 ? _slots_19_io_uop_exc_cause : _GEN_386 ? _slots_18_io_uop_exc_cause : _GEN_372 ? _slots_17_io_uop_exc_cause : _GEN_358 ? _slots_16_io_uop_exc_cause : _GEN_344 ? _slots_15_io_uop_exc_cause : _GEN_330 ? _slots_14_io_uop_exc_cause : _GEN_316 ? _slots_13_io_uop_exc_cause : _GEN_302 ? _slots_12_io_uop_exc_cause : _GEN_288 ? _slots_11_io_uop_exc_cause : _GEN_274 ? _slots_10_io_uop_exc_cause : _GEN_260 ? _slots_9_io_uop_exc_cause : _GEN_246 ? _slots_8_io_uop_exc_cause : _GEN_232 ? _slots_7_io_uop_exc_cause : _GEN_218 ? _slots_6_io_uop_exc_cause : _GEN_204 ? _slots_5_io_uop_exc_cause : _GEN_190 ? _slots_4_io_uop_exc_cause : _GEN_176 ? _slots_3_io_uop_exc_cause : _GEN_162 ? _slots_2_io_uop_exc_cause : _GEN_148 ? _slots_1_io_uop_exc_cause : _GEN_141 ? _slots_0_io_uop_exc_cause : 64'h0;
  assign io_iss_uops_0_bypassable = _GEN_677 ? _slots_39_io_uop_bypassable : _GEN_666 ? _slots_38_io_uop_bypassable : _GEN_652 ? _slots_37_io_uop_bypassable : _GEN_638 ? _slots_36_io_uop_bypassable : _GEN_624 ? _slots_35_io_uop_bypassable : _GEN_610 ? _slots_34_io_uop_bypassable : _GEN_596 ? _slots_33_io_uop_bypassable : _GEN_582 ? _slots_32_io_uop_bypassable : _GEN_568 ? _slots_31_io_uop_bypassable : _GEN_554 ? _slots_30_io_uop_bypassable : _GEN_540 ? _slots_29_io_uop_bypassable : _GEN_526 ? _slots_28_io_uop_bypassable : _GEN_512 ? _slots_27_io_uop_bypassable : _GEN_498 ? _slots_26_io_uop_bypassable : _GEN_484 ? _slots_25_io_uop_bypassable : _GEN_470 ? _slots_24_io_uop_bypassable : _GEN_456 ? _slots_23_io_uop_bypassable : _GEN_442 ? _slots_22_io_uop_bypassable : _GEN_428 ? _slots_21_io_uop_bypassable : _GEN_414 ? _slots_20_io_uop_bypassable : _GEN_400 ? _slots_19_io_uop_bypassable : _GEN_386 ? _slots_18_io_uop_bypassable : _GEN_372 ? _slots_17_io_uop_bypassable : _GEN_358 ? _slots_16_io_uop_bypassable : _GEN_344 ? _slots_15_io_uop_bypassable : _GEN_330 ? _slots_14_io_uop_bypassable : _GEN_316 ? _slots_13_io_uop_bypassable : _GEN_302 ? _slots_12_io_uop_bypassable : _GEN_288 ? _slots_11_io_uop_bypassable : _GEN_274 ? _slots_10_io_uop_bypassable : _GEN_260 ? _slots_9_io_uop_bypassable : _GEN_246 ? _slots_8_io_uop_bypassable : _GEN_232 ? _slots_7_io_uop_bypassable : _GEN_218 ? _slots_6_io_uop_bypassable : _GEN_204 ? _slots_5_io_uop_bypassable : _GEN_190 ? _slots_4_io_uop_bypassable : _GEN_176 ? _slots_3_io_uop_bypassable : _GEN_162 ? _slots_2_io_uop_bypassable : _GEN_148 ? _slots_1_io_uop_bypassable : _GEN_141 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_0_mem_cmd = _GEN_677 ? _slots_39_io_uop_mem_cmd : _GEN_666 ? _slots_38_io_uop_mem_cmd : _GEN_652 ? _slots_37_io_uop_mem_cmd : _GEN_638 ? _slots_36_io_uop_mem_cmd : _GEN_624 ? _slots_35_io_uop_mem_cmd : _GEN_610 ? _slots_34_io_uop_mem_cmd : _GEN_596 ? _slots_33_io_uop_mem_cmd : _GEN_582 ? _slots_32_io_uop_mem_cmd : _GEN_568 ? _slots_31_io_uop_mem_cmd : _GEN_554 ? _slots_30_io_uop_mem_cmd : _GEN_540 ? _slots_29_io_uop_mem_cmd : _GEN_526 ? _slots_28_io_uop_mem_cmd : _GEN_512 ? _slots_27_io_uop_mem_cmd : _GEN_498 ? _slots_26_io_uop_mem_cmd : _GEN_484 ? _slots_25_io_uop_mem_cmd : _GEN_470 ? _slots_24_io_uop_mem_cmd : _GEN_456 ? _slots_23_io_uop_mem_cmd : _GEN_442 ? _slots_22_io_uop_mem_cmd : _GEN_428 ? _slots_21_io_uop_mem_cmd : _GEN_414 ? _slots_20_io_uop_mem_cmd : _GEN_400 ? _slots_19_io_uop_mem_cmd : _GEN_386 ? _slots_18_io_uop_mem_cmd : _GEN_372 ? _slots_17_io_uop_mem_cmd : _GEN_358 ? _slots_16_io_uop_mem_cmd : _GEN_344 ? _slots_15_io_uop_mem_cmd : _GEN_330 ? _slots_14_io_uop_mem_cmd : _GEN_316 ? _slots_13_io_uop_mem_cmd : _GEN_302 ? _slots_12_io_uop_mem_cmd : _GEN_288 ? _slots_11_io_uop_mem_cmd : _GEN_274 ? _slots_10_io_uop_mem_cmd : _GEN_260 ? _slots_9_io_uop_mem_cmd : _GEN_246 ? _slots_8_io_uop_mem_cmd : _GEN_232 ? _slots_7_io_uop_mem_cmd : _GEN_218 ? _slots_6_io_uop_mem_cmd : _GEN_204 ? _slots_5_io_uop_mem_cmd : _GEN_190 ? _slots_4_io_uop_mem_cmd : _GEN_176 ? _slots_3_io_uop_mem_cmd : _GEN_162 ? _slots_2_io_uop_mem_cmd : _GEN_148 ? _slots_1_io_uop_mem_cmd : _GEN_141 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_0_mem_size = _GEN_677 ? _slots_39_io_uop_mem_size : _GEN_666 ? _slots_38_io_uop_mem_size : _GEN_652 ? _slots_37_io_uop_mem_size : _GEN_638 ? _slots_36_io_uop_mem_size : _GEN_624 ? _slots_35_io_uop_mem_size : _GEN_610 ? _slots_34_io_uop_mem_size : _GEN_596 ? _slots_33_io_uop_mem_size : _GEN_582 ? _slots_32_io_uop_mem_size : _GEN_568 ? _slots_31_io_uop_mem_size : _GEN_554 ? _slots_30_io_uop_mem_size : _GEN_540 ? _slots_29_io_uop_mem_size : _GEN_526 ? _slots_28_io_uop_mem_size : _GEN_512 ? _slots_27_io_uop_mem_size : _GEN_498 ? _slots_26_io_uop_mem_size : _GEN_484 ? _slots_25_io_uop_mem_size : _GEN_470 ? _slots_24_io_uop_mem_size : _GEN_456 ? _slots_23_io_uop_mem_size : _GEN_442 ? _slots_22_io_uop_mem_size : _GEN_428 ? _slots_21_io_uop_mem_size : _GEN_414 ? _slots_20_io_uop_mem_size : _GEN_400 ? _slots_19_io_uop_mem_size : _GEN_386 ? _slots_18_io_uop_mem_size : _GEN_372 ? _slots_17_io_uop_mem_size : _GEN_358 ? _slots_16_io_uop_mem_size : _GEN_344 ? _slots_15_io_uop_mem_size : _GEN_330 ? _slots_14_io_uop_mem_size : _GEN_316 ? _slots_13_io_uop_mem_size : _GEN_302 ? _slots_12_io_uop_mem_size : _GEN_288 ? _slots_11_io_uop_mem_size : _GEN_274 ? _slots_10_io_uop_mem_size : _GEN_260 ? _slots_9_io_uop_mem_size : _GEN_246 ? _slots_8_io_uop_mem_size : _GEN_232 ? _slots_7_io_uop_mem_size : _GEN_218 ? _slots_6_io_uop_mem_size : _GEN_204 ? _slots_5_io_uop_mem_size : _GEN_190 ? _slots_4_io_uop_mem_size : _GEN_176 ? _slots_3_io_uop_mem_size : _GEN_162 ? _slots_2_io_uop_mem_size : _GEN_148 ? _slots_1_io_uop_mem_size : _GEN_141 ? _slots_0_io_uop_mem_size : 2'h0;
  assign io_iss_uops_0_mem_signed = _GEN_677 ? _slots_39_io_uop_mem_signed : _GEN_666 ? _slots_38_io_uop_mem_signed : _GEN_652 ? _slots_37_io_uop_mem_signed : _GEN_638 ? _slots_36_io_uop_mem_signed : _GEN_624 ? _slots_35_io_uop_mem_signed : _GEN_610 ? _slots_34_io_uop_mem_signed : _GEN_596 ? _slots_33_io_uop_mem_signed : _GEN_582 ? _slots_32_io_uop_mem_signed : _GEN_568 ? _slots_31_io_uop_mem_signed : _GEN_554 ? _slots_30_io_uop_mem_signed : _GEN_540 ? _slots_29_io_uop_mem_signed : _GEN_526 ? _slots_28_io_uop_mem_signed : _GEN_512 ? _slots_27_io_uop_mem_signed : _GEN_498 ? _slots_26_io_uop_mem_signed : _GEN_484 ? _slots_25_io_uop_mem_signed : _GEN_470 ? _slots_24_io_uop_mem_signed : _GEN_456 ? _slots_23_io_uop_mem_signed : _GEN_442 ? _slots_22_io_uop_mem_signed : _GEN_428 ? _slots_21_io_uop_mem_signed : _GEN_414 ? _slots_20_io_uop_mem_signed : _GEN_400 ? _slots_19_io_uop_mem_signed : _GEN_386 ? _slots_18_io_uop_mem_signed : _GEN_372 ? _slots_17_io_uop_mem_signed : _GEN_358 ? _slots_16_io_uop_mem_signed : _GEN_344 ? _slots_15_io_uop_mem_signed : _GEN_330 ? _slots_14_io_uop_mem_signed : _GEN_316 ? _slots_13_io_uop_mem_signed : _GEN_302 ? _slots_12_io_uop_mem_signed : _GEN_288 ? _slots_11_io_uop_mem_signed : _GEN_274 ? _slots_10_io_uop_mem_signed : _GEN_260 ? _slots_9_io_uop_mem_signed : _GEN_246 ? _slots_8_io_uop_mem_signed : _GEN_232 ? _slots_7_io_uop_mem_signed : _GEN_218 ? _slots_6_io_uop_mem_signed : _GEN_204 ? _slots_5_io_uop_mem_signed : _GEN_190 ? _slots_4_io_uop_mem_signed : _GEN_176 ? _slots_3_io_uop_mem_signed : _GEN_162 ? _slots_2_io_uop_mem_signed : _GEN_148 ? _slots_1_io_uop_mem_signed : _GEN_141 & _slots_0_io_uop_mem_signed;
  assign io_iss_uops_0_is_fence = _GEN_677 ? _slots_39_io_uop_is_fence : _GEN_666 ? _slots_38_io_uop_is_fence : _GEN_652 ? _slots_37_io_uop_is_fence : _GEN_638 ? _slots_36_io_uop_is_fence : _GEN_624 ? _slots_35_io_uop_is_fence : _GEN_610 ? _slots_34_io_uop_is_fence : _GEN_596 ? _slots_33_io_uop_is_fence : _GEN_582 ? _slots_32_io_uop_is_fence : _GEN_568 ? _slots_31_io_uop_is_fence : _GEN_554 ? _slots_30_io_uop_is_fence : _GEN_540 ? _slots_29_io_uop_is_fence : _GEN_526 ? _slots_28_io_uop_is_fence : _GEN_512 ? _slots_27_io_uop_is_fence : _GEN_498 ? _slots_26_io_uop_is_fence : _GEN_484 ? _slots_25_io_uop_is_fence : _GEN_470 ? _slots_24_io_uop_is_fence : _GEN_456 ? _slots_23_io_uop_is_fence : _GEN_442 ? _slots_22_io_uop_is_fence : _GEN_428 ? _slots_21_io_uop_is_fence : _GEN_414 ? _slots_20_io_uop_is_fence : _GEN_400 ? _slots_19_io_uop_is_fence : _GEN_386 ? _slots_18_io_uop_is_fence : _GEN_372 ? _slots_17_io_uop_is_fence : _GEN_358 ? _slots_16_io_uop_is_fence : _GEN_344 ? _slots_15_io_uop_is_fence : _GEN_330 ? _slots_14_io_uop_is_fence : _GEN_316 ? _slots_13_io_uop_is_fence : _GEN_302 ? _slots_12_io_uop_is_fence : _GEN_288 ? _slots_11_io_uop_is_fence : _GEN_274 ? _slots_10_io_uop_is_fence : _GEN_260 ? _slots_9_io_uop_is_fence : _GEN_246 ? _slots_8_io_uop_is_fence : _GEN_232 ? _slots_7_io_uop_is_fence : _GEN_218 ? _slots_6_io_uop_is_fence : _GEN_204 ? _slots_5_io_uop_is_fence : _GEN_190 ? _slots_4_io_uop_is_fence : _GEN_176 ? _slots_3_io_uop_is_fence : _GEN_162 ? _slots_2_io_uop_is_fence : _GEN_148 ? _slots_1_io_uop_is_fence : _GEN_141 & _slots_0_io_uop_is_fence;
  assign io_iss_uops_0_is_fencei = _GEN_677 ? _slots_39_io_uop_is_fencei : _GEN_666 ? _slots_38_io_uop_is_fencei : _GEN_652 ? _slots_37_io_uop_is_fencei : _GEN_638 ? _slots_36_io_uop_is_fencei : _GEN_624 ? _slots_35_io_uop_is_fencei : _GEN_610 ? _slots_34_io_uop_is_fencei : _GEN_596 ? _slots_33_io_uop_is_fencei : _GEN_582 ? _slots_32_io_uop_is_fencei : _GEN_568 ? _slots_31_io_uop_is_fencei : _GEN_554 ? _slots_30_io_uop_is_fencei : _GEN_540 ? _slots_29_io_uop_is_fencei : _GEN_526 ? _slots_28_io_uop_is_fencei : _GEN_512 ? _slots_27_io_uop_is_fencei : _GEN_498 ? _slots_26_io_uop_is_fencei : _GEN_484 ? _slots_25_io_uop_is_fencei : _GEN_470 ? _slots_24_io_uop_is_fencei : _GEN_456 ? _slots_23_io_uop_is_fencei : _GEN_442 ? _slots_22_io_uop_is_fencei : _GEN_428 ? _slots_21_io_uop_is_fencei : _GEN_414 ? _slots_20_io_uop_is_fencei : _GEN_400 ? _slots_19_io_uop_is_fencei : _GEN_386 ? _slots_18_io_uop_is_fencei : _GEN_372 ? _slots_17_io_uop_is_fencei : _GEN_358 ? _slots_16_io_uop_is_fencei : _GEN_344 ? _slots_15_io_uop_is_fencei : _GEN_330 ? _slots_14_io_uop_is_fencei : _GEN_316 ? _slots_13_io_uop_is_fencei : _GEN_302 ? _slots_12_io_uop_is_fencei : _GEN_288 ? _slots_11_io_uop_is_fencei : _GEN_274 ? _slots_10_io_uop_is_fencei : _GEN_260 ? _slots_9_io_uop_is_fencei : _GEN_246 ? _slots_8_io_uop_is_fencei : _GEN_232 ? _slots_7_io_uop_is_fencei : _GEN_218 ? _slots_6_io_uop_is_fencei : _GEN_204 ? _slots_5_io_uop_is_fencei : _GEN_190 ? _slots_4_io_uop_is_fencei : _GEN_176 ? _slots_3_io_uop_is_fencei : _GEN_162 ? _slots_2_io_uop_is_fencei : _GEN_148 ? _slots_1_io_uop_is_fencei : _GEN_141 & _slots_0_io_uop_is_fencei;
  assign io_iss_uops_0_is_amo = _GEN_677 ? _slots_39_io_uop_is_amo : _GEN_666 ? _slots_38_io_uop_is_amo : _GEN_652 ? _slots_37_io_uop_is_amo : _GEN_638 ? _slots_36_io_uop_is_amo : _GEN_624 ? _slots_35_io_uop_is_amo : _GEN_610 ? _slots_34_io_uop_is_amo : _GEN_596 ? _slots_33_io_uop_is_amo : _GEN_582 ? _slots_32_io_uop_is_amo : _GEN_568 ? _slots_31_io_uop_is_amo : _GEN_554 ? _slots_30_io_uop_is_amo : _GEN_540 ? _slots_29_io_uop_is_amo : _GEN_526 ? _slots_28_io_uop_is_amo : _GEN_512 ? _slots_27_io_uop_is_amo : _GEN_498 ? _slots_26_io_uop_is_amo : _GEN_484 ? _slots_25_io_uop_is_amo : _GEN_470 ? _slots_24_io_uop_is_amo : _GEN_456 ? _slots_23_io_uop_is_amo : _GEN_442 ? _slots_22_io_uop_is_amo : _GEN_428 ? _slots_21_io_uop_is_amo : _GEN_414 ? _slots_20_io_uop_is_amo : _GEN_400 ? _slots_19_io_uop_is_amo : _GEN_386 ? _slots_18_io_uop_is_amo : _GEN_372 ? _slots_17_io_uop_is_amo : _GEN_358 ? _slots_16_io_uop_is_amo : _GEN_344 ? _slots_15_io_uop_is_amo : _GEN_330 ? _slots_14_io_uop_is_amo : _GEN_316 ? _slots_13_io_uop_is_amo : _GEN_302 ? _slots_12_io_uop_is_amo : _GEN_288 ? _slots_11_io_uop_is_amo : _GEN_274 ? _slots_10_io_uop_is_amo : _GEN_260 ? _slots_9_io_uop_is_amo : _GEN_246 ? _slots_8_io_uop_is_amo : _GEN_232 ? _slots_7_io_uop_is_amo : _GEN_218 ? _slots_6_io_uop_is_amo : _GEN_204 ? _slots_5_io_uop_is_amo : _GEN_190 ? _slots_4_io_uop_is_amo : _GEN_176 ? _slots_3_io_uop_is_amo : _GEN_162 ? _slots_2_io_uop_is_amo : _GEN_148 ? _slots_1_io_uop_is_amo : _GEN_141 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_0_uses_ldq = _GEN_677 ? _slots_39_io_uop_uses_ldq : _GEN_666 ? _slots_38_io_uop_uses_ldq : _GEN_652 ? _slots_37_io_uop_uses_ldq : _GEN_638 ? _slots_36_io_uop_uses_ldq : _GEN_624 ? _slots_35_io_uop_uses_ldq : _GEN_610 ? _slots_34_io_uop_uses_ldq : _GEN_596 ? _slots_33_io_uop_uses_ldq : _GEN_582 ? _slots_32_io_uop_uses_ldq : _GEN_568 ? _slots_31_io_uop_uses_ldq : _GEN_554 ? _slots_30_io_uop_uses_ldq : _GEN_540 ? _slots_29_io_uop_uses_ldq : _GEN_526 ? _slots_28_io_uop_uses_ldq : _GEN_512 ? _slots_27_io_uop_uses_ldq : _GEN_498 ? _slots_26_io_uop_uses_ldq : _GEN_484 ? _slots_25_io_uop_uses_ldq : _GEN_470 ? _slots_24_io_uop_uses_ldq : _GEN_456 ? _slots_23_io_uop_uses_ldq : _GEN_442 ? _slots_22_io_uop_uses_ldq : _GEN_428 ? _slots_21_io_uop_uses_ldq : _GEN_414 ? _slots_20_io_uop_uses_ldq : _GEN_400 ? _slots_19_io_uop_uses_ldq : _GEN_386 ? _slots_18_io_uop_uses_ldq : _GEN_372 ? _slots_17_io_uop_uses_ldq : _GEN_358 ? _slots_16_io_uop_uses_ldq : _GEN_344 ? _slots_15_io_uop_uses_ldq : _GEN_330 ? _slots_14_io_uop_uses_ldq : _GEN_316 ? _slots_13_io_uop_uses_ldq : _GEN_302 ? _slots_12_io_uop_uses_ldq : _GEN_288 ? _slots_11_io_uop_uses_ldq : _GEN_274 ? _slots_10_io_uop_uses_ldq : _GEN_260 ? _slots_9_io_uop_uses_ldq : _GEN_246 ? _slots_8_io_uop_uses_ldq : _GEN_232 ? _slots_7_io_uop_uses_ldq : _GEN_218 ? _slots_6_io_uop_uses_ldq : _GEN_204 ? _slots_5_io_uop_uses_ldq : _GEN_190 ? _slots_4_io_uop_uses_ldq : _GEN_176 ? _slots_3_io_uop_uses_ldq : _GEN_162 ? _slots_2_io_uop_uses_ldq : _GEN_148 ? _slots_1_io_uop_uses_ldq : _GEN_141 & _slots_0_io_uop_uses_ldq;
  assign io_iss_uops_0_uses_stq = _GEN_677 ? _slots_39_io_uop_uses_stq : _GEN_666 ? _slots_38_io_uop_uses_stq : _GEN_652 ? _slots_37_io_uop_uses_stq : _GEN_638 ? _slots_36_io_uop_uses_stq : _GEN_624 ? _slots_35_io_uop_uses_stq : _GEN_610 ? _slots_34_io_uop_uses_stq : _GEN_596 ? _slots_33_io_uop_uses_stq : _GEN_582 ? _slots_32_io_uop_uses_stq : _GEN_568 ? _slots_31_io_uop_uses_stq : _GEN_554 ? _slots_30_io_uop_uses_stq : _GEN_540 ? _slots_29_io_uop_uses_stq : _GEN_526 ? _slots_28_io_uop_uses_stq : _GEN_512 ? _slots_27_io_uop_uses_stq : _GEN_498 ? _slots_26_io_uop_uses_stq : _GEN_484 ? _slots_25_io_uop_uses_stq : _GEN_470 ? _slots_24_io_uop_uses_stq : _GEN_456 ? _slots_23_io_uop_uses_stq : _GEN_442 ? _slots_22_io_uop_uses_stq : _GEN_428 ? _slots_21_io_uop_uses_stq : _GEN_414 ? _slots_20_io_uop_uses_stq : _GEN_400 ? _slots_19_io_uop_uses_stq : _GEN_386 ? _slots_18_io_uop_uses_stq : _GEN_372 ? _slots_17_io_uop_uses_stq : _GEN_358 ? _slots_16_io_uop_uses_stq : _GEN_344 ? _slots_15_io_uop_uses_stq : _GEN_330 ? _slots_14_io_uop_uses_stq : _GEN_316 ? _slots_13_io_uop_uses_stq : _GEN_302 ? _slots_12_io_uop_uses_stq : _GEN_288 ? _slots_11_io_uop_uses_stq : _GEN_274 ? _slots_10_io_uop_uses_stq : _GEN_260 ? _slots_9_io_uop_uses_stq : _GEN_246 ? _slots_8_io_uop_uses_stq : _GEN_232 ? _slots_7_io_uop_uses_stq : _GEN_218 ? _slots_6_io_uop_uses_stq : _GEN_204 ? _slots_5_io_uop_uses_stq : _GEN_190 ? _slots_4_io_uop_uses_stq : _GEN_176 ? _slots_3_io_uop_uses_stq : _GEN_162 ? _slots_2_io_uop_uses_stq : _GEN_148 ? _slots_1_io_uop_uses_stq : _GEN_141 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_0_is_sys_pc2epc = _GEN_677 ? _slots_39_io_uop_is_sys_pc2epc : _GEN_666 ? _slots_38_io_uop_is_sys_pc2epc : _GEN_652 ? _slots_37_io_uop_is_sys_pc2epc : _GEN_638 ? _slots_36_io_uop_is_sys_pc2epc : _GEN_624 ? _slots_35_io_uop_is_sys_pc2epc : _GEN_610 ? _slots_34_io_uop_is_sys_pc2epc : _GEN_596 ? _slots_33_io_uop_is_sys_pc2epc : _GEN_582 ? _slots_32_io_uop_is_sys_pc2epc : _GEN_568 ? _slots_31_io_uop_is_sys_pc2epc : _GEN_554 ? _slots_30_io_uop_is_sys_pc2epc : _GEN_540 ? _slots_29_io_uop_is_sys_pc2epc : _GEN_526 ? _slots_28_io_uop_is_sys_pc2epc : _GEN_512 ? _slots_27_io_uop_is_sys_pc2epc : _GEN_498 ? _slots_26_io_uop_is_sys_pc2epc : _GEN_484 ? _slots_25_io_uop_is_sys_pc2epc : _GEN_470 ? _slots_24_io_uop_is_sys_pc2epc : _GEN_456 ? _slots_23_io_uop_is_sys_pc2epc : _GEN_442 ? _slots_22_io_uop_is_sys_pc2epc : _GEN_428 ? _slots_21_io_uop_is_sys_pc2epc : _GEN_414 ? _slots_20_io_uop_is_sys_pc2epc : _GEN_400 ? _slots_19_io_uop_is_sys_pc2epc : _GEN_386 ? _slots_18_io_uop_is_sys_pc2epc : _GEN_372 ? _slots_17_io_uop_is_sys_pc2epc : _GEN_358 ? _slots_16_io_uop_is_sys_pc2epc : _GEN_344 ? _slots_15_io_uop_is_sys_pc2epc : _GEN_330 ? _slots_14_io_uop_is_sys_pc2epc : _GEN_316 ? _slots_13_io_uop_is_sys_pc2epc : _GEN_302 ? _slots_12_io_uop_is_sys_pc2epc : _GEN_288 ? _slots_11_io_uop_is_sys_pc2epc : _GEN_274 ? _slots_10_io_uop_is_sys_pc2epc : _GEN_260 ? _slots_9_io_uop_is_sys_pc2epc : _GEN_246 ? _slots_8_io_uop_is_sys_pc2epc : _GEN_232 ? _slots_7_io_uop_is_sys_pc2epc : _GEN_218 ? _slots_6_io_uop_is_sys_pc2epc : _GEN_204 ? _slots_5_io_uop_is_sys_pc2epc : _GEN_190 ? _slots_4_io_uop_is_sys_pc2epc : _GEN_176 ? _slots_3_io_uop_is_sys_pc2epc : _GEN_162 ? _slots_2_io_uop_is_sys_pc2epc : _GEN_148 ? _slots_1_io_uop_is_sys_pc2epc : _GEN_141 & _slots_0_io_uop_is_sys_pc2epc;
  assign io_iss_uops_0_is_unique = _GEN_677 ? _slots_39_io_uop_is_unique : _GEN_666 ? _slots_38_io_uop_is_unique : _GEN_652 ? _slots_37_io_uop_is_unique : _GEN_638 ? _slots_36_io_uop_is_unique : _GEN_624 ? _slots_35_io_uop_is_unique : _GEN_610 ? _slots_34_io_uop_is_unique : _GEN_596 ? _slots_33_io_uop_is_unique : _GEN_582 ? _slots_32_io_uop_is_unique : _GEN_568 ? _slots_31_io_uop_is_unique : _GEN_554 ? _slots_30_io_uop_is_unique : _GEN_540 ? _slots_29_io_uop_is_unique : _GEN_526 ? _slots_28_io_uop_is_unique : _GEN_512 ? _slots_27_io_uop_is_unique : _GEN_498 ? _slots_26_io_uop_is_unique : _GEN_484 ? _slots_25_io_uop_is_unique : _GEN_470 ? _slots_24_io_uop_is_unique : _GEN_456 ? _slots_23_io_uop_is_unique : _GEN_442 ? _slots_22_io_uop_is_unique : _GEN_428 ? _slots_21_io_uop_is_unique : _GEN_414 ? _slots_20_io_uop_is_unique : _GEN_400 ? _slots_19_io_uop_is_unique : _GEN_386 ? _slots_18_io_uop_is_unique : _GEN_372 ? _slots_17_io_uop_is_unique : _GEN_358 ? _slots_16_io_uop_is_unique : _GEN_344 ? _slots_15_io_uop_is_unique : _GEN_330 ? _slots_14_io_uop_is_unique : _GEN_316 ? _slots_13_io_uop_is_unique : _GEN_302 ? _slots_12_io_uop_is_unique : _GEN_288 ? _slots_11_io_uop_is_unique : _GEN_274 ? _slots_10_io_uop_is_unique : _GEN_260 ? _slots_9_io_uop_is_unique : _GEN_246 ? _slots_8_io_uop_is_unique : _GEN_232 ? _slots_7_io_uop_is_unique : _GEN_218 ? _slots_6_io_uop_is_unique : _GEN_204 ? _slots_5_io_uop_is_unique : _GEN_190 ? _slots_4_io_uop_is_unique : _GEN_176 ? _slots_3_io_uop_is_unique : _GEN_162 ? _slots_2_io_uop_is_unique : _GEN_148 ? _slots_1_io_uop_is_unique : _GEN_141 & _slots_0_io_uop_is_unique;
  assign io_iss_uops_0_flush_on_commit = _GEN_677 ? _slots_39_io_uop_flush_on_commit : _GEN_666 ? _slots_38_io_uop_flush_on_commit : _GEN_652 ? _slots_37_io_uop_flush_on_commit : _GEN_638 ? _slots_36_io_uop_flush_on_commit : _GEN_624 ? _slots_35_io_uop_flush_on_commit : _GEN_610 ? _slots_34_io_uop_flush_on_commit : _GEN_596 ? _slots_33_io_uop_flush_on_commit : _GEN_582 ? _slots_32_io_uop_flush_on_commit : _GEN_568 ? _slots_31_io_uop_flush_on_commit : _GEN_554 ? _slots_30_io_uop_flush_on_commit : _GEN_540 ? _slots_29_io_uop_flush_on_commit : _GEN_526 ? _slots_28_io_uop_flush_on_commit : _GEN_512 ? _slots_27_io_uop_flush_on_commit : _GEN_498 ? _slots_26_io_uop_flush_on_commit : _GEN_484 ? _slots_25_io_uop_flush_on_commit : _GEN_470 ? _slots_24_io_uop_flush_on_commit : _GEN_456 ? _slots_23_io_uop_flush_on_commit : _GEN_442 ? _slots_22_io_uop_flush_on_commit : _GEN_428 ? _slots_21_io_uop_flush_on_commit : _GEN_414 ? _slots_20_io_uop_flush_on_commit : _GEN_400 ? _slots_19_io_uop_flush_on_commit : _GEN_386 ? _slots_18_io_uop_flush_on_commit : _GEN_372 ? _slots_17_io_uop_flush_on_commit : _GEN_358 ? _slots_16_io_uop_flush_on_commit : _GEN_344 ? _slots_15_io_uop_flush_on_commit : _GEN_330 ? _slots_14_io_uop_flush_on_commit : _GEN_316 ? _slots_13_io_uop_flush_on_commit : _GEN_302 ? _slots_12_io_uop_flush_on_commit : _GEN_288 ? _slots_11_io_uop_flush_on_commit : _GEN_274 ? _slots_10_io_uop_flush_on_commit : _GEN_260 ? _slots_9_io_uop_flush_on_commit : _GEN_246 ? _slots_8_io_uop_flush_on_commit : _GEN_232 ? _slots_7_io_uop_flush_on_commit : _GEN_218 ? _slots_6_io_uop_flush_on_commit : _GEN_204 ? _slots_5_io_uop_flush_on_commit : _GEN_190 ? _slots_4_io_uop_flush_on_commit : _GEN_176 ? _slots_3_io_uop_flush_on_commit : _GEN_162 ? _slots_2_io_uop_flush_on_commit : _GEN_148 ? _slots_1_io_uop_flush_on_commit : _GEN_141 & _slots_0_io_uop_flush_on_commit;
  assign io_iss_uops_0_ldst_is_rs1 = _GEN_677 ? _slots_39_io_uop_ldst_is_rs1 : _GEN_666 ? _slots_38_io_uop_ldst_is_rs1 : _GEN_652 ? _slots_37_io_uop_ldst_is_rs1 : _GEN_638 ? _slots_36_io_uop_ldst_is_rs1 : _GEN_624 ? _slots_35_io_uop_ldst_is_rs1 : _GEN_610 ? _slots_34_io_uop_ldst_is_rs1 : _GEN_596 ? _slots_33_io_uop_ldst_is_rs1 : _GEN_582 ? _slots_32_io_uop_ldst_is_rs1 : _GEN_568 ? _slots_31_io_uop_ldst_is_rs1 : _GEN_554 ? _slots_30_io_uop_ldst_is_rs1 : _GEN_540 ? _slots_29_io_uop_ldst_is_rs1 : _GEN_526 ? _slots_28_io_uop_ldst_is_rs1 : _GEN_512 ? _slots_27_io_uop_ldst_is_rs1 : _GEN_498 ? _slots_26_io_uop_ldst_is_rs1 : _GEN_484 ? _slots_25_io_uop_ldst_is_rs1 : _GEN_470 ? _slots_24_io_uop_ldst_is_rs1 : _GEN_456 ? _slots_23_io_uop_ldst_is_rs1 : _GEN_442 ? _slots_22_io_uop_ldst_is_rs1 : _GEN_428 ? _slots_21_io_uop_ldst_is_rs1 : _GEN_414 ? _slots_20_io_uop_ldst_is_rs1 : _GEN_400 ? _slots_19_io_uop_ldst_is_rs1 : _GEN_386 ? _slots_18_io_uop_ldst_is_rs1 : _GEN_372 ? _slots_17_io_uop_ldst_is_rs1 : _GEN_358 ? _slots_16_io_uop_ldst_is_rs1 : _GEN_344 ? _slots_15_io_uop_ldst_is_rs1 : _GEN_330 ? _slots_14_io_uop_ldst_is_rs1 : _GEN_316 ? _slots_13_io_uop_ldst_is_rs1 : _GEN_302 ? _slots_12_io_uop_ldst_is_rs1 : _GEN_288 ? _slots_11_io_uop_ldst_is_rs1 : _GEN_274 ? _slots_10_io_uop_ldst_is_rs1 : _GEN_260 ? _slots_9_io_uop_ldst_is_rs1 : _GEN_246 ? _slots_8_io_uop_ldst_is_rs1 : _GEN_232 ? _slots_7_io_uop_ldst_is_rs1 : _GEN_218 ? _slots_6_io_uop_ldst_is_rs1 : _GEN_204 ? _slots_5_io_uop_ldst_is_rs1 : _GEN_190 ? _slots_4_io_uop_ldst_is_rs1 : _GEN_176 ? _slots_3_io_uop_ldst_is_rs1 : _GEN_162 ? _slots_2_io_uop_ldst_is_rs1 : _GEN_148 ? _slots_1_io_uop_ldst_is_rs1 : _GEN_141 & _slots_0_io_uop_ldst_is_rs1;
  assign io_iss_uops_0_ldst = _GEN_677 ? _slots_39_io_uop_ldst : _GEN_666 ? _slots_38_io_uop_ldst : _GEN_652 ? _slots_37_io_uop_ldst : _GEN_638 ? _slots_36_io_uop_ldst : _GEN_624 ? _slots_35_io_uop_ldst : _GEN_610 ? _slots_34_io_uop_ldst : _GEN_596 ? _slots_33_io_uop_ldst : _GEN_582 ? _slots_32_io_uop_ldst : _GEN_568 ? _slots_31_io_uop_ldst : _GEN_554 ? _slots_30_io_uop_ldst : _GEN_540 ? _slots_29_io_uop_ldst : _GEN_526 ? _slots_28_io_uop_ldst : _GEN_512 ? _slots_27_io_uop_ldst : _GEN_498 ? _slots_26_io_uop_ldst : _GEN_484 ? _slots_25_io_uop_ldst : _GEN_470 ? _slots_24_io_uop_ldst : _GEN_456 ? _slots_23_io_uop_ldst : _GEN_442 ? _slots_22_io_uop_ldst : _GEN_428 ? _slots_21_io_uop_ldst : _GEN_414 ? _slots_20_io_uop_ldst : _GEN_400 ? _slots_19_io_uop_ldst : _GEN_386 ? _slots_18_io_uop_ldst : _GEN_372 ? _slots_17_io_uop_ldst : _GEN_358 ? _slots_16_io_uop_ldst : _GEN_344 ? _slots_15_io_uop_ldst : _GEN_330 ? _slots_14_io_uop_ldst : _GEN_316 ? _slots_13_io_uop_ldst : _GEN_302 ? _slots_12_io_uop_ldst : _GEN_288 ? _slots_11_io_uop_ldst : _GEN_274 ? _slots_10_io_uop_ldst : _GEN_260 ? _slots_9_io_uop_ldst : _GEN_246 ? _slots_8_io_uop_ldst : _GEN_232 ? _slots_7_io_uop_ldst : _GEN_218 ? _slots_6_io_uop_ldst : _GEN_204 ? _slots_5_io_uop_ldst : _GEN_190 ? _slots_4_io_uop_ldst : _GEN_176 ? _slots_3_io_uop_ldst : _GEN_162 ? _slots_2_io_uop_ldst : _GEN_148 ? _slots_1_io_uop_ldst : _GEN_141 ? _slots_0_io_uop_ldst : 6'h0;
  assign io_iss_uops_0_lrs1 = _GEN_677 ? _slots_39_io_uop_lrs1 : _GEN_666 ? _slots_38_io_uop_lrs1 : _GEN_652 ? _slots_37_io_uop_lrs1 : _GEN_638 ? _slots_36_io_uop_lrs1 : _GEN_624 ? _slots_35_io_uop_lrs1 : _GEN_610 ? _slots_34_io_uop_lrs1 : _GEN_596 ? _slots_33_io_uop_lrs1 : _GEN_582 ? _slots_32_io_uop_lrs1 : _GEN_568 ? _slots_31_io_uop_lrs1 : _GEN_554 ? _slots_30_io_uop_lrs1 : _GEN_540 ? _slots_29_io_uop_lrs1 : _GEN_526 ? _slots_28_io_uop_lrs1 : _GEN_512 ? _slots_27_io_uop_lrs1 : _GEN_498 ? _slots_26_io_uop_lrs1 : _GEN_484 ? _slots_25_io_uop_lrs1 : _GEN_470 ? _slots_24_io_uop_lrs1 : _GEN_456 ? _slots_23_io_uop_lrs1 : _GEN_442 ? _slots_22_io_uop_lrs1 : _GEN_428 ? _slots_21_io_uop_lrs1 : _GEN_414 ? _slots_20_io_uop_lrs1 : _GEN_400 ? _slots_19_io_uop_lrs1 : _GEN_386 ? _slots_18_io_uop_lrs1 : _GEN_372 ? _slots_17_io_uop_lrs1 : _GEN_358 ? _slots_16_io_uop_lrs1 : _GEN_344 ? _slots_15_io_uop_lrs1 : _GEN_330 ? _slots_14_io_uop_lrs1 : _GEN_316 ? _slots_13_io_uop_lrs1 : _GEN_302 ? _slots_12_io_uop_lrs1 : _GEN_288 ? _slots_11_io_uop_lrs1 : _GEN_274 ? _slots_10_io_uop_lrs1 : _GEN_260 ? _slots_9_io_uop_lrs1 : _GEN_246 ? _slots_8_io_uop_lrs1 : _GEN_232 ? _slots_7_io_uop_lrs1 : _GEN_218 ? _slots_6_io_uop_lrs1 : _GEN_204 ? _slots_5_io_uop_lrs1 : _GEN_190 ? _slots_4_io_uop_lrs1 : _GEN_176 ? _slots_3_io_uop_lrs1 : _GEN_162 ? _slots_2_io_uop_lrs1 : _GEN_148 ? _slots_1_io_uop_lrs1 : _GEN_141 ? _slots_0_io_uop_lrs1 : 6'h0;
  assign io_iss_uops_0_lrs2 = _GEN_677 ? _slots_39_io_uop_lrs2 : _GEN_666 ? _slots_38_io_uop_lrs2 : _GEN_652 ? _slots_37_io_uop_lrs2 : _GEN_638 ? _slots_36_io_uop_lrs2 : _GEN_624 ? _slots_35_io_uop_lrs2 : _GEN_610 ? _slots_34_io_uop_lrs2 : _GEN_596 ? _slots_33_io_uop_lrs2 : _GEN_582 ? _slots_32_io_uop_lrs2 : _GEN_568 ? _slots_31_io_uop_lrs2 : _GEN_554 ? _slots_30_io_uop_lrs2 : _GEN_540 ? _slots_29_io_uop_lrs2 : _GEN_526 ? _slots_28_io_uop_lrs2 : _GEN_512 ? _slots_27_io_uop_lrs2 : _GEN_498 ? _slots_26_io_uop_lrs2 : _GEN_484 ? _slots_25_io_uop_lrs2 : _GEN_470 ? _slots_24_io_uop_lrs2 : _GEN_456 ? _slots_23_io_uop_lrs2 : _GEN_442 ? _slots_22_io_uop_lrs2 : _GEN_428 ? _slots_21_io_uop_lrs2 : _GEN_414 ? _slots_20_io_uop_lrs2 : _GEN_400 ? _slots_19_io_uop_lrs2 : _GEN_386 ? _slots_18_io_uop_lrs2 : _GEN_372 ? _slots_17_io_uop_lrs2 : _GEN_358 ? _slots_16_io_uop_lrs2 : _GEN_344 ? _slots_15_io_uop_lrs2 : _GEN_330 ? _slots_14_io_uop_lrs2 : _GEN_316 ? _slots_13_io_uop_lrs2 : _GEN_302 ? _slots_12_io_uop_lrs2 : _GEN_288 ? _slots_11_io_uop_lrs2 : _GEN_274 ? _slots_10_io_uop_lrs2 : _GEN_260 ? _slots_9_io_uop_lrs2 : _GEN_246 ? _slots_8_io_uop_lrs2 : _GEN_232 ? _slots_7_io_uop_lrs2 : _GEN_218 ? _slots_6_io_uop_lrs2 : _GEN_204 ? _slots_5_io_uop_lrs2 : _GEN_190 ? _slots_4_io_uop_lrs2 : _GEN_176 ? _slots_3_io_uop_lrs2 : _GEN_162 ? _slots_2_io_uop_lrs2 : _GEN_148 ? _slots_1_io_uop_lrs2 : _GEN_141 ? _slots_0_io_uop_lrs2 : 6'h0;
  assign io_iss_uops_0_lrs3 = _GEN_677 ? _slots_39_io_uop_lrs3 : _GEN_666 ? _slots_38_io_uop_lrs3 : _GEN_652 ? _slots_37_io_uop_lrs3 : _GEN_638 ? _slots_36_io_uop_lrs3 : _GEN_624 ? _slots_35_io_uop_lrs3 : _GEN_610 ? _slots_34_io_uop_lrs3 : _GEN_596 ? _slots_33_io_uop_lrs3 : _GEN_582 ? _slots_32_io_uop_lrs3 : _GEN_568 ? _slots_31_io_uop_lrs3 : _GEN_554 ? _slots_30_io_uop_lrs3 : _GEN_540 ? _slots_29_io_uop_lrs3 : _GEN_526 ? _slots_28_io_uop_lrs3 : _GEN_512 ? _slots_27_io_uop_lrs3 : _GEN_498 ? _slots_26_io_uop_lrs3 : _GEN_484 ? _slots_25_io_uop_lrs3 : _GEN_470 ? _slots_24_io_uop_lrs3 : _GEN_456 ? _slots_23_io_uop_lrs3 : _GEN_442 ? _slots_22_io_uop_lrs3 : _GEN_428 ? _slots_21_io_uop_lrs3 : _GEN_414 ? _slots_20_io_uop_lrs3 : _GEN_400 ? _slots_19_io_uop_lrs3 : _GEN_386 ? _slots_18_io_uop_lrs3 : _GEN_372 ? _slots_17_io_uop_lrs3 : _GEN_358 ? _slots_16_io_uop_lrs3 : _GEN_344 ? _slots_15_io_uop_lrs3 : _GEN_330 ? _slots_14_io_uop_lrs3 : _GEN_316 ? _slots_13_io_uop_lrs3 : _GEN_302 ? _slots_12_io_uop_lrs3 : _GEN_288 ? _slots_11_io_uop_lrs3 : _GEN_274 ? _slots_10_io_uop_lrs3 : _GEN_260 ? _slots_9_io_uop_lrs3 : _GEN_246 ? _slots_8_io_uop_lrs3 : _GEN_232 ? _slots_7_io_uop_lrs3 : _GEN_218 ? _slots_6_io_uop_lrs3 : _GEN_204 ? _slots_5_io_uop_lrs3 : _GEN_190 ? _slots_4_io_uop_lrs3 : _GEN_176 ? _slots_3_io_uop_lrs3 : _GEN_162 ? _slots_2_io_uop_lrs3 : _GEN_148 ? _slots_1_io_uop_lrs3 : _GEN_141 ? _slots_0_io_uop_lrs3 : 6'h0;
  assign io_iss_uops_0_ldst_val = _GEN_677 ? _slots_39_io_uop_ldst_val : _GEN_666 ? _slots_38_io_uop_ldst_val : _GEN_652 ? _slots_37_io_uop_ldst_val : _GEN_638 ? _slots_36_io_uop_ldst_val : _GEN_624 ? _slots_35_io_uop_ldst_val : _GEN_610 ? _slots_34_io_uop_ldst_val : _GEN_596 ? _slots_33_io_uop_ldst_val : _GEN_582 ? _slots_32_io_uop_ldst_val : _GEN_568 ? _slots_31_io_uop_ldst_val : _GEN_554 ? _slots_30_io_uop_ldst_val : _GEN_540 ? _slots_29_io_uop_ldst_val : _GEN_526 ? _slots_28_io_uop_ldst_val : _GEN_512 ? _slots_27_io_uop_ldst_val : _GEN_498 ? _slots_26_io_uop_ldst_val : _GEN_484 ? _slots_25_io_uop_ldst_val : _GEN_470 ? _slots_24_io_uop_ldst_val : _GEN_456 ? _slots_23_io_uop_ldst_val : _GEN_442 ? _slots_22_io_uop_ldst_val : _GEN_428 ? _slots_21_io_uop_ldst_val : _GEN_414 ? _slots_20_io_uop_ldst_val : _GEN_400 ? _slots_19_io_uop_ldst_val : _GEN_386 ? _slots_18_io_uop_ldst_val : _GEN_372 ? _slots_17_io_uop_ldst_val : _GEN_358 ? _slots_16_io_uop_ldst_val : _GEN_344 ? _slots_15_io_uop_ldst_val : _GEN_330 ? _slots_14_io_uop_ldst_val : _GEN_316 ? _slots_13_io_uop_ldst_val : _GEN_302 ? _slots_12_io_uop_ldst_val : _GEN_288 ? _slots_11_io_uop_ldst_val : _GEN_274 ? _slots_10_io_uop_ldst_val : _GEN_260 ? _slots_9_io_uop_ldst_val : _GEN_246 ? _slots_8_io_uop_ldst_val : _GEN_232 ? _slots_7_io_uop_ldst_val : _GEN_218 ? _slots_6_io_uop_ldst_val : _GEN_204 ? _slots_5_io_uop_ldst_val : _GEN_190 ? _slots_4_io_uop_ldst_val : _GEN_176 ? _slots_3_io_uop_ldst_val : _GEN_162 ? _slots_2_io_uop_ldst_val : _GEN_148 ? _slots_1_io_uop_ldst_val : _GEN_141 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_0_dst_rtype = _GEN_677 ? _slots_39_io_uop_dst_rtype : _GEN_666 ? _slots_38_io_uop_dst_rtype : _GEN_652 ? _slots_37_io_uop_dst_rtype : _GEN_638 ? _slots_36_io_uop_dst_rtype : _GEN_624 ? _slots_35_io_uop_dst_rtype : _GEN_610 ? _slots_34_io_uop_dst_rtype : _GEN_596 ? _slots_33_io_uop_dst_rtype : _GEN_582 ? _slots_32_io_uop_dst_rtype : _GEN_568 ? _slots_31_io_uop_dst_rtype : _GEN_554 ? _slots_30_io_uop_dst_rtype : _GEN_540 ? _slots_29_io_uop_dst_rtype : _GEN_526 ? _slots_28_io_uop_dst_rtype : _GEN_512 ? _slots_27_io_uop_dst_rtype : _GEN_498 ? _slots_26_io_uop_dst_rtype : _GEN_484 ? _slots_25_io_uop_dst_rtype : _GEN_470 ? _slots_24_io_uop_dst_rtype : _GEN_456 ? _slots_23_io_uop_dst_rtype : _GEN_442 ? _slots_22_io_uop_dst_rtype : _GEN_428 ? _slots_21_io_uop_dst_rtype : _GEN_414 ? _slots_20_io_uop_dst_rtype : _GEN_400 ? _slots_19_io_uop_dst_rtype : _GEN_386 ? _slots_18_io_uop_dst_rtype : _GEN_372 ? _slots_17_io_uop_dst_rtype : _GEN_358 ? _slots_16_io_uop_dst_rtype : _GEN_344 ? _slots_15_io_uop_dst_rtype : _GEN_330 ? _slots_14_io_uop_dst_rtype : _GEN_316 ? _slots_13_io_uop_dst_rtype : _GEN_302 ? _slots_12_io_uop_dst_rtype : _GEN_288 ? _slots_11_io_uop_dst_rtype : _GEN_274 ? _slots_10_io_uop_dst_rtype : _GEN_260 ? _slots_9_io_uop_dst_rtype : _GEN_246 ? _slots_8_io_uop_dst_rtype : _GEN_232 ? _slots_7_io_uop_dst_rtype : _GEN_218 ? _slots_6_io_uop_dst_rtype : _GEN_204 ? _slots_5_io_uop_dst_rtype : _GEN_190 ? _slots_4_io_uop_dst_rtype : _GEN_176 ? _slots_3_io_uop_dst_rtype : _GEN_162 ? _slots_2_io_uop_dst_rtype : _GEN_148 ? _slots_1_io_uop_dst_rtype : _GEN_141 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_0_lrs1_rtype = _GEN_677 ? _slots_39_io_uop_lrs1_rtype : _GEN_666 ? _slots_38_io_uop_lrs1_rtype : _GEN_652 ? _slots_37_io_uop_lrs1_rtype : _GEN_638 ? _slots_36_io_uop_lrs1_rtype : _GEN_624 ? _slots_35_io_uop_lrs1_rtype : _GEN_610 ? _slots_34_io_uop_lrs1_rtype : _GEN_596 ? _slots_33_io_uop_lrs1_rtype : _GEN_582 ? _slots_32_io_uop_lrs1_rtype : _GEN_568 ? _slots_31_io_uop_lrs1_rtype : _GEN_554 ? _slots_30_io_uop_lrs1_rtype : _GEN_540 ? _slots_29_io_uop_lrs1_rtype : _GEN_526 ? _slots_28_io_uop_lrs1_rtype : _GEN_512 ? _slots_27_io_uop_lrs1_rtype : _GEN_498 ? _slots_26_io_uop_lrs1_rtype : _GEN_484 ? _slots_25_io_uop_lrs1_rtype : _GEN_470 ? _slots_24_io_uop_lrs1_rtype : _GEN_456 ? _slots_23_io_uop_lrs1_rtype : _GEN_442 ? _slots_22_io_uop_lrs1_rtype : _GEN_428 ? _slots_21_io_uop_lrs1_rtype : _GEN_414 ? _slots_20_io_uop_lrs1_rtype : _GEN_400 ? _slots_19_io_uop_lrs1_rtype : _GEN_386 ? _slots_18_io_uop_lrs1_rtype : _GEN_372 ? _slots_17_io_uop_lrs1_rtype : _GEN_358 ? _slots_16_io_uop_lrs1_rtype : _GEN_344 ? _slots_15_io_uop_lrs1_rtype : _GEN_330 ? _slots_14_io_uop_lrs1_rtype : _GEN_316 ? _slots_13_io_uop_lrs1_rtype : _GEN_302 ? _slots_12_io_uop_lrs1_rtype : _GEN_288 ? _slots_11_io_uop_lrs1_rtype : _GEN_274 ? _slots_10_io_uop_lrs1_rtype : _GEN_260 ? _slots_9_io_uop_lrs1_rtype : _GEN_246 ? _slots_8_io_uop_lrs1_rtype : _GEN_232 ? _slots_7_io_uop_lrs1_rtype : _GEN_218 ? _slots_6_io_uop_lrs1_rtype : _GEN_204 ? _slots_5_io_uop_lrs1_rtype : _GEN_190 ? _slots_4_io_uop_lrs1_rtype : _GEN_176 ? _slots_3_io_uop_lrs1_rtype : _GEN_162 ? _slots_2_io_uop_lrs1_rtype : _GEN_148 ? _slots_1_io_uop_lrs1_rtype : _GEN_141 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_0_lrs2_rtype = _GEN_677 ? _slots_39_io_uop_lrs2_rtype : _GEN_666 ? _slots_38_io_uop_lrs2_rtype : _GEN_652 ? _slots_37_io_uop_lrs2_rtype : _GEN_638 ? _slots_36_io_uop_lrs2_rtype : _GEN_624 ? _slots_35_io_uop_lrs2_rtype : _GEN_610 ? _slots_34_io_uop_lrs2_rtype : _GEN_596 ? _slots_33_io_uop_lrs2_rtype : _GEN_582 ? _slots_32_io_uop_lrs2_rtype : _GEN_568 ? _slots_31_io_uop_lrs2_rtype : _GEN_554 ? _slots_30_io_uop_lrs2_rtype : _GEN_540 ? _slots_29_io_uop_lrs2_rtype : _GEN_526 ? _slots_28_io_uop_lrs2_rtype : _GEN_512 ? _slots_27_io_uop_lrs2_rtype : _GEN_498 ? _slots_26_io_uop_lrs2_rtype : _GEN_484 ? _slots_25_io_uop_lrs2_rtype : _GEN_470 ? _slots_24_io_uop_lrs2_rtype : _GEN_456 ? _slots_23_io_uop_lrs2_rtype : _GEN_442 ? _slots_22_io_uop_lrs2_rtype : _GEN_428 ? _slots_21_io_uop_lrs2_rtype : _GEN_414 ? _slots_20_io_uop_lrs2_rtype : _GEN_400 ? _slots_19_io_uop_lrs2_rtype : _GEN_386 ? _slots_18_io_uop_lrs2_rtype : _GEN_372 ? _slots_17_io_uop_lrs2_rtype : _GEN_358 ? _slots_16_io_uop_lrs2_rtype : _GEN_344 ? _slots_15_io_uop_lrs2_rtype : _GEN_330 ? _slots_14_io_uop_lrs2_rtype : _GEN_316 ? _slots_13_io_uop_lrs2_rtype : _GEN_302 ? _slots_12_io_uop_lrs2_rtype : _GEN_288 ? _slots_11_io_uop_lrs2_rtype : _GEN_274 ? _slots_10_io_uop_lrs2_rtype : _GEN_260 ? _slots_9_io_uop_lrs2_rtype : _GEN_246 ? _slots_8_io_uop_lrs2_rtype : _GEN_232 ? _slots_7_io_uop_lrs2_rtype : _GEN_218 ? _slots_6_io_uop_lrs2_rtype : _GEN_204 ? _slots_5_io_uop_lrs2_rtype : _GEN_190 ? _slots_4_io_uop_lrs2_rtype : _GEN_176 ? _slots_3_io_uop_lrs2_rtype : _GEN_162 ? _slots_2_io_uop_lrs2_rtype : _GEN_148 ? _slots_1_io_uop_lrs2_rtype : _GEN_141 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_0_frs3_en = _GEN_677 ? _slots_39_io_uop_frs3_en : _GEN_666 ? _slots_38_io_uop_frs3_en : _GEN_652 ? _slots_37_io_uop_frs3_en : _GEN_638 ? _slots_36_io_uop_frs3_en : _GEN_624 ? _slots_35_io_uop_frs3_en : _GEN_610 ? _slots_34_io_uop_frs3_en : _GEN_596 ? _slots_33_io_uop_frs3_en : _GEN_582 ? _slots_32_io_uop_frs3_en : _GEN_568 ? _slots_31_io_uop_frs3_en : _GEN_554 ? _slots_30_io_uop_frs3_en : _GEN_540 ? _slots_29_io_uop_frs3_en : _GEN_526 ? _slots_28_io_uop_frs3_en : _GEN_512 ? _slots_27_io_uop_frs3_en : _GEN_498 ? _slots_26_io_uop_frs3_en : _GEN_484 ? _slots_25_io_uop_frs3_en : _GEN_470 ? _slots_24_io_uop_frs3_en : _GEN_456 ? _slots_23_io_uop_frs3_en : _GEN_442 ? _slots_22_io_uop_frs3_en : _GEN_428 ? _slots_21_io_uop_frs3_en : _GEN_414 ? _slots_20_io_uop_frs3_en : _GEN_400 ? _slots_19_io_uop_frs3_en : _GEN_386 ? _slots_18_io_uop_frs3_en : _GEN_372 ? _slots_17_io_uop_frs3_en : _GEN_358 ? _slots_16_io_uop_frs3_en : _GEN_344 ? _slots_15_io_uop_frs3_en : _GEN_330 ? _slots_14_io_uop_frs3_en : _GEN_316 ? _slots_13_io_uop_frs3_en : _GEN_302 ? _slots_12_io_uop_frs3_en : _GEN_288 ? _slots_11_io_uop_frs3_en : _GEN_274 ? _slots_10_io_uop_frs3_en : _GEN_260 ? _slots_9_io_uop_frs3_en : _GEN_246 ? _slots_8_io_uop_frs3_en : _GEN_232 ? _slots_7_io_uop_frs3_en : _GEN_218 ? _slots_6_io_uop_frs3_en : _GEN_204 ? _slots_5_io_uop_frs3_en : _GEN_190 ? _slots_4_io_uop_frs3_en : _GEN_176 ? _slots_3_io_uop_frs3_en : _GEN_162 ? _slots_2_io_uop_frs3_en : _GEN_148 ? _slots_1_io_uop_frs3_en : _GEN_141 & _slots_0_io_uop_frs3_en;
  assign io_iss_uops_0_fp_val = _GEN_677 ? _slots_39_io_uop_fp_val : _GEN_666 ? _slots_38_io_uop_fp_val : _GEN_652 ? _slots_37_io_uop_fp_val : _GEN_638 ? _slots_36_io_uop_fp_val : _GEN_624 ? _slots_35_io_uop_fp_val : _GEN_610 ? _slots_34_io_uop_fp_val : _GEN_596 ? _slots_33_io_uop_fp_val : _GEN_582 ? _slots_32_io_uop_fp_val : _GEN_568 ? _slots_31_io_uop_fp_val : _GEN_554 ? _slots_30_io_uop_fp_val : _GEN_540 ? _slots_29_io_uop_fp_val : _GEN_526 ? _slots_28_io_uop_fp_val : _GEN_512 ? _slots_27_io_uop_fp_val : _GEN_498 ? _slots_26_io_uop_fp_val : _GEN_484 ? _slots_25_io_uop_fp_val : _GEN_470 ? _slots_24_io_uop_fp_val : _GEN_456 ? _slots_23_io_uop_fp_val : _GEN_442 ? _slots_22_io_uop_fp_val : _GEN_428 ? _slots_21_io_uop_fp_val : _GEN_414 ? _slots_20_io_uop_fp_val : _GEN_400 ? _slots_19_io_uop_fp_val : _GEN_386 ? _slots_18_io_uop_fp_val : _GEN_372 ? _slots_17_io_uop_fp_val : _GEN_358 ? _slots_16_io_uop_fp_val : _GEN_344 ? _slots_15_io_uop_fp_val : _GEN_330 ? _slots_14_io_uop_fp_val : _GEN_316 ? _slots_13_io_uop_fp_val : _GEN_302 ? _slots_12_io_uop_fp_val : _GEN_288 ? _slots_11_io_uop_fp_val : _GEN_274 ? _slots_10_io_uop_fp_val : _GEN_260 ? _slots_9_io_uop_fp_val : _GEN_246 ? _slots_8_io_uop_fp_val : _GEN_232 ? _slots_7_io_uop_fp_val : _GEN_218 ? _slots_6_io_uop_fp_val : _GEN_204 ? _slots_5_io_uop_fp_val : _GEN_190 ? _slots_4_io_uop_fp_val : _GEN_176 ? _slots_3_io_uop_fp_val : _GEN_162 ? _slots_2_io_uop_fp_val : _GEN_148 ? _slots_1_io_uop_fp_val : _GEN_141 & _slots_0_io_uop_fp_val;
  assign io_iss_uops_0_fp_single = _GEN_677 ? _slots_39_io_uop_fp_single : _GEN_666 ? _slots_38_io_uop_fp_single : _GEN_652 ? _slots_37_io_uop_fp_single : _GEN_638 ? _slots_36_io_uop_fp_single : _GEN_624 ? _slots_35_io_uop_fp_single : _GEN_610 ? _slots_34_io_uop_fp_single : _GEN_596 ? _slots_33_io_uop_fp_single : _GEN_582 ? _slots_32_io_uop_fp_single : _GEN_568 ? _slots_31_io_uop_fp_single : _GEN_554 ? _slots_30_io_uop_fp_single : _GEN_540 ? _slots_29_io_uop_fp_single : _GEN_526 ? _slots_28_io_uop_fp_single : _GEN_512 ? _slots_27_io_uop_fp_single : _GEN_498 ? _slots_26_io_uop_fp_single : _GEN_484 ? _slots_25_io_uop_fp_single : _GEN_470 ? _slots_24_io_uop_fp_single : _GEN_456 ? _slots_23_io_uop_fp_single : _GEN_442 ? _slots_22_io_uop_fp_single : _GEN_428 ? _slots_21_io_uop_fp_single : _GEN_414 ? _slots_20_io_uop_fp_single : _GEN_400 ? _slots_19_io_uop_fp_single : _GEN_386 ? _slots_18_io_uop_fp_single : _GEN_372 ? _slots_17_io_uop_fp_single : _GEN_358 ? _slots_16_io_uop_fp_single : _GEN_344 ? _slots_15_io_uop_fp_single : _GEN_330 ? _slots_14_io_uop_fp_single : _GEN_316 ? _slots_13_io_uop_fp_single : _GEN_302 ? _slots_12_io_uop_fp_single : _GEN_288 ? _slots_11_io_uop_fp_single : _GEN_274 ? _slots_10_io_uop_fp_single : _GEN_260 ? _slots_9_io_uop_fp_single : _GEN_246 ? _slots_8_io_uop_fp_single : _GEN_232 ? _slots_7_io_uop_fp_single : _GEN_218 ? _slots_6_io_uop_fp_single : _GEN_204 ? _slots_5_io_uop_fp_single : _GEN_190 ? _slots_4_io_uop_fp_single : _GEN_176 ? _slots_3_io_uop_fp_single : _GEN_162 ? _slots_2_io_uop_fp_single : _GEN_148 ? _slots_1_io_uop_fp_single : _GEN_141 & _slots_0_io_uop_fp_single;
  assign io_iss_uops_0_xcpt_pf_if = _GEN_677 ? _slots_39_io_uop_xcpt_pf_if : _GEN_666 ? _slots_38_io_uop_xcpt_pf_if : _GEN_652 ? _slots_37_io_uop_xcpt_pf_if : _GEN_638 ? _slots_36_io_uop_xcpt_pf_if : _GEN_624 ? _slots_35_io_uop_xcpt_pf_if : _GEN_610 ? _slots_34_io_uop_xcpt_pf_if : _GEN_596 ? _slots_33_io_uop_xcpt_pf_if : _GEN_582 ? _slots_32_io_uop_xcpt_pf_if : _GEN_568 ? _slots_31_io_uop_xcpt_pf_if : _GEN_554 ? _slots_30_io_uop_xcpt_pf_if : _GEN_540 ? _slots_29_io_uop_xcpt_pf_if : _GEN_526 ? _slots_28_io_uop_xcpt_pf_if : _GEN_512 ? _slots_27_io_uop_xcpt_pf_if : _GEN_498 ? _slots_26_io_uop_xcpt_pf_if : _GEN_484 ? _slots_25_io_uop_xcpt_pf_if : _GEN_470 ? _slots_24_io_uop_xcpt_pf_if : _GEN_456 ? _slots_23_io_uop_xcpt_pf_if : _GEN_442 ? _slots_22_io_uop_xcpt_pf_if : _GEN_428 ? _slots_21_io_uop_xcpt_pf_if : _GEN_414 ? _slots_20_io_uop_xcpt_pf_if : _GEN_400 ? _slots_19_io_uop_xcpt_pf_if : _GEN_386 ? _slots_18_io_uop_xcpt_pf_if : _GEN_372 ? _slots_17_io_uop_xcpt_pf_if : _GEN_358 ? _slots_16_io_uop_xcpt_pf_if : _GEN_344 ? _slots_15_io_uop_xcpt_pf_if : _GEN_330 ? _slots_14_io_uop_xcpt_pf_if : _GEN_316 ? _slots_13_io_uop_xcpt_pf_if : _GEN_302 ? _slots_12_io_uop_xcpt_pf_if : _GEN_288 ? _slots_11_io_uop_xcpt_pf_if : _GEN_274 ? _slots_10_io_uop_xcpt_pf_if : _GEN_260 ? _slots_9_io_uop_xcpt_pf_if : _GEN_246 ? _slots_8_io_uop_xcpt_pf_if : _GEN_232 ? _slots_7_io_uop_xcpt_pf_if : _GEN_218 ? _slots_6_io_uop_xcpt_pf_if : _GEN_204 ? _slots_5_io_uop_xcpt_pf_if : _GEN_190 ? _slots_4_io_uop_xcpt_pf_if : _GEN_176 ? _slots_3_io_uop_xcpt_pf_if : _GEN_162 ? _slots_2_io_uop_xcpt_pf_if : _GEN_148 ? _slots_1_io_uop_xcpt_pf_if : _GEN_141 & _slots_0_io_uop_xcpt_pf_if;
  assign io_iss_uops_0_xcpt_ae_if = _GEN_677 ? _slots_39_io_uop_xcpt_ae_if : _GEN_666 ? _slots_38_io_uop_xcpt_ae_if : _GEN_652 ? _slots_37_io_uop_xcpt_ae_if : _GEN_638 ? _slots_36_io_uop_xcpt_ae_if : _GEN_624 ? _slots_35_io_uop_xcpt_ae_if : _GEN_610 ? _slots_34_io_uop_xcpt_ae_if : _GEN_596 ? _slots_33_io_uop_xcpt_ae_if : _GEN_582 ? _slots_32_io_uop_xcpt_ae_if : _GEN_568 ? _slots_31_io_uop_xcpt_ae_if : _GEN_554 ? _slots_30_io_uop_xcpt_ae_if : _GEN_540 ? _slots_29_io_uop_xcpt_ae_if : _GEN_526 ? _slots_28_io_uop_xcpt_ae_if : _GEN_512 ? _slots_27_io_uop_xcpt_ae_if : _GEN_498 ? _slots_26_io_uop_xcpt_ae_if : _GEN_484 ? _slots_25_io_uop_xcpt_ae_if : _GEN_470 ? _slots_24_io_uop_xcpt_ae_if : _GEN_456 ? _slots_23_io_uop_xcpt_ae_if : _GEN_442 ? _slots_22_io_uop_xcpt_ae_if : _GEN_428 ? _slots_21_io_uop_xcpt_ae_if : _GEN_414 ? _slots_20_io_uop_xcpt_ae_if : _GEN_400 ? _slots_19_io_uop_xcpt_ae_if : _GEN_386 ? _slots_18_io_uop_xcpt_ae_if : _GEN_372 ? _slots_17_io_uop_xcpt_ae_if : _GEN_358 ? _slots_16_io_uop_xcpt_ae_if : _GEN_344 ? _slots_15_io_uop_xcpt_ae_if : _GEN_330 ? _slots_14_io_uop_xcpt_ae_if : _GEN_316 ? _slots_13_io_uop_xcpt_ae_if : _GEN_302 ? _slots_12_io_uop_xcpt_ae_if : _GEN_288 ? _slots_11_io_uop_xcpt_ae_if : _GEN_274 ? _slots_10_io_uop_xcpt_ae_if : _GEN_260 ? _slots_9_io_uop_xcpt_ae_if : _GEN_246 ? _slots_8_io_uop_xcpt_ae_if : _GEN_232 ? _slots_7_io_uop_xcpt_ae_if : _GEN_218 ? _slots_6_io_uop_xcpt_ae_if : _GEN_204 ? _slots_5_io_uop_xcpt_ae_if : _GEN_190 ? _slots_4_io_uop_xcpt_ae_if : _GEN_176 ? _slots_3_io_uop_xcpt_ae_if : _GEN_162 ? _slots_2_io_uop_xcpt_ae_if : _GEN_148 ? _slots_1_io_uop_xcpt_ae_if : _GEN_141 & _slots_0_io_uop_xcpt_ae_if;
  assign io_iss_uops_0_xcpt_ma_if = _GEN_677 ? _slots_39_io_uop_xcpt_ma_if : _GEN_666 ? _slots_38_io_uop_xcpt_ma_if : _GEN_652 ? _slots_37_io_uop_xcpt_ma_if : _GEN_638 ? _slots_36_io_uop_xcpt_ma_if : _GEN_624 ? _slots_35_io_uop_xcpt_ma_if : _GEN_610 ? _slots_34_io_uop_xcpt_ma_if : _GEN_596 ? _slots_33_io_uop_xcpt_ma_if : _GEN_582 ? _slots_32_io_uop_xcpt_ma_if : _GEN_568 ? _slots_31_io_uop_xcpt_ma_if : _GEN_554 ? _slots_30_io_uop_xcpt_ma_if : _GEN_540 ? _slots_29_io_uop_xcpt_ma_if : _GEN_526 ? _slots_28_io_uop_xcpt_ma_if : _GEN_512 ? _slots_27_io_uop_xcpt_ma_if : _GEN_498 ? _slots_26_io_uop_xcpt_ma_if : _GEN_484 ? _slots_25_io_uop_xcpt_ma_if : _GEN_470 ? _slots_24_io_uop_xcpt_ma_if : _GEN_456 ? _slots_23_io_uop_xcpt_ma_if : _GEN_442 ? _slots_22_io_uop_xcpt_ma_if : _GEN_428 ? _slots_21_io_uop_xcpt_ma_if : _GEN_414 ? _slots_20_io_uop_xcpt_ma_if : _GEN_400 ? _slots_19_io_uop_xcpt_ma_if : _GEN_386 ? _slots_18_io_uop_xcpt_ma_if : _GEN_372 ? _slots_17_io_uop_xcpt_ma_if : _GEN_358 ? _slots_16_io_uop_xcpt_ma_if : _GEN_344 ? _slots_15_io_uop_xcpt_ma_if : _GEN_330 ? _slots_14_io_uop_xcpt_ma_if : _GEN_316 ? _slots_13_io_uop_xcpt_ma_if : _GEN_302 ? _slots_12_io_uop_xcpt_ma_if : _GEN_288 ? _slots_11_io_uop_xcpt_ma_if : _GEN_274 ? _slots_10_io_uop_xcpt_ma_if : _GEN_260 ? _slots_9_io_uop_xcpt_ma_if : _GEN_246 ? _slots_8_io_uop_xcpt_ma_if : _GEN_232 ? _slots_7_io_uop_xcpt_ma_if : _GEN_218 ? _slots_6_io_uop_xcpt_ma_if : _GEN_204 ? _slots_5_io_uop_xcpt_ma_if : _GEN_190 ? _slots_4_io_uop_xcpt_ma_if : _GEN_176 ? _slots_3_io_uop_xcpt_ma_if : _GEN_162 ? _slots_2_io_uop_xcpt_ma_if : _GEN_148 ? _slots_1_io_uop_xcpt_ma_if : _GEN_141 & _slots_0_io_uop_xcpt_ma_if;
  assign io_iss_uops_0_bp_debug_if = _GEN_677 ? _slots_39_io_uop_bp_debug_if : _GEN_666 ? _slots_38_io_uop_bp_debug_if : _GEN_652 ? _slots_37_io_uop_bp_debug_if : _GEN_638 ? _slots_36_io_uop_bp_debug_if : _GEN_624 ? _slots_35_io_uop_bp_debug_if : _GEN_610 ? _slots_34_io_uop_bp_debug_if : _GEN_596 ? _slots_33_io_uop_bp_debug_if : _GEN_582 ? _slots_32_io_uop_bp_debug_if : _GEN_568 ? _slots_31_io_uop_bp_debug_if : _GEN_554 ? _slots_30_io_uop_bp_debug_if : _GEN_540 ? _slots_29_io_uop_bp_debug_if : _GEN_526 ? _slots_28_io_uop_bp_debug_if : _GEN_512 ? _slots_27_io_uop_bp_debug_if : _GEN_498 ? _slots_26_io_uop_bp_debug_if : _GEN_484 ? _slots_25_io_uop_bp_debug_if : _GEN_470 ? _slots_24_io_uop_bp_debug_if : _GEN_456 ? _slots_23_io_uop_bp_debug_if : _GEN_442 ? _slots_22_io_uop_bp_debug_if : _GEN_428 ? _slots_21_io_uop_bp_debug_if : _GEN_414 ? _slots_20_io_uop_bp_debug_if : _GEN_400 ? _slots_19_io_uop_bp_debug_if : _GEN_386 ? _slots_18_io_uop_bp_debug_if : _GEN_372 ? _slots_17_io_uop_bp_debug_if : _GEN_358 ? _slots_16_io_uop_bp_debug_if : _GEN_344 ? _slots_15_io_uop_bp_debug_if : _GEN_330 ? _slots_14_io_uop_bp_debug_if : _GEN_316 ? _slots_13_io_uop_bp_debug_if : _GEN_302 ? _slots_12_io_uop_bp_debug_if : _GEN_288 ? _slots_11_io_uop_bp_debug_if : _GEN_274 ? _slots_10_io_uop_bp_debug_if : _GEN_260 ? _slots_9_io_uop_bp_debug_if : _GEN_246 ? _slots_8_io_uop_bp_debug_if : _GEN_232 ? _slots_7_io_uop_bp_debug_if : _GEN_218 ? _slots_6_io_uop_bp_debug_if : _GEN_204 ? _slots_5_io_uop_bp_debug_if : _GEN_190 ? _slots_4_io_uop_bp_debug_if : _GEN_176 ? _slots_3_io_uop_bp_debug_if : _GEN_162 ? _slots_2_io_uop_bp_debug_if : _GEN_148 ? _slots_1_io_uop_bp_debug_if : _GEN_141 & _slots_0_io_uop_bp_debug_if;
  assign io_iss_uops_0_bp_xcpt_if = _GEN_677 ? _slots_39_io_uop_bp_xcpt_if : _GEN_666 ? _slots_38_io_uop_bp_xcpt_if : _GEN_652 ? _slots_37_io_uop_bp_xcpt_if : _GEN_638 ? _slots_36_io_uop_bp_xcpt_if : _GEN_624 ? _slots_35_io_uop_bp_xcpt_if : _GEN_610 ? _slots_34_io_uop_bp_xcpt_if : _GEN_596 ? _slots_33_io_uop_bp_xcpt_if : _GEN_582 ? _slots_32_io_uop_bp_xcpt_if : _GEN_568 ? _slots_31_io_uop_bp_xcpt_if : _GEN_554 ? _slots_30_io_uop_bp_xcpt_if : _GEN_540 ? _slots_29_io_uop_bp_xcpt_if : _GEN_526 ? _slots_28_io_uop_bp_xcpt_if : _GEN_512 ? _slots_27_io_uop_bp_xcpt_if : _GEN_498 ? _slots_26_io_uop_bp_xcpt_if : _GEN_484 ? _slots_25_io_uop_bp_xcpt_if : _GEN_470 ? _slots_24_io_uop_bp_xcpt_if : _GEN_456 ? _slots_23_io_uop_bp_xcpt_if : _GEN_442 ? _slots_22_io_uop_bp_xcpt_if : _GEN_428 ? _slots_21_io_uop_bp_xcpt_if : _GEN_414 ? _slots_20_io_uop_bp_xcpt_if : _GEN_400 ? _slots_19_io_uop_bp_xcpt_if : _GEN_386 ? _slots_18_io_uop_bp_xcpt_if : _GEN_372 ? _slots_17_io_uop_bp_xcpt_if : _GEN_358 ? _slots_16_io_uop_bp_xcpt_if : _GEN_344 ? _slots_15_io_uop_bp_xcpt_if : _GEN_330 ? _slots_14_io_uop_bp_xcpt_if : _GEN_316 ? _slots_13_io_uop_bp_xcpt_if : _GEN_302 ? _slots_12_io_uop_bp_xcpt_if : _GEN_288 ? _slots_11_io_uop_bp_xcpt_if : _GEN_274 ? _slots_10_io_uop_bp_xcpt_if : _GEN_260 ? _slots_9_io_uop_bp_xcpt_if : _GEN_246 ? _slots_8_io_uop_bp_xcpt_if : _GEN_232 ? _slots_7_io_uop_bp_xcpt_if : _GEN_218 ? _slots_6_io_uop_bp_xcpt_if : _GEN_204 ? _slots_5_io_uop_bp_xcpt_if : _GEN_190 ? _slots_4_io_uop_bp_xcpt_if : _GEN_176 ? _slots_3_io_uop_bp_xcpt_if : _GEN_162 ? _slots_2_io_uop_bp_xcpt_if : _GEN_148 ? _slots_1_io_uop_bp_xcpt_if : _GEN_141 & _slots_0_io_uop_bp_xcpt_if;
  assign io_iss_uops_0_debug_fsrc = _GEN_677 ? _slots_39_io_uop_debug_fsrc : _GEN_666 ? _slots_38_io_uop_debug_fsrc : _GEN_652 ? _slots_37_io_uop_debug_fsrc : _GEN_638 ? _slots_36_io_uop_debug_fsrc : _GEN_624 ? _slots_35_io_uop_debug_fsrc : _GEN_610 ? _slots_34_io_uop_debug_fsrc : _GEN_596 ? _slots_33_io_uop_debug_fsrc : _GEN_582 ? _slots_32_io_uop_debug_fsrc : _GEN_568 ? _slots_31_io_uop_debug_fsrc : _GEN_554 ? _slots_30_io_uop_debug_fsrc : _GEN_540 ? _slots_29_io_uop_debug_fsrc : _GEN_526 ? _slots_28_io_uop_debug_fsrc : _GEN_512 ? _slots_27_io_uop_debug_fsrc : _GEN_498 ? _slots_26_io_uop_debug_fsrc : _GEN_484 ? _slots_25_io_uop_debug_fsrc : _GEN_470 ? _slots_24_io_uop_debug_fsrc : _GEN_456 ? _slots_23_io_uop_debug_fsrc : _GEN_442 ? _slots_22_io_uop_debug_fsrc : _GEN_428 ? _slots_21_io_uop_debug_fsrc : _GEN_414 ? _slots_20_io_uop_debug_fsrc : _GEN_400 ? _slots_19_io_uop_debug_fsrc : _GEN_386 ? _slots_18_io_uop_debug_fsrc : _GEN_372 ? _slots_17_io_uop_debug_fsrc : _GEN_358 ? _slots_16_io_uop_debug_fsrc : _GEN_344 ? _slots_15_io_uop_debug_fsrc : _GEN_330 ? _slots_14_io_uop_debug_fsrc : _GEN_316 ? _slots_13_io_uop_debug_fsrc : _GEN_302 ? _slots_12_io_uop_debug_fsrc : _GEN_288 ? _slots_11_io_uop_debug_fsrc : _GEN_274 ? _slots_10_io_uop_debug_fsrc : _GEN_260 ? _slots_9_io_uop_debug_fsrc : _GEN_246 ? _slots_8_io_uop_debug_fsrc : _GEN_232 ? _slots_7_io_uop_debug_fsrc : _GEN_218 ? _slots_6_io_uop_debug_fsrc : _GEN_204 ? _slots_5_io_uop_debug_fsrc : _GEN_190 ? _slots_4_io_uop_debug_fsrc : _GEN_176 ? _slots_3_io_uop_debug_fsrc : _GEN_162 ? _slots_2_io_uop_debug_fsrc : _GEN_148 ? _slots_1_io_uop_debug_fsrc : _GEN_141 ? _slots_0_io_uop_debug_fsrc : 2'h0;
  assign io_iss_uops_0_debug_tsrc = _GEN_677 ? _slots_39_io_uop_debug_tsrc : _GEN_666 ? _slots_38_io_uop_debug_tsrc : _GEN_652 ? _slots_37_io_uop_debug_tsrc : _GEN_638 ? _slots_36_io_uop_debug_tsrc : _GEN_624 ? _slots_35_io_uop_debug_tsrc : _GEN_610 ? _slots_34_io_uop_debug_tsrc : _GEN_596 ? _slots_33_io_uop_debug_tsrc : _GEN_582 ? _slots_32_io_uop_debug_tsrc : _GEN_568 ? _slots_31_io_uop_debug_tsrc : _GEN_554 ? _slots_30_io_uop_debug_tsrc : _GEN_540 ? _slots_29_io_uop_debug_tsrc : _GEN_526 ? _slots_28_io_uop_debug_tsrc : _GEN_512 ? _slots_27_io_uop_debug_tsrc : _GEN_498 ? _slots_26_io_uop_debug_tsrc : _GEN_484 ? _slots_25_io_uop_debug_tsrc : _GEN_470 ? _slots_24_io_uop_debug_tsrc : _GEN_456 ? _slots_23_io_uop_debug_tsrc : _GEN_442 ? _slots_22_io_uop_debug_tsrc : _GEN_428 ? _slots_21_io_uop_debug_tsrc : _GEN_414 ? _slots_20_io_uop_debug_tsrc : _GEN_400 ? _slots_19_io_uop_debug_tsrc : _GEN_386 ? _slots_18_io_uop_debug_tsrc : _GEN_372 ? _slots_17_io_uop_debug_tsrc : _GEN_358 ? _slots_16_io_uop_debug_tsrc : _GEN_344 ? _slots_15_io_uop_debug_tsrc : _GEN_330 ? _slots_14_io_uop_debug_tsrc : _GEN_316 ? _slots_13_io_uop_debug_tsrc : _GEN_302 ? _slots_12_io_uop_debug_tsrc : _GEN_288 ? _slots_11_io_uop_debug_tsrc : _GEN_274 ? _slots_10_io_uop_debug_tsrc : _GEN_260 ? _slots_9_io_uop_debug_tsrc : _GEN_246 ? _slots_8_io_uop_debug_tsrc : _GEN_232 ? _slots_7_io_uop_debug_tsrc : _GEN_218 ? _slots_6_io_uop_debug_tsrc : _GEN_204 ? _slots_5_io_uop_debug_tsrc : _GEN_190 ? _slots_4_io_uop_debug_tsrc : _GEN_176 ? _slots_3_io_uop_debug_tsrc : _GEN_162 ? _slots_2_io_uop_debug_tsrc : _GEN_148 ? _slots_1_io_uop_debug_tsrc : _GEN_141 ? _slots_0_io_uop_debug_tsrc : 2'h0;
  assign io_iss_uops_1_uopc = _GEN_679 ? _slots_39_io_uop_uopc : _GEN_669 ? _slots_38_io_uop_uopc : _GEN_656 ? _slots_37_io_uop_uopc : _GEN_642 ? _slots_36_io_uop_uopc : _GEN_628 ? _slots_35_io_uop_uopc : _GEN_614 ? _slots_34_io_uop_uopc : _GEN_600 ? _slots_33_io_uop_uopc : _GEN_586 ? _slots_32_io_uop_uopc : _GEN_572 ? _slots_31_io_uop_uopc : _GEN_558 ? _slots_30_io_uop_uopc : _GEN_544 ? _slots_29_io_uop_uopc : _GEN_530 ? _slots_28_io_uop_uopc : _GEN_516 ? _slots_27_io_uop_uopc : _GEN_502 ? _slots_26_io_uop_uopc : _GEN_488 ? _slots_25_io_uop_uopc : _GEN_474 ? _slots_24_io_uop_uopc : _GEN_460 ? _slots_23_io_uop_uopc : _GEN_446 ? _slots_22_io_uop_uopc : _GEN_432 ? _slots_21_io_uop_uopc : _GEN_418 ? _slots_20_io_uop_uopc : _GEN_404 ? _slots_19_io_uop_uopc : _GEN_390 ? _slots_18_io_uop_uopc : _GEN_376 ? _slots_17_io_uop_uopc : _GEN_362 ? _slots_16_io_uop_uopc : _GEN_348 ? _slots_15_io_uop_uopc : _GEN_334 ? _slots_14_io_uop_uopc : _GEN_320 ? _slots_13_io_uop_uopc : _GEN_306 ? _slots_12_io_uop_uopc : _GEN_292 ? _slots_11_io_uop_uopc : _GEN_278 ? _slots_10_io_uop_uopc : _GEN_264 ? _slots_9_io_uop_uopc : _GEN_250 ? _slots_8_io_uop_uopc : _GEN_236 ? _slots_7_io_uop_uopc : _GEN_222 ? _slots_6_io_uop_uopc : _GEN_208 ? _slots_5_io_uop_uopc : _GEN_194 ? _slots_4_io_uop_uopc : _GEN_180 ? _slots_3_io_uop_uopc : _GEN_166 ? _slots_2_io_uop_uopc : _GEN_152 ? _slots_1_io_uop_uopc : _GEN_143 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_1_is_rvc = _GEN_679 ? _slots_39_io_uop_is_rvc : _GEN_669 ? _slots_38_io_uop_is_rvc : _GEN_656 ? _slots_37_io_uop_is_rvc : _GEN_642 ? _slots_36_io_uop_is_rvc : _GEN_628 ? _slots_35_io_uop_is_rvc : _GEN_614 ? _slots_34_io_uop_is_rvc : _GEN_600 ? _slots_33_io_uop_is_rvc : _GEN_586 ? _slots_32_io_uop_is_rvc : _GEN_572 ? _slots_31_io_uop_is_rvc : _GEN_558 ? _slots_30_io_uop_is_rvc : _GEN_544 ? _slots_29_io_uop_is_rvc : _GEN_530 ? _slots_28_io_uop_is_rvc : _GEN_516 ? _slots_27_io_uop_is_rvc : _GEN_502 ? _slots_26_io_uop_is_rvc : _GEN_488 ? _slots_25_io_uop_is_rvc : _GEN_474 ? _slots_24_io_uop_is_rvc : _GEN_460 ? _slots_23_io_uop_is_rvc : _GEN_446 ? _slots_22_io_uop_is_rvc : _GEN_432 ? _slots_21_io_uop_is_rvc : _GEN_418 ? _slots_20_io_uop_is_rvc : _GEN_404 ? _slots_19_io_uop_is_rvc : _GEN_390 ? _slots_18_io_uop_is_rvc : _GEN_376 ? _slots_17_io_uop_is_rvc : _GEN_362 ? _slots_16_io_uop_is_rvc : _GEN_348 ? _slots_15_io_uop_is_rvc : _GEN_334 ? _slots_14_io_uop_is_rvc : _GEN_320 ? _slots_13_io_uop_is_rvc : _GEN_306 ? _slots_12_io_uop_is_rvc : _GEN_292 ? _slots_11_io_uop_is_rvc : _GEN_278 ? _slots_10_io_uop_is_rvc : _GEN_264 ? _slots_9_io_uop_is_rvc : _GEN_250 ? _slots_8_io_uop_is_rvc : _GEN_236 ? _slots_7_io_uop_is_rvc : _GEN_222 ? _slots_6_io_uop_is_rvc : _GEN_208 ? _slots_5_io_uop_is_rvc : _GEN_194 ? _slots_4_io_uop_is_rvc : _GEN_180 ? _slots_3_io_uop_is_rvc : _GEN_166 ? _slots_2_io_uop_is_rvc : _GEN_152 ? _slots_1_io_uop_is_rvc : _GEN_143 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_1_fu_code = _GEN_679 ? _slots_39_io_uop_fu_code : _GEN_669 ? _slots_38_io_uop_fu_code : _GEN_656 ? _slots_37_io_uop_fu_code : _GEN_642 ? _slots_36_io_uop_fu_code : _GEN_628 ? _slots_35_io_uop_fu_code : _GEN_614 ? _slots_34_io_uop_fu_code : _GEN_600 ? _slots_33_io_uop_fu_code : _GEN_586 ? _slots_32_io_uop_fu_code : _GEN_572 ? _slots_31_io_uop_fu_code : _GEN_558 ? _slots_30_io_uop_fu_code : _GEN_544 ? _slots_29_io_uop_fu_code : _GEN_530 ? _slots_28_io_uop_fu_code : _GEN_516 ? _slots_27_io_uop_fu_code : _GEN_502 ? _slots_26_io_uop_fu_code : _GEN_488 ? _slots_25_io_uop_fu_code : _GEN_474 ? _slots_24_io_uop_fu_code : _GEN_460 ? _slots_23_io_uop_fu_code : _GEN_446 ? _slots_22_io_uop_fu_code : _GEN_432 ? _slots_21_io_uop_fu_code : _GEN_418 ? _slots_20_io_uop_fu_code : _GEN_404 ? _slots_19_io_uop_fu_code : _GEN_390 ? _slots_18_io_uop_fu_code : _GEN_376 ? _slots_17_io_uop_fu_code : _GEN_362 ? _slots_16_io_uop_fu_code : _GEN_348 ? _slots_15_io_uop_fu_code : _GEN_334 ? _slots_14_io_uop_fu_code : _GEN_320 ? _slots_13_io_uop_fu_code : _GEN_306 ? _slots_12_io_uop_fu_code : _GEN_292 ? _slots_11_io_uop_fu_code : _GEN_278 ? _slots_10_io_uop_fu_code : _GEN_264 ? _slots_9_io_uop_fu_code : _GEN_250 ? _slots_8_io_uop_fu_code : _GEN_236 ? _slots_7_io_uop_fu_code : _GEN_222 ? _slots_6_io_uop_fu_code : _GEN_208 ? _slots_5_io_uop_fu_code : _GEN_194 ? _slots_4_io_uop_fu_code : _GEN_180 ? _slots_3_io_uop_fu_code : _GEN_166 ? _slots_2_io_uop_fu_code : _GEN_152 ? _slots_1_io_uop_fu_code : _GEN_143 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_1_iw_p1_poisoned = _GEN_679 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_669 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_656 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_642 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_628 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_614 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_600 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_586 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_572 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_558 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_544 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_530 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_516 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_502 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_488 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_474 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_460 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_446 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_432 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_418 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_404 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_390 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_376 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_362 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_348 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_334 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_320 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_306 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_292 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_278 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_264 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_250 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_236 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_222 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_208 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_194 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_180 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_166 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_152 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_143 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_1_iw_p2_poisoned = _GEN_679 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_669 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_656 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_642 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_628 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_614 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_600 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_586 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_572 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_558 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_544 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_530 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_516 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_502 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_488 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_474 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_460 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_446 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_432 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_418 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_404 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_390 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_376 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_362 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_348 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_334 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_320 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_306 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_292 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_278 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_264 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_250 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_236 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_222 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_208 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_194 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_180 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_166 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_152 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_143 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_1_is_br = _GEN_679 ? _slots_39_io_uop_is_br : _GEN_669 ? _slots_38_io_uop_is_br : _GEN_656 ? _slots_37_io_uop_is_br : _GEN_642 ? _slots_36_io_uop_is_br : _GEN_628 ? _slots_35_io_uop_is_br : _GEN_614 ? _slots_34_io_uop_is_br : _GEN_600 ? _slots_33_io_uop_is_br : _GEN_586 ? _slots_32_io_uop_is_br : _GEN_572 ? _slots_31_io_uop_is_br : _GEN_558 ? _slots_30_io_uop_is_br : _GEN_544 ? _slots_29_io_uop_is_br : _GEN_530 ? _slots_28_io_uop_is_br : _GEN_516 ? _slots_27_io_uop_is_br : _GEN_502 ? _slots_26_io_uop_is_br : _GEN_488 ? _slots_25_io_uop_is_br : _GEN_474 ? _slots_24_io_uop_is_br : _GEN_460 ? _slots_23_io_uop_is_br : _GEN_446 ? _slots_22_io_uop_is_br : _GEN_432 ? _slots_21_io_uop_is_br : _GEN_418 ? _slots_20_io_uop_is_br : _GEN_404 ? _slots_19_io_uop_is_br : _GEN_390 ? _slots_18_io_uop_is_br : _GEN_376 ? _slots_17_io_uop_is_br : _GEN_362 ? _slots_16_io_uop_is_br : _GEN_348 ? _slots_15_io_uop_is_br : _GEN_334 ? _slots_14_io_uop_is_br : _GEN_320 ? _slots_13_io_uop_is_br : _GEN_306 ? _slots_12_io_uop_is_br : _GEN_292 ? _slots_11_io_uop_is_br : _GEN_278 ? _slots_10_io_uop_is_br : _GEN_264 ? _slots_9_io_uop_is_br : _GEN_250 ? _slots_8_io_uop_is_br : _GEN_236 ? _slots_7_io_uop_is_br : _GEN_222 ? _slots_6_io_uop_is_br : _GEN_208 ? _slots_5_io_uop_is_br : _GEN_194 ? _slots_4_io_uop_is_br : _GEN_180 ? _slots_3_io_uop_is_br : _GEN_166 ? _slots_2_io_uop_is_br : _GEN_152 ? _slots_1_io_uop_is_br : _GEN_143 & _slots_0_io_uop_is_br;
  assign io_iss_uops_1_is_jalr = _GEN_679 ? _slots_39_io_uop_is_jalr : _GEN_669 ? _slots_38_io_uop_is_jalr : _GEN_656 ? _slots_37_io_uop_is_jalr : _GEN_642 ? _slots_36_io_uop_is_jalr : _GEN_628 ? _slots_35_io_uop_is_jalr : _GEN_614 ? _slots_34_io_uop_is_jalr : _GEN_600 ? _slots_33_io_uop_is_jalr : _GEN_586 ? _slots_32_io_uop_is_jalr : _GEN_572 ? _slots_31_io_uop_is_jalr : _GEN_558 ? _slots_30_io_uop_is_jalr : _GEN_544 ? _slots_29_io_uop_is_jalr : _GEN_530 ? _slots_28_io_uop_is_jalr : _GEN_516 ? _slots_27_io_uop_is_jalr : _GEN_502 ? _slots_26_io_uop_is_jalr : _GEN_488 ? _slots_25_io_uop_is_jalr : _GEN_474 ? _slots_24_io_uop_is_jalr : _GEN_460 ? _slots_23_io_uop_is_jalr : _GEN_446 ? _slots_22_io_uop_is_jalr : _GEN_432 ? _slots_21_io_uop_is_jalr : _GEN_418 ? _slots_20_io_uop_is_jalr : _GEN_404 ? _slots_19_io_uop_is_jalr : _GEN_390 ? _slots_18_io_uop_is_jalr : _GEN_376 ? _slots_17_io_uop_is_jalr : _GEN_362 ? _slots_16_io_uop_is_jalr : _GEN_348 ? _slots_15_io_uop_is_jalr : _GEN_334 ? _slots_14_io_uop_is_jalr : _GEN_320 ? _slots_13_io_uop_is_jalr : _GEN_306 ? _slots_12_io_uop_is_jalr : _GEN_292 ? _slots_11_io_uop_is_jalr : _GEN_278 ? _slots_10_io_uop_is_jalr : _GEN_264 ? _slots_9_io_uop_is_jalr : _GEN_250 ? _slots_8_io_uop_is_jalr : _GEN_236 ? _slots_7_io_uop_is_jalr : _GEN_222 ? _slots_6_io_uop_is_jalr : _GEN_208 ? _slots_5_io_uop_is_jalr : _GEN_194 ? _slots_4_io_uop_is_jalr : _GEN_180 ? _slots_3_io_uop_is_jalr : _GEN_166 ? _slots_2_io_uop_is_jalr : _GEN_152 ? _slots_1_io_uop_is_jalr : _GEN_143 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_1_is_jal = _GEN_679 ? _slots_39_io_uop_is_jal : _GEN_669 ? _slots_38_io_uop_is_jal : _GEN_656 ? _slots_37_io_uop_is_jal : _GEN_642 ? _slots_36_io_uop_is_jal : _GEN_628 ? _slots_35_io_uop_is_jal : _GEN_614 ? _slots_34_io_uop_is_jal : _GEN_600 ? _slots_33_io_uop_is_jal : _GEN_586 ? _slots_32_io_uop_is_jal : _GEN_572 ? _slots_31_io_uop_is_jal : _GEN_558 ? _slots_30_io_uop_is_jal : _GEN_544 ? _slots_29_io_uop_is_jal : _GEN_530 ? _slots_28_io_uop_is_jal : _GEN_516 ? _slots_27_io_uop_is_jal : _GEN_502 ? _slots_26_io_uop_is_jal : _GEN_488 ? _slots_25_io_uop_is_jal : _GEN_474 ? _slots_24_io_uop_is_jal : _GEN_460 ? _slots_23_io_uop_is_jal : _GEN_446 ? _slots_22_io_uop_is_jal : _GEN_432 ? _slots_21_io_uop_is_jal : _GEN_418 ? _slots_20_io_uop_is_jal : _GEN_404 ? _slots_19_io_uop_is_jal : _GEN_390 ? _slots_18_io_uop_is_jal : _GEN_376 ? _slots_17_io_uop_is_jal : _GEN_362 ? _slots_16_io_uop_is_jal : _GEN_348 ? _slots_15_io_uop_is_jal : _GEN_334 ? _slots_14_io_uop_is_jal : _GEN_320 ? _slots_13_io_uop_is_jal : _GEN_306 ? _slots_12_io_uop_is_jal : _GEN_292 ? _slots_11_io_uop_is_jal : _GEN_278 ? _slots_10_io_uop_is_jal : _GEN_264 ? _slots_9_io_uop_is_jal : _GEN_250 ? _slots_8_io_uop_is_jal : _GEN_236 ? _slots_7_io_uop_is_jal : _GEN_222 ? _slots_6_io_uop_is_jal : _GEN_208 ? _slots_5_io_uop_is_jal : _GEN_194 ? _slots_4_io_uop_is_jal : _GEN_180 ? _slots_3_io_uop_is_jal : _GEN_166 ? _slots_2_io_uop_is_jal : _GEN_152 ? _slots_1_io_uop_is_jal : _GEN_143 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_1_is_sfb = _GEN_679 ? _slots_39_io_uop_is_sfb : _GEN_669 ? _slots_38_io_uop_is_sfb : _GEN_656 ? _slots_37_io_uop_is_sfb : _GEN_642 ? _slots_36_io_uop_is_sfb : _GEN_628 ? _slots_35_io_uop_is_sfb : _GEN_614 ? _slots_34_io_uop_is_sfb : _GEN_600 ? _slots_33_io_uop_is_sfb : _GEN_586 ? _slots_32_io_uop_is_sfb : _GEN_572 ? _slots_31_io_uop_is_sfb : _GEN_558 ? _slots_30_io_uop_is_sfb : _GEN_544 ? _slots_29_io_uop_is_sfb : _GEN_530 ? _slots_28_io_uop_is_sfb : _GEN_516 ? _slots_27_io_uop_is_sfb : _GEN_502 ? _slots_26_io_uop_is_sfb : _GEN_488 ? _slots_25_io_uop_is_sfb : _GEN_474 ? _slots_24_io_uop_is_sfb : _GEN_460 ? _slots_23_io_uop_is_sfb : _GEN_446 ? _slots_22_io_uop_is_sfb : _GEN_432 ? _slots_21_io_uop_is_sfb : _GEN_418 ? _slots_20_io_uop_is_sfb : _GEN_404 ? _slots_19_io_uop_is_sfb : _GEN_390 ? _slots_18_io_uop_is_sfb : _GEN_376 ? _slots_17_io_uop_is_sfb : _GEN_362 ? _slots_16_io_uop_is_sfb : _GEN_348 ? _slots_15_io_uop_is_sfb : _GEN_334 ? _slots_14_io_uop_is_sfb : _GEN_320 ? _slots_13_io_uop_is_sfb : _GEN_306 ? _slots_12_io_uop_is_sfb : _GEN_292 ? _slots_11_io_uop_is_sfb : _GEN_278 ? _slots_10_io_uop_is_sfb : _GEN_264 ? _slots_9_io_uop_is_sfb : _GEN_250 ? _slots_8_io_uop_is_sfb : _GEN_236 ? _slots_7_io_uop_is_sfb : _GEN_222 ? _slots_6_io_uop_is_sfb : _GEN_208 ? _slots_5_io_uop_is_sfb : _GEN_194 ? _slots_4_io_uop_is_sfb : _GEN_180 ? _slots_3_io_uop_is_sfb : _GEN_166 ? _slots_2_io_uop_is_sfb : _GEN_152 ? _slots_1_io_uop_is_sfb : _GEN_143 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_1_br_mask = _GEN_679 ? _slots_39_io_uop_br_mask : _GEN_669 ? _slots_38_io_uop_br_mask : _GEN_656 ? _slots_37_io_uop_br_mask : _GEN_642 ? _slots_36_io_uop_br_mask : _GEN_628 ? _slots_35_io_uop_br_mask : _GEN_614 ? _slots_34_io_uop_br_mask : _GEN_600 ? _slots_33_io_uop_br_mask : _GEN_586 ? _slots_32_io_uop_br_mask : _GEN_572 ? _slots_31_io_uop_br_mask : _GEN_558 ? _slots_30_io_uop_br_mask : _GEN_544 ? _slots_29_io_uop_br_mask : _GEN_530 ? _slots_28_io_uop_br_mask : _GEN_516 ? _slots_27_io_uop_br_mask : _GEN_502 ? _slots_26_io_uop_br_mask : _GEN_488 ? _slots_25_io_uop_br_mask : _GEN_474 ? _slots_24_io_uop_br_mask : _GEN_460 ? _slots_23_io_uop_br_mask : _GEN_446 ? _slots_22_io_uop_br_mask : _GEN_432 ? _slots_21_io_uop_br_mask : _GEN_418 ? _slots_20_io_uop_br_mask : _GEN_404 ? _slots_19_io_uop_br_mask : _GEN_390 ? _slots_18_io_uop_br_mask : _GEN_376 ? _slots_17_io_uop_br_mask : _GEN_362 ? _slots_16_io_uop_br_mask : _GEN_348 ? _slots_15_io_uop_br_mask : _GEN_334 ? _slots_14_io_uop_br_mask : _GEN_320 ? _slots_13_io_uop_br_mask : _GEN_306 ? _slots_12_io_uop_br_mask : _GEN_292 ? _slots_11_io_uop_br_mask : _GEN_278 ? _slots_10_io_uop_br_mask : _GEN_264 ? _slots_9_io_uop_br_mask : _GEN_250 ? _slots_8_io_uop_br_mask : _GEN_236 ? _slots_7_io_uop_br_mask : _GEN_222 ? _slots_6_io_uop_br_mask : _GEN_208 ? _slots_5_io_uop_br_mask : _GEN_194 ? _slots_4_io_uop_br_mask : _GEN_180 ? _slots_3_io_uop_br_mask : _GEN_166 ? _slots_2_io_uop_br_mask : _GEN_152 ? _slots_1_io_uop_br_mask : _GEN_143 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_1_br_tag = _GEN_679 ? _slots_39_io_uop_br_tag : _GEN_669 ? _slots_38_io_uop_br_tag : _GEN_656 ? _slots_37_io_uop_br_tag : _GEN_642 ? _slots_36_io_uop_br_tag : _GEN_628 ? _slots_35_io_uop_br_tag : _GEN_614 ? _slots_34_io_uop_br_tag : _GEN_600 ? _slots_33_io_uop_br_tag : _GEN_586 ? _slots_32_io_uop_br_tag : _GEN_572 ? _slots_31_io_uop_br_tag : _GEN_558 ? _slots_30_io_uop_br_tag : _GEN_544 ? _slots_29_io_uop_br_tag : _GEN_530 ? _slots_28_io_uop_br_tag : _GEN_516 ? _slots_27_io_uop_br_tag : _GEN_502 ? _slots_26_io_uop_br_tag : _GEN_488 ? _slots_25_io_uop_br_tag : _GEN_474 ? _slots_24_io_uop_br_tag : _GEN_460 ? _slots_23_io_uop_br_tag : _GEN_446 ? _slots_22_io_uop_br_tag : _GEN_432 ? _slots_21_io_uop_br_tag : _GEN_418 ? _slots_20_io_uop_br_tag : _GEN_404 ? _slots_19_io_uop_br_tag : _GEN_390 ? _slots_18_io_uop_br_tag : _GEN_376 ? _slots_17_io_uop_br_tag : _GEN_362 ? _slots_16_io_uop_br_tag : _GEN_348 ? _slots_15_io_uop_br_tag : _GEN_334 ? _slots_14_io_uop_br_tag : _GEN_320 ? _slots_13_io_uop_br_tag : _GEN_306 ? _slots_12_io_uop_br_tag : _GEN_292 ? _slots_11_io_uop_br_tag : _GEN_278 ? _slots_10_io_uop_br_tag : _GEN_264 ? _slots_9_io_uop_br_tag : _GEN_250 ? _slots_8_io_uop_br_tag : _GEN_236 ? _slots_7_io_uop_br_tag : _GEN_222 ? _slots_6_io_uop_br_tag : _GEN_208 ? _slots_5_io_uop_br_tag : _GEN_194 ? _slots_4_io_uop_br_tag : _GEN_180 ? _slots_3_io_uop_br_tag : _GEN_166 ? _slots_2_io_uop_br_tag : _GEN_152 ? _slots_1_io_uop_br_tag : _GEN_143 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_1_ftq_idx = _GEN_679 ? _slots_39_io_uop_ftq_idx : _GEN_669 ? _slots_38_io_uop_ftq_idx : _GEN_656 ? _slots_37_io_uop_ftq_idx : _GEN_642 ? _slots_36_io_uop_ftq_idx : _GEN_628 ? _slots_35_io_uop_ftq_idx : _GEN_614 ? _slots_34_io_uop_ftq_idx : _GEN_600 ? _slots_33_io_uop_ftq_idx : _GEN_586 ? _slots_32_io_uop_ftq_idx : _GEN_572 ? _slots_31_io_uop_ftq_idx : _GEN_558 ? _slots_30_io_uop_ftq_idx : _GEN_544 ? _slots_29_io_uop_ftq_idx : _GEN_530 ? _slots_28_io_uop_ftq_idx : _GEN_516 ? _slots_27_io_uop_ftq_idx : _GEN_502 ? _slots_26_io_uop_ftq_idx : _GEN_488 ? _slots_25_io_uop_ftq_idx : _GEN_474 ? _slots_24_io_uop_ftq_idx : _GEN_460 ? _slots_23_io_uop_ftq_idx : _GEN_446 ? _slots_22_io_uop_ftq_idx : _GEN_432 ? _slots_21_io_uop_ftq_idx : _GEN_418 ? _slots_20_io_uop_ftq_idx : _GEN_404 ? _slots_19_io_uop_ftq_idx : _GEN_390 ? _slots_18_io_uop_ftq_idx : _GEN_376 ? _slots_17_io_uop_ftq_idx : _GEN_362 ? _slots_16_io_uop_ftq_idx : _GEN_348 ? _slots_15_io_uop_ftq_idx : _GEN_334 ? _slots_14_io_uop_ftq_idx : _GEN_320 ? _slots_13_io_uop_ftq_idx : _GEN_306 ? _slots_12_io_uop_ftq_idx : _GEN_292 ? _slots_11_io_uop_ftq_idx : _GEN_278 ? _slots_10_io_uop_ftq_idx : _GEN_264 ? _slots_9_io_uop_ftq_idx : _GEN_250 ? _slots_8_io_uop_ftq_idx : _GEN_236 ? _slots_7_io_uop_ftq_idx : _GEN_222 ? _slots_6_io_uop_ftq_idx : _GEN_208 ? _slots_5_io_uop_ftq_idx : _GEN_194 ? _slots_4_io_uop_ftq_idx : _GEN_180 ? _slots_3_io_uop_ftq_idx : _GEN_166 ? _slots_2_io_uop_ftq_idx : _GEN_152 ? _slots_1_io_uop_ftq_idx : _GEN_143 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_1_edge_inst = _GEN_679 ? _slots_39_io_uop_edge_inst : _GEN_669 ? _slots_38_io_uop_edge_inst : _GEN_656 ? _slots_37_io_uop_edge_inst : _GEN_642 ? _slots_36_io_uop_edge_inst : _GEN_628 ? _slots_35_io_uop_edge_inst : _GEN_614 ? _slots_34_io_uop_edge_inst : _GEN_600 ? _slots_33_io_uop_edge_inst : _GEN_586 ? _slots_32_io_uop_edge_inst : _GEN_572 ? _slots_31_io_uop_edge_inst : _GEN_558 ? _slots_30_io_uop_edge_inst : _GEN_544 ? _slots_29_io_uop_edge_inst : _GEN_530 ? _slots_28_io_uop_edge_inst : _GEN_516 ? _slots_27_io_uop_edge_inst : _GEN_502 ? _slots_26_io_uop_edge_inst : _GEN_488 ? _slots_25_io_uop_edge_inst : _GEN_474 ? _slots_24_io_uop_edge_inst : _GEN_460 ? _slots_23_io_uop_edge_inst : _GEN_446 ? _slots_22_io_uop_edge_inst : _GEN_432 ? _slots_21_io_uop_edge_inst : _GEN_418 ? _slots_20_io_uop_edge_inst : _GEN_404 ? _slots_19_io_uop_edge_inst : _GEN_390 ? _slots_18_io_uop_edge_inst : _GEN_376 ? _slots_17_io_uop_edge_inst : _GEN_362 ? _slots_16_io_uop_edge_inst : _GEN_348 ? _slots_15_io_uop_edge_inst : _GEN_334 ? _slots_14_io_uop_edge_inst : _GEN_320 ? _slots_13_io_uop_edge_inst : _GEN_306 ? _slots_12_io_uop_edge_inst : _GEN_292 ? _slots_11_io_uop_edge_inst : _GEN_278 ? _slots_10_io_uop_edge_inst : _GEN_264 ? _slots_9_io_uop_edge_inst : _GEN_250 ? _slots_8_io_uop_edge_inst : _GEN_236 ? _slots_7_io_uop_edge_inst : _GEN_222 ? _slots_6_io_uop_edge_inst : _GEN_208 ? _slots_5_io_uop_edge_inst : _GEN_194 ? _slots_4_io_uop_edge_inst : _GEN_180 ? _slots_3_io_uop_edge_inst : _GEN_166 ? _slots_2_io_uop_edge_inst : _GEN_152 ? _slots_1_io_uop_edge_inst : _GEN_143 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_1_pc_lob = _GEN_679 ? _slots_39_io_uop_pc_lob : _GEN_669 ? _slots_38_io_uop_pc_lob : _GEN_656 ? _slots_37_io_uop_pc_lob : _GEN_642 ? _slots_36_io_uop_pc_lob : _GEN_628 ? _slots_35_io_uop_pc_lob : _GEN_614 ? _slots_34_io_uop_pc_lob : _GEN_600 ? _slots_33_io_uop_pc_lob : _GEN_586 ? _slots_32_io_uop_pc_lob : _GEN_572 ? _slots_31_io_uop_pc_lob : _GEN_558 ? _slots_30_io_uop_pc_lob : _GEN_544 ? _slots_29_io_uop_pc_lob : _GEN_530 ? _slots_28_io_uop_pc_lob : _GEN_516 ? _slots_27_io_uop_pc_lob : _GEN_502 ? _slots_26_io_uop_pc_lob : _GEN_488 ? _slots_25_io_uop_pc_lob : _GEN_474 ? _slots_24_io_uop_pc_lob : _GEN_460 ? _slots_23_io_uop_pc_lob : _GEN_446 ? _slots_22_io_uop_pc_lob : _GEN_432 ? _slots_21_io_uop_pc_lob : _GEN_418 ? _slots_20_io_uop_pc_lob : _GEN_404 ? _slots_19_io_uop_pc_lob : _GEN_390 ? _slots_18_io_uop_pc_lob : _GEN_376 ? _slots_17_io_uop_pc_lob : _GEN_362 ? _slots_16_io_uop_pc_lob : _GEN_348 ? _slots_15_io_uop_pc_lob : _GEN_334 ? _slots_14_io_uop_pc_lob : _GEN_320 ? _slots_13_io_uop_pc_lob : _GEN_306 ? _slots_12_io_uop_pc_lob : _GEN_292 ? _slots_11_io_uop_pc_lob : _GEN_278 ? _slots_10_io_uop_pc_lob : _GEN_264 ? _slots_9_io_uop_pc_lob : _GEN_250 ? _slots_8_io_uop_pc_lob : _GEN_236 ? _slots_7_io_uop_pc_lob : _GEN_222 ? _slots_6_io_uop_pc_lob : _GEN_208 ? _slots_5_io_uop_pc_lob : _GEN_194 ? _slots_4_io_uop_pc_lob : _GEN_180 ? _slots_3_io_uop_pc_lob : _GEN_166 ? _slots_2_io_uop_pc_lob : _GEN_152 ? _slots_1_io_uop_pc_lob : _GEN_143 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_1_taken = _GEN_679 ? _slots_39_io_uop_taken : _GEN_669 ? _slots_38_io_uop_taken : _GEN_656 ? _slots_37_io_uop_taken : _GEN_642 ? _slots_36_io_uop_taken : _GEN_628 ? _slots_35_io_uop_taken : _GEN_614 ? _slots_34_io_uop_taken : _GEN_600 ? _slots_33_io_uop_taken : _GEN_586 ? _slots_32_io_uop_taken : _GEN_572 ? _slots_31_io_uop_taken : _GEN_558 ? _slots_30_io_uop_taken : _GEN_544 ? _slots_29_io_uop_taken : _GEN_530 ? _slots_28_io_uop_taken : _GEN_516 ? _slots_27_io_uop_taken : _GEN_502 ? _slots_26_io_uop_taken : _GEN_488 ? _slots_25_io_uop_taken : _GEN_474 ? _slots_24_io_uop_taken : _GEN_460 ? _slots_23_io_uop_taken : _GEN_446 ? _slots_22_io_uop_taken : _GEN_432 ? _slots_21_io_uop_taken : _GEN_418 ? _slots_20_io_uop_taken : _GEN_404 ? _slots_19_io_uop_taken : _GEN_390 ? _slots_18_io_uop_taken : _GEN_376 ? _slots_17_io_uop_taken : _GEN_362 ? _slots_16_io_uop_taken : _GEN_348 ? _slots_15_io_uop_taken : _GEN_334 ? _slots_14_io_uop_taken : _GEN_320 ? _slots_13_io_uop_taken : _GEN_306 ? _slots_12_io_uop_taken : _GEN_292 ? _slots_11_io_uop_taken : _GEN_278 ? _slots_10_io_uop_taken : _GEN_264 ? _slots_9_io_uop_taken : _GEN_250 ? _slots_8_io_uop_taken : _GEN_236 ? _slots_7_io_uop_taken : _GEN_222 ? _slots_6_io_uop_taken : _GEN_208 ? _slots_5_io_uop_taken : _GEN_194 ? _slots_4_io_uop_taken : _GEN_180 ? _slots_3_io_uop_taken : _GEN_166 ? _slots_2_io_uop_taken : _GEN_152 ? _slots_1_io_uop_taken : _GEN_143 & _slots_0_io_uop_taken;
  assign io_iss_uops_1_imm_packed = _GEN_679 ? _slots_39_io_uop_imm_packed : _GEN_669 ? _slots_38_io_uop_imm_packed : _GEN_656 ? _slots_37_io_uop_imm_packed : _GEN_642 ? _slots_36_io_uop_imm_packed : _GEN_628 ? _slots_35_io_uop_imm_packed : _GEN_614 ? _slots_34_io_uop_imm_packed : _GEN_600 ? _slots_33_io_uop_imm_packed : _GEN_586 ? _slots_32_io_uop_imm_packed : _GEN_572 ? _slots_31_io_uop_imm_packed : _GEN_558 ? _slots_30_io_uop_imm_packed : _GEN_544 ? _slots_29_io_uop_imm_packed : _GEN_530 ? _slots_28_io_uop_imm_packed : _GEN_516 ? _slots_27_io_uop_imm_packed : _GEN_502 ? _slots_26_io_uop_imm_packed : _GEN_488 ? _slots_25_io_uop_imm_packed : _GEN_474 ? _slots_24_io_uop_imm_packed : _GEN_460 ? _slots_23_io_uop_imm_packed : _GEN_446 ? _slots_22_io_uop_imm_packed : _GEN_432 ? _slots_21_io_uop_imm_packed : _GEN_418 ? _slots_20_io_uop_imm_packed : _GEN_404 ? _slots_19_io_uop_imm_packed : _GEN_390 ? _slots_18_io_uop_imm_packed : _GEN_376 ? _slots_17_io_uop_imm_packed : _GEN_362 ? _slots_16_io_uop_imm_packed : _GEN_348 ? _slots_15_io_uop_imm_packed : _GEN_334 ? _slots_14_io_uop_imm_packed : _GEN_320 ? _slots_13_io_uop_imm_packed : _GEN_306 ? _slots_12_io_uop_imm_packed : _GEN_292 ? _slots_11_io_uop_imm_packed : _GEN_278 ? _slots_10_io_uop_imm_packed : _GEN_264 ? _slots_9_io_uop_imm_packed : _GEN_250 ? _slots_8_io_uop_imm_packed : _GEN_236 ? _slots_7_io_uop_imm_packed : _GEN_222 ? _slots_6_io_uop_imm_packed : _GEN_208 ? _slots_5_io_uop_imm_packed : _GEN_194 ? _slots_4_io_uop_imm_packed : _GEN_180 ? _slots_3_io_uop_imm_packed : _GEN_166 ? _slots_2_io_uop_imm_packed : _GEN_152 ? _slots_1_io_uop_imm_packed : _GEN_143 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_1_rob_idx = _GEN_679 ? _slots_39_io_uop_rob_idx : _GEN_669 ? _slots_38_io_uop_rob_idx : _GEN_656 ? _slots_37_io_uop_rob_idx : _GEN_642 ? _slots_36_io_uop_rob_idx : _GEN_628 ? _slots_35_io_uop_rob_idx : _GEN_614 ? _slots_34_io_uop_rob_idx : _GEN_600 ? _slots_33_io_uop_rob_idx : _GEN_586 ? _slots_32_io_uop_rob_idx : _GEN_572 ? _slots_31_io_uop_rob_idx : _GEN_558 ? _slots_30_io_uop_rob_idx : _GEN_544 ? _slots_29_io_uop_rob_idx : _GEN_530 ? _slots_28_io_uop_rob_idx : _GEN_516 ? _slots_27_io_uop_rob_idx : _GEN_502 ? _slots_26_io_uop_rob_idx : _GEN_488 ? _slots_25_io_uop_rob_idx : _GEN_474 ? _slots_24_io_uop_rob_idx : _GEN_460 ? _slots_23_io_uop_rob_idx : _GEN_446 ? _slots_22_io_uop_rob_idx : _GEN_432 ? _slots_21_io_uop_rob_idx : _GEN_418 ? _slots_20_io_uop_rob_idx : _GEN_404 ? _slots_19_io_uop_rob_idx : _GEN_390 ? _slots_18_io_uop_rob_idx : _GEN_376 ? _slots_17_io_uop_rob_idx : _GEN_362 ? _slots_16_io_uop_rob_idx : _GEN_348 ? _slots_15_io_uop_rob_idx : _GEN_334 ? _slots_14_io_uop_rob_idx : _GEN_320 ? _slots_13_io_uop_rob_idx : _GEN_306 ? _slots_12_io_uop_rob_idx : _GEN_292 ? _slots_11_io_uop_rob_idx : _GEN_278 ? _slots_10_io_uop_rob_idx : _GEN_264 ? _slots_9_io_uop_rob_idx : _GEN_250 ? _slots_8_io_uop_rob_idx : _GEN_236 ? _slots_7_io_uop_rob_idx : _GEN_222 ? _slots_6_io_uop_rob_idx : _GEN_208 ? _slots_5_io_uop_rob_idx : _GEN_194 ? _slots_4_io_uop_rob_idx : _GEN_180 ? _slots_3_io_uop_rob_idx : _GEN_166 ? _slots_2_io_uop_rob_idx : _GEN_152 ? _slots_1_io_uop_rob_idx : _GEN_143 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_1_ldq_idx = _GEN_679 ? _slots_39_io_uop_ldq_idx : _GEN_669 ? _slots_38_io_uop_ldq_idx : _GEN_656 ? _slots_37_io_uop_ldq_idx : _GEN_642 ? _slots_36_io_uop_ldq_idx : _GEN_628 ? _slots_35_io_uop_ldq_idx : _GEN_614 ? _slots_34_io_uop_ldq_idx : _GEN_600 ? _slots_33_io_uop_ldq_idx : _GEN_586 ? _slots_32_io_uop_ldq_idx : _GEN_572 ? _slots_31_io_uop_ldq_idx : _GEN_558 ? _slots_30_io_uop_ldq_idx : _GEN_544 ? _slots_29_io_uop_ldq_idx : _GEN_530 ? _slots_28_io_uop_ldq_idx : _GEN_516 ? _slots_27_io_uop_ldq_idx : _GEN_502 ? _slots_26_io_uop_ldq_idx : _GEN_488 ? _slots_25_io_uop_ldq_idx : _GEN_474 ? _slots_24_io_uop_ldq_idx : _GEN_460 ? _slots_23_io_uop_ldq_idx : _GEN_446 ? _slots_22_io_uop_ldq_idx : _GEN_432 ? _slots_21_io_uop_ldq_idx : _GEN_418 ? _slots_20_io_uop_ldq_idx : _GEN_404 ? _slots_19_io_uop_ldq_idx : _GEN_390 ? _slots_18_io_uop_ldq_idx : _GEN_376 ? _slots_17_io_uop_ldq_idx : _GEN_362 ? _slots_16_io_uop_ldq_idx : _GEN_348 ? _slots_15_io_uop_ldq_idx : _GEN_334 ? _slots_14_io_uop_ldq_idx : _GEN_320 ? _slots_13_io_uop_ldq_idx : _GEN_306 ? _slots_12_io_uop_ldq_idx : _GEN_292 ? _slots_11_io_uop_ldq_idx : _GEN_278 ? _slots_10_io_uop_ldq_idx : _GEN_264 ? _slots_9_io_uop_ldq_idx : _GEN_250 ? _slots_8_io_uop_ldq_idx : _GEN_236 ? _slots_7_io_uop_ldq_idx : _GEN_222 ? _slots_6_io_uop_ldq_idx : _GEN_208 ? _slots_5_io_uop_ldq_idx : _GEN_194 ? _slots_4_io_uop_ldq_idx : _GEN_180 ? _slots_3_io_uop_ldq_idx : _GEN_166 ? _slots_2_io_uop_ldq_idx : _GEN_152 ? _slots_1_io_uop_ldq_idx : _GEN_143 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_1_stq_idx = _GEN_679 ? _slots_39_io_uop_stq_idx : _GEN_669 ? _slots_38_io_uop_stq_idx : _GEN_656 ? _slots_37_io_uop_stq_idx : _GEN_642 ? _slots_36_io_uop_stq_idx : _GEN_628 ? _slots_35_io_uop_stq_idx : _GEN_614 ? _slots_34_io_uop_stq_idx : _GEN_600 ? _slots_33_io_uop_stq_idx : _GEN_586 ? _slots_32_io_uop_stq_idx : _GEN_572 ? _slots_31_io_uop_stq_idx : _GEN_558 ? _slots_30_io_uop_stq_idx : _GEN_544 ? _slots_29_io_uop_stq_idx : _GEN_530 ? _slots_28_io_uop_stq_idx : _GEN_516 ? _slots_27_io_uop_stq_idx : _GEN_502 ? _slots_26_io_uop_stq_idx : _GEN_488 ? _slots_25_io_uop_stq_idx : _GEN_474 ? _slots_24_io_uop_stq_idx : _GEN_460 ? _slots_23_io_uop_stq_idx : _GEN_446 ? _slots_22_io_uop_stq_idx : _GEN_432 ? _slots_21_io_uop_stq_idx : _GEN_418 ? _slots_20_io_uop_stq_idx : _GEN_404 ? _slots_19_io_uop_stq_idx : _GEN_390 ? _slots_18_io_uop_stq_idx : _GEN_376 ? _slots_17_io_uop_stq_idx : _GEN_362 ? _slots_16_io_uop_stq_idx : _GEN_348 ? _slots_15_io_uop_stq_idx : _GEN_334 ? _slots_14_io_uop_stq_idx : _GEN_320 ? _slots_13_io_uop_stq_idx : _GEN_306 ? _slots_12_io_uop_stq_idx : _GEN_292 ? _slots_11_io_uop_stq_idx : _GEN_278 ? _slots_10_io_uop_stq_idx : _GEN_264 ? _slots_9_io_uop_stq_idx : _GEN_250 ? _slots_8_io_uop_stq_idx : _GEN_236 ? _slots_7_io_uop_stq_idx : _GEN_222 ? _slots_6_io_uop_stq_idx : _GEN_208 ? _slots_5_io_uop_stq_idx : _GEN_194 ? _slots_4_io_uop_stq_idx : _GEN_180 ? _slots_3_io_uop_stq_idx : _GEN_166 ? _slots_2_io_uop_stq_idx : _GEN_152 ? _slots_1_io_uop_stq_idx : _GEN_143 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_1_pdst = _GEN_679 ? _slots_39_io_uop_pdst : _GEN_669 ? _slots_38_io_uop_pdst : _GEN_656 ? _slots_37_io_uop_pdst : _GEN_642 ? _slots_36_io_uop_pdst : _GEN_628 ? _slots_35_io_uop_pdst : _GEN_614 ? _slots_34_io_uop_pdst : _GEN_600 ? _slots_33_io_uop_pdst : _GEN_586 ? _slots_32_io_uop_pdst : _GEN_572 ? _slots_31_io_uop_pdst : _GEN_558 ? _slots_30_io_uop_pdst : _GEN_544 ? _slots_29_io_uop_pdst : _GEN_530 ? _slots_28_io_uop_pdst : _GEN_516 ? _slots_27_io_uop_pdst : _GEN_502 ? _slots_26_io_uop_pdst : _GEN_488 ? _slots_25_io_uop_pdst : _GEN_474 ? _slots_24_io_uop_pdst : _GEN_460 ? _slots_23_io_uop_pdst : _GEN_446 ? _slots_22_io_uop_pdst : _GEN_432 ? _slots_21_io_uop_pdst : _GEN_418 ? _slots_20_io_uop_pdst : _GEN_404 ? _slots_19_io_uop_pdst : _GEN_390 ? _slots_18_io_uop_pdst : _GEN_376 ? _slots_17_io_uop_pdst : _GEN_362 ? _slots_16_io_uop_pdst : _GEN_348 ? _slots_15_io_uop_pdst : _GEN_334 ? _slots_14_io_uop_pdst : _GEN_320 ? _slots_13_io_uop_pdst : _GEN_306 ? _slots_12_io_uop_pdst : _GEN_292 ? _slots_11_io_uop_pdst : _GEN_278 ? _slots_10_io_uop_pdst : _GEN_264 ? _slots_9_io_uop_pdst : _GEN_250 ? _slots_8_io_uop_pdst : _GEN_236 ? _slots_7_io_uop_pdst : _GEN_222 ? _slots_6_io_uop_pdst : _GEN_208 ? _slots_5_io_uop_pdst : _GEN_194 ? _slots_4_io_uop_pdst : _GEN_180 ? _slots_3_io_uop_pdst : _GEN_166 ? _slots_2_io_uop_pdst : _GEN_152 ? _slots_1_io_uop_pdst : _GEN_143 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_1_prs1 = _GEN_679 ? _slots_39_io_uop_prs1 : _GEN_669 ? _slots_38_io_uop_prs1 : _GEN_656 ? _slots_37_io_uop_prs1 : _GEN_642 ? _slots_36_io_uop_prs1 : _GEN_628 ? _slots_35_io_uop_prs1 : _GEN_614 ? _slots_34_io_uop_prs1 : _GEN_600 ? _slots_33_io_uop_prs1 : _GEN_586 ? _slots_32_io_uop_prs1 : _GEN_572 ? _slots_31_io_uop_prs1 : _GEN_558 ? _slots_30_io_uop_prs1 : _GEN_544 ? _slots_29_io_uop_prs1 : _GEN_530 ? _slots_28_io_uop_prs1 : _GEN_516 ? _slots_27_io_uop_prs1 : _GEN_502 ? _slots_26_io_uop_prs1 : _GEN_488 ? _slots_25_io_uop_prs1 : _GEN_474 ? _slots_24_io_uop_prs1 : _GEN_460 ? _slots_23_io_uop_prs1 : _GEN_446 ? _slots_22_io_uop_prs1 : _GEN_432 ? _slots_21_io_uop_prs1 : _GEN_418 ? _slots_20_io_uop_prs1 : _GEN_404 ? _slots_19_io_uop_prs1 : _GEN_390 ? _slots_18_io_uop_prs1 : _GEN_376 ? _slots_17_io_uop_prs1 : _GEN_362 ? _slots_16_io_uop_prs1 : _GEN_348 ? _slots_15_io_uop_prs1 : _GEN_334 ? _slots_14_io_uop_prs1 : _GEN_320 ? _slots_13_io_uop_prs1 : _GEN_306 ? _slots_12_io_uop_prs1 : _GEN_292 ? _slots_11_io_uop_prs1 : _GEN_278 ? _slots_10_io_uop_prs1 : _GEN_264 ? _slots_9_io_uop_prs1 : _GEN_250 ? _slots_8_io_uop_prs1 : _GEN_236 ? _slots_7_io_uop_prs1 : _GEN_222 ? _slots_6_io_uop_prs1 : _GEN_208 ? _slots_5_io_uop_prs1 : _GEN_194 ? _slots_4_io_uop_prs1 : _GEN_180 ? _slots_3_io_uop_prs1 : _GEN_166 ? _slots_2_io_uop_prs1 : _GEN_152 ? _slots_1_io_uop_prs1 : _GEN_143 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_1_prs2 = _GEN_679 ? _slots_39_io_uop_prs2 : _GEN_669 ? _slots_38_io_uop_prs2 : _GEN_656 ? _slots_37_io_uop_prs2 : _GEN_642 ? _slots_36_io_uop_prs2 : _GEN_628 ? _slots_35_io_uop_prs2 : _GEN_614 ? _slots_34_io_uop_prs2 : _GEN_600 ? _slots_33_io_uop_prs2 : _GEN_586 ? _slots_32_io_uop_prs2 : _GEN_572 ? _slots_31_io_uop_prs2 : _GEN_558 ? _slots_30_io_uop_prs2 : _GEN_544 ? _slots_29_io_uop_prs2 : _GEN_530 ? _slots_28_io_uop_prs2 : _GEN_516 ? _slots_27_io_uop_prs2 : _GEN_502 ? _slots_26_io_uop_prs2 : _GEN_488 ? _slots_25_io_uop_prs2 : _GEN_474 ? _slots_24_io_uop_prs2 : _GEN_460 ? _slots_23_io_uop_prs2 : _GEN_446 ? _slots_22_io_uop_prs2 : _GEN_432 ? _slots_21_io_uop_prs2 : _GEN_418 ? _slots_20_io_uop_prs2 : _GEN_404 ? _slots_19_io_uop_prs2 : _GEN_390 ? _slots_18_io_uop_prs2 : _GEN_376 ? _slots_17_io_uop_prs2 : _GEN_362 ? _slots_16_io_uop_prs2 : _GEN_348 ? _slots_15_io_uop_prs2 : _GEN_334 ? _slots_14_io_uop_prs2 : _GEN_320 ? _slots_13_io_uop_prs2 : _GEN_306 ? _slots_12_io_uop_prs2 : _GEN_292 ? _slots_11_io_uop_prs2 : _GEN_278 ? _slots_10_io_uop_prs2 : _GEN_264 ? _slots_9_io_uop_prs2 : _GEN_250 ? _slots_8_io_uop_prs2 : _GEN_236 ? _slots_7_io_uop_prs2 : _GEN_222 ? _slots_6_io_uop_prs2 : _GEN_208 ? _slots_5_io_uop_prs2 : _GEN_194 ? _slots_4_io_uop_prs2 : _GEN_180 ? _slots_3_io_uop_prs2 : _GEN_166 ? _slots_2_io_uop_prs2 : _GEN_152 ? _slots_1_io_uop_prs2 : _GEN_143 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_1_bypassable = _GEN_679 ? _slots_39_io_uop_bypassable : _GEN_669 ? _slots_38_io_uop_bypassable : _GEN_656 ? _slots_37_io_uop_bypassable : _GEN_642 ? _slots_36_io_uop_bypassable : _GEN_628 ? _slots_35_io_uop_bypassable : _GEN_614 ? _slots_34_io_uop_bypassable : _GEN_600 ? _slots_33_io_uop_bypassable : _GEN_586 ? _slots_32_io_uop_bypassable : _GEN_572 ? _slots_31_io_uop_bypassable : _GEN_558 ? _slots_30_io_uop_bypassable : _GEN_544 ? _slots_29_io_uop_bypassable : _GEN_530 ? _slots_28_io_uop_bypassable : _GEN_516 ? _slots_27_io_uop_bypassable : _GEN_502 ? _slots_26_io_uop_bypassable : _GEN_488 ? _slots_25_io_uop_bypassable : _GEN_474 ? _slots_24_io_uop_bypassable : _GEN_460 ? _slots_23_io_uop_bypassable : _GEN_446 ? _slots_22_io_uop_bypassable : _GEN_432 ? _slots_21_io_uop_bypassable : _GEN_418 ? _slots_20_io_uop_bypassable : _GEN_404 ? _slots_19_io_uop_bypassable : _GEN_390 ? _slots_18_io_uop_bypassable : _GEN_376 ? _slots_17_io_uop_bypassable : _GEN_362 ? _slots_16_io_uop_bypassable : _GEN_348 ? _slots_15_io_uop_bypassable : _GEN_334 ? _slots_14_io_uop_bypassable : _GEN_320 ? _slots_13_io_uop_bypassable : _GEN_306 ? _slots_12_io_uop_bypassable : _GEN_292 ? _slots_11_io_uop_bypassable : _GEN_278 ? _slots_10_io_uop_bypassable : _GEN_264 ? _slots_9_io_uop_bypassable : _GEN_250 ? _slots_8_io_uop_bypassable : _GEN_236 ? _slots_7_io_uop_bypassable : _GEN_222 ? _slots_6_io_uop_bypassable : _GEN_208 ? _slots_5_io_uop_bypassable : _GEN_194 ? _slots_4_io_uop_bypassable : _GEN_180 ? _slots_3_io_uop_bypassable : _GEN_166 ? _slots_2_io_uop_bypassable : _GEN_152 ? _slots_1_io_uop_bypassable : _GEN_143 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_1_mem_cmd = _GEN_679 ? _slots_39_io_uop_mem_cmd : _GEN_669 ? _slots_38_io_uop_mem_cmd : _GEN_656 ? _slots_37_io_uop_mem_cmd : _GEN_642 ? _slots_36_io_uop_mem_cmd : _GEN_628 ? _slots_35_io_uop_mem_cmd : _GEN_614 ? _slots_34_io_uop_mem_cmd : _GEN_600 ? _slots_33_io_uop_mem_cmd : _GEN_586 ? _slots_32_io_uop_mem_cmd : _GEN_572 ? _slots_31_io_uop_mem_cmd : _GEN_558 ? _slots_30_io_uop_mem_cmd : _GEN_544 ? _slots_29_io_uop_mem_cmd : _GEN_530 ? _slots_28_io_uop_mem_cmd : _GEN_516 ? _slots_27_io_uop_mem_cmd : _GEN_502 ? _slots_26_io_uop_mem_cmd : _GEN_488 ? _slots_25_io_uop_mem_cmd : _GEN_474 ? _slots_24_io_uop_mem_cmd : _GEN_460 ? _slots_23_io_uop_mem_cmd : _GEN_446 ? _slots_22_io_uop_mem_cmd : _GEN_432 ? _slots_21_io_uop_mem_cmd : _GEN_418 ? _slots_20_io_uop_mem_cmd : _GEN_404 ? _slots_19_io_uop_mem_cmd : _GEN_390 ? _slots_18_io_uop_mem_cmd : _GEN_376 ? _slots_17_io_uop_mem_cmd : _GEN_362 ? _slots_16_io_uop_mem_cmd : _GEN_348 ? _slots_15_io_uop_mem_cmd : _GEN_334 ? _slots_14_io_uop_mem_cmd : _GEN_320 ? _slots_13_io_uop_mem_cmd : _GEN_306 ? _slots_12_io_uop_mem_cmd : _GEN_292 ? _slots_11_io_uop_mem_cmd : _GEN_278 ? _slots_10_io_uop_mem_cmd : _GEN_264 ? _slots_9_io_uop_mem_cmd : _GEN_250 ? _slots_8_io_uop_mem_cmd : _GEN_236 ? _slots_7_io_uop_mem_cmd : _GEN_222 ? _slots_6_io_uop_mem_cmd : _GEN_208 ? _slots_5_io_uop_mem_cmd : _GEN_194 ? _slots_4_io_uop_mem_cmd : _GEN_180 ? _slots_3_io_uop_mem_cmd : _GEN_166 ? _slots_2_io_uop_mem_cmd : _GEN_152 ? _slots_1_io_uop_mem_cmd : _GEN_143 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_1_is_amo = _GEN_679 ? _slots_39_io_uop_is_amo : _GEN_669 ? _slots_38_io_uop_is_amo : _GEN_656 ? _slots_37_io_uop_is_amo : _GEN_642 ? _slots_36_io_uop_is_amo : _GEN_628 ? _slots_35_io_uop_is_amo : _GEN_614 ? _slots_34_io_uop_is_amo : _GEN_600 ? _slots_33_io_uop_is_amo : _GEN_586 ? _slots_32_io_uop_is_amo : _GEN_572 ? _slots_31_io_uop_is_amo : _GEN_558 ? _slots_30_io_uop_is_amo : _GEN_544 ? _slots_29_io_uop_is_amo : _GEN_530 ? _slots_28_io_uop_is_amo : _GEN_516 ? _slots_27_io_uop_is_amo : _GEN_502 ? _slots_26_io_uop_is_amo : _GEN_488 ? _slots_25_io_uop_is_amo : _GEN_474 ? _slots_24_io_uop_is_amo : _GEN_460 ? _slots_23_io_uop_is_amo : _GEN_446 ? _slots_22_io_uop_is_amo : _GEN_432 ? _slots_21_io_uop_is_amo : _GEN_418 ? _slots_20_io_uop_is_amo : _GEN_404 ? _slots_19_io_uop_is_amo : _GEN_390 ? _slots_18_io_uop_is_amo : _GEN_376 ? _slots_17_io_uop_is_amo : _GEN_362 ? _slots_16_io_uop_is_amo : _GEN_348 ? _slots_15_io_uop_is_amo : _GEN_334 ? _slots_14_io_uop_is_amo : _GEN_320 ? _slots_13_io_uop_is_amo : _GEN_306 ? _slots_12_io_uop_is_amo : _GEN_292 ? _slots_11_io_uop_is_amo : _GEN_278 ? _slots_10_io_uop_is_amo : _GEN_264 ? _slots_9_io_uop_is_amo : _GEN_250 ? _slots_8_io_uop_is_amo : _GEN_236 ? _slots_7_io_uop_is_amo : _GEN_222 ? _slots_6_io_uop_is_amo : _GEN_208 ? _slots_5_io_uop_is_amo : _GEN_194 ? _slots_4_io_uop_is_amo : _GEN_180 ? _slots_3_io_uop_is_amo : _GEN_166 ? _slots_2_io_uop_is_amo : _GEN_152 ? _slots_1_io_uop_is_amo : _GEN_143 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_1_uses_stq = _GEN_679 ? _slots_39_io_uop_uses_stq : _GEN_669 ? _slots_38_io_uop_uses_stq : _GEN_656 ? _slots_37_io_uop_uses_stq : _GEN_642 ? _slots_36_io_uop_uses_stq : _GEN_628 ? _slots_35_io_uop_uses_stq : _GEN_614 ? _slots_34_io_uop_uses_stq : _GEN_600 ? _slots_33_io_uop_uses_stq : _GEN_586 ? _slots_32_io_uop_uses_stq : _GEN_572 ? _slots_31_io_uop_uses_stq : _GEN_558 ? _slots_30_io_uop_uses_stq : _GEN_544 ? _slots_29_io_uop_uses_stq : _GEN_530 ? _slots_28_io_uop_uses_stq : _GEN_516 ? _slots_27_io_uop_uses_stq : _GEN_502 ? _slots_26_io_uop_uses_stq : _GEN_488 ? _slots_25_io_uop_uses_stq : _GEN_474 ? _slots_24_io_uop_uses_stq : _GEN_460 ? _slots_23_io_uop_uses_stq : _GEN_446 ? _slots_22_io_uop_uses_stq : _GEN_432 ? _slots_21_io_uop_uses_stq : _GEN_418 ? _slots_20_io_uop_uses_stq : _GEN_404 ? _slots_19_io_uop_uses_stq : _GEN_390 ? _slots_18_io_uop_uses_stq : _GEN_376 ? _slots_17_io_uop_uses_stq : _GEN_362 ? _slots_16_io_uop_uses_stq : _GEN_348 ? _slots_15_io_uop_uses_stq : _GEN_334 ? _slots_14_io_uop_uses_stq : _GEN_320 ? _slots_13_io_uop_uses_stq : _GEN_306 ? _slots_12_io_uop_uses_stq : _GEN_292 ? _slots_11_io_uop_uses_stq : _GEN_278 ? _slots_10_io_uop_uses_stq : _GEN_264 ? _slots_9_io_uop_uses_stq : _GEN_250 ? _slots_8_io_uop_uses_stq : _GEN_236 ? _slots_7_io_uop_uses_stq : _GEN_222 ? _slots_6_io_uop_uses_stq : _GEN_208 ? _slots_5_io_uop_uses_stq : _GEN_194 ? _slots_4_io_uop_uses_stq : _GEN_180 ? _slots_3_io_uop_uses_stq : _GEN_166 ? _slots_2_io_uop_uses_stq : _GEN_152 ? _slots_1_io_uop_uses_stq : _GEN_143 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_1_ldst_val = _GEN_679 ? _slots_39_io_uop_ldst_val : _GEN_669 ? _slots_38_io_uop_ldst_val : _GEN_656 ? _slots_37_io_uop_ldst_val : _GEN_642 ? _slots_36_io_uop_ldst_val : _GEN_628 ? _slots_35_io_uop_ldst_val : _GEN_614 ? _slots_34_io_uop_ldst_val : _GEN_600 ? _slots_33_io_uop_ldst_val : _GEN_586 ? _slots_32_io_uop_ldst_val : _GEN_572 ? _slots_31_io_uop_ldst_val : _GEN_558 ? _slots_30_io_uop_ldst_val : _GEN_544 ? _slots_29_io_uop_ldst_val : _GEN_530 ? _slots_28_io_uop_ldst_val : _GEN_516 ? _slots_27_io_uop_ldst_val : _GEN_502 ? _slots_26_io_uop_ldst_val : _GEN_488 ? _slots_25_io_uop_ldst_val : _GEN_474 ? _slots_24_io_uop_ldst_val : _GEN_460 ? _slots_23_io_uop_ldst_val : _GEN_446 ? _slots_22_io_uop_ldst_val : _GEN_432 ? _slots_21_io_uop_ldst_val : _GEN_418 ? _slots_20_io_uop_ldst_val : _GEN_404 ? _slots_19_io_uop_ldst_val : _GEN_390 ? _slots_18_io_uop_ldst_val : _GEN_376 ? _slots_17_io_uop_ldst_val : _GEN_362 ? _slots_16_io_uop_ldst_val : _GEN_348 ? _slots_15_io_uop_ldst_val : _GEN_334 ? _slots_14_io_uop_ldst_val : _GEN_320 ? _slots_13_io_uop_ldst_val : _GEN_306 ? _slots_12_io_uop_ldst_val : _GEN_292 ? _slots_11_io_uop_ldst_val : _GEN_278 ? _slots_10_io_uop_ldst_val : _GEN_264 ? _slots_9_io_uop_ldst_val : _GEN_250 ? _slots_8_io_uop_ldst_val : _GEN_236 ? _slots_7_io_uop_ldst_val : _GEN_222 ? _slots_6_io_uop_ldst_val : _GEN_208 ? _slots_5_io_uop_ldst_val : _GEN_194 ? _slots_4_io_uop_ldst_val : _GEN_180 ? _slots_3_io_uop_ldst_val : _GEN_166 ? _slots_2_io_uop_ldst_val : _GEN_152 ? _slots_1_io_uop_ldst_val : _GEN_143 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_1_dst_rtype = _GEN_679 ? _slots_39_io_uop_dst_rtype : _GEN_669 ? _slots_38_io_uop_dst_rtype : _GEN_656 ? _slots_37_io_uop_dst_rtype : _GEN_642 ? _slots_36_io_uop_dst_rtype : _GEN_628 ? _slots_35_io_uop_dst_rtype : _GEN_614 ? _slots_34_io_uop_dst_rtype : _GEN_600 ? _slots_33_io_uop_dst_rtype : _GEN_586 ? _slots_32_io_uop_dst_rtype : _GEN_572 ? _slots_31_io_uop_dst_rtype : _GEN_558 ? _slots_30_io_uop_dst_rtype : _GEN_544 ? _slots_29_io_uop_dst_rtype : _GEN_530 ? _slots_28_io_uop_dst_rtype : _GEN_516 ? _slots_27_io_uop_dst_rtype : _GEN_502 ? _slots_26_io_uop_dst_rtype : _GEN_488 ? _slots_25_io_uop_dst_rtype : _GEN_474 ? _slots_24_io_uop_dst_rtype : _GEN_460 ? _slots_23_io_uop_dst_rtype : _GEN_446 ? _slots_22_io_uop_dst_rtype : _GEN_432 ? _slots_21_io_uop_dst_rtype : _GEN_418 ? _slots_20_io_uop_dst_rtype : _GEN_404 ? _slots_19_io_uop_dst_rtype : _GEN_390 ? _slots_18_io_uop_dst_rtype : _GEN_376 ? _slots_17_io_uop_dst_rtype : _GEN_362 ? _slots_16_io_uop_dst_rtype : _GEN_348 ? _slots_15_io_uop_dst_rtype : _GEN_334 ? _slots_14_io_uop_dst_rtype : _GEN_320 ? _slots_13_io_uop_dst_rtype : _GEN_306 ? _slots_12_io_uop_dst_rtype : _GEN_292 ? _slots_11_io_uop_dst_rtype : _GEN_278 ? _slots_10_io_uop_dst_rtype : _GEN_264 ? _slots_9_io_uop_dst_rtype : _GEN_250 ? _slots_8_io_uop_dst_rtype : _GEN_236 ? _slots_7_io_uop_dst_rtype : _GEN_222 ? _slots_6_io_uop_dst_rtype : _GEN_208 ? _slots_5_io_uop_dst_rtype : _GEN_194 ? _slots_4_io_uop_dst_rtype : _GEN_180 ? _slots_3_io_uop_dst_rtype : _GEN_166 ? _slots_2_io_uop_dst_rtype : _GEN_152 ? _slots_1_io_uop_dst_rtype : _GEN_143 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_1_lrs1_rtype = _GEN_679 ? _slots_39_io_uop_lrs1_rtype : _GEN_669 ? _slots_38_io_uop_lrs1_rtype : _GEN_656 ? _slots_37_io_uop_lrs1_rtype : _GEN_642 ? _slots_36_io_uop_lrs1_rtype : _GEN_628 ? _slots_35_io_uop_lrs1_rtype : _GEN_614 ? _slots_34_io_uop_lrs1_rtype : _GEN_600 ? _slots_33_io_uop_lrs1_rtype : _GEN_586 ? _slots_32_io_uop_lrs1_rtype : _GEN_572 ? _slots_31_io_uop_lrs1_rtype : _GEN_558 ? _slots_30_io_uop_lrs1_rtype : _GEN_544 ? _slots_29_io_uop_lrs1_rtype : _GEN_530 ? _slots_28_io_uop_lrs1_rtype : _GEN_516 ? _slots_27_io_uop_lrs1_rtype : _GEN_502 ? _slots_26_io_uop_lrs1_rtype : _GEN_488 ? _slots_25_io_uop_lrs1_rtype : _GEN_474 ? _slots_24_io_uop_lrs1_rtype : _GEN_460 ? _slots_23_io_uop_lrs1_rtype : _GEN_446 ? _slots_22_io_uop_lrs1_rtype : _GEN_432 ? _slots_21_io_uop_lrs1_rtype : _GEN_418 ? _slots_20_io_uop_lrs1_rtype : _GEN_404 ? _slots_19_io_uop_lrs1_rtype : _GEN_390 ? _slots_18_io_uop_lrs1_rtype : _GEN_376 ? _slots_17_io_uop_lrs1_rtype : _GEN_362 ? _slots_16_io_uop_lrs1_rtype : _GEN_348 ? _slots_15_io_uop_lrs1_rtype : _GEN_334 ? _slots_14_io_uop_lrs1_rtype : _GEN_320 ? _slots_13_io_uop_lrs1_rtype : _GEN_306 ? _slots_12_io_uop_lrs1_rtype : _GEN_292 ? _slots_11_io_uop_lrs1_rtype : _GEN_278 ? _slots_10_io_uop_lrs1_rtype : _GEN_264 ? _slots_9_io_uop_lrs1_rtype : _GEN_250 ? _slots_8_io_uop_lrs1_rtype : _GEN_236 ? _slots_7_io_uop_lrs1_rtype : _GEN_222 ? _slots_6_io_uop_lrs1_rtype : _GEN_208 ? _slots_5_io_uop_lrs1_rtype : _GEN_194 ? _slots_4_io_uop_lrs1_rtype : _GEN_180 ? _slots_3_io_uop_lrs1_rtype : _GEN_166 ? _slots_2_io_uop_lrs1_rtype : _GEN_152 ? _slots_1_io_uop_lrs1_rtype : _GEN_143 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_1_lrs2_rtype = _GEN_679 ? _slots_39_io_uop_lrs2_rtype : _GEN_669 ? _slots_38_io_uop_lrs2_rtype : _GEN_656 ? _slots_37_io_uop_lrs2_rtype : _GEN_642 ? _slots_36_io_uop_lrs2_rtype : _GEN_628 ? _slots_35_io_uop_lrs2_rtype : _GEN_614 ? _slots_34_io_uop_lrs2_rtype : _GEN_600 ? _slots_33_io_uop_lrs2_rtype : _GEN_586 ? _slots_32_io_uop_lrs2_rtype : _GEN_572 ? _slots_31_io_uop_lrs2_rtype : _GEN_558 ? _slots_30_io_uop_lrs2_rtype : _GEN_544 ? _slots_29_io_uop_lrs2_rtype : _GEN_530 ? _slots_28_io_uop_lrs2_rtype : _GEN_516 ? _slots_27_io_uop_lrs2_rtype : _GEN_502 ? _slots_26_io_uop_lrs2_rtype : _GEN_488 ? _slots_25_io_uop_lrs2_rtype : _GEN_474 ? _slots_24_io_uop_lrs2_rtype : _GEN_460 ? _slots_23_io_uop_lrs2_rtype : _GEN_446 ? _slots_22_io_uop_lrs2_rtype : _GEN_432 ? _slots_21_io_uop_lrs2_rtype : _GEN_418 ? _slots_20_io_uop_lrs2_rtype : _GEN_404 ? _slots_19_io_uop_lrs2_rtype : _GEN_390 ? _slots_18_io_uop_lrs2_rtype : _GEN_376 ? _slots_17_io_uop_lrs2_rtype : _GEN_362 ? _slots_16_io_uop_lrs2_rtype : _GEN_348 ? _slots_15_io_uop_lrs2_rtype : _GEN_334 ? _slots_14_io_uop_lrs2_rtype : _GEN_320 ? _slots_13_io_uop_lrs2_rtype : _GEN_306 ? _slots_12_io_uop_lrs2_rtype : _GEN_292 ? _slots_11_io_uop_lrs2_rtype : _GEN_278 ? _slots_10_io_uop_lrs2_rtype : _GEN_264 ? _slots_9_io_uop_lrs2_rtype : _GEN_250 ? _slots_8_io_uop_lrs2_rtype : _GEN_236 ? _slots_7_io_uop_lrs2_rtype : _GEN_222 ? _slots_6_io_uop_lrs2_rtype : _GEN_208 ? _slots_5_io_uop_lrs2_rtype : _GEN_194 ? _slots_4_io_uop_lrs2_rtype : _GEN_180 ? _slots_3_io_uop_lrs2_rtype : _GEN_166 ? _slots_2_io_uop_lrs2_rtype : _GEN_152 ? _slots_1_io_uop_lrs2_rtype : _GEN_143 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_2_uopc = _GEN_681 ? _slots_39_io_uop_uopc : _GEN_673 ? _slots_38_io_uop_uopc : _GEN_660 ? _slots_37_io_uop_uopc : _GEN_646 ? _slots_36_io_uop_uopc : _GEN_632 ? _slots_35_io_uop_uopc : _GEN_618 ? _slots_34_io_uop_uopc : _GEN_604 ? _slots_33_io_uop_uopc : _GEN_590 ? _slots_32_io_uop_uopc : _GEN_576 ? _slots_31_io_uop_uopc : _GEN_562 ? _slots_30_io_uop_uopc : _GEN_548 ? _slots_29_io_uop_uopc : _GEN_534 ? _slots_28_io_uop_uopc : _GEN_520 ? _slots_27_io_uop_uopc : _GEN_506 ? _slots_26_io_uop_uopc : _GEN_492 ? _slots_25_io_uop_uopc : _GEN_478 ? _slots_24_io_uop_uopc : _GEN_464 ? _slots_23_io_uop_uopc : _GEN_450 ? _slots_22_io_uop_uopc : _GEN_436 ? _slots_21_io_uop_uopc : _GEN_422 ? _slots_20_io_uop_uopc : _GEN_408 ? _slots_19_io_uop_uopc : _GEN_394 ? _slots_18_io_uop_uopc : _GEN_380 ? _slots_17_io_uop_uopc : _GEN_366 ? _slots_16_io_uop_uopc : _GEN_352 ? _slots_15_io_uop_uopc : _GEN_338 ? _slots_14_io_uop_uopc : _GEN_324 ? _slots_13_io_uop_uopc : _GEN_310 ? _slots_12_io_uop_uopc : _GEN_296 ? _slots_11_io_uop_uopc : _GEN_282 ? _slots_10_io_uop_uopc : _GEN_268 ? _slots_9_io_uop_uopc : _GEN_254 ? _slots_8_io_uop_uopc : _GEN_240 ? _slots_7_io_uop_uopc : _GEN_226 ? _slots_6_io_uop_uopc : _GEN_212 ? _slots_5_io_uop_uopc : _GEN_198 ? _slots_4_io_uop_uopc : _GEN_184 ? _slots_3_io_uop_uopc : _GEN_170 ? _slots_2_io_uop_uopc : _GEN_156 ? _slots_1_io_uop_uopc : _GEN_145 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_2_is_rvc = _GEN_681 ? _slots_39_io_uop_is_rvc : _GEN_673 ? _slots_38_io_uop_is_rvc : _GEN_660 ? _slots_37_io_uop_is_rvc : _GEN_646 ? _slots_36_io_uop_is_rvc : _GEN_632 ? _slots_35_io_uop_is_rvc : _GEN_618 ? _slots_34_io_uop_is_rvc : _GEN_604 ? _slots_33_io_uop_is_rvc : _GEN_590 ? _slots_32_io_uop_is_rvc : _GEN_576 ? _slots_31_io_uop_is_rvc : _GEN_562 ? _slots_30_io_uop_is_rvc : _GEN_548 ? _slots_29_io_uop_is_rvc : _GEN_534 ? _slots_28_io_uop_is_rvc : _GEN_520 ? _slots_27_io_uop_is_rvc : _GEN_506 ? _slots_26_io_uop_is_rvc : _GEN_492 ? _slots_25_io_uop_is_rvc : _GEN_478 ? _slots_24_io_uop_is_rvc : _GEN_464 ? _slots_23_io_uop_is_rvc : _GEN_450 ? _slots_22_io_uop_is_rvc : _GEN_436 ? _slots_21_io_uop_is_rvc : _GEN_422 ? _slots_20_io_uop_is_rvc : _GEN_408 ? _slots_19_io_uop_is_rvc : _GEN_394 ? _slots_18_io_uop_is_rvc : _GEN_380 ? _slots_17_io_uop_is_rvc : _GEN_366 ? _slots_16_io_uop_is_rvc : _GEN_352 ? _slots_15_io_uop_is_rvc : _GEN_338 ? _slots_14_io_uop_is_rvc : _GEN_324 ? _slots_13_io_uop_is_rvc : _GEN_310 ? _slots_12_io_uop_is_rvc : _GEN_296 ? _slots_11_io_uop_is_rvc : _GEN_282 ? _slots_10_io_uop_is_rvc : _GEN_268 ? _slots_9_io_uop_is_rvc : _GEN_254 ? _slots_8_io_uop_is_rvc : _GEN_240 ? _slots_7_io_uop_is_rvc : _GEN_226 ? _slots_6_io_uop_is_rvc : _GEN_212 ? _slots_5_io_uop_is_rvc : _GEN_198 ? _slots_4_io_uop_is_rvc : _GEN_184 ? _slots_3_io_uop_is_rvc : _GEN_170 ? _slots_2_io_uop_is_rvc : _GEN_156 ? _slots_1_io_uop_is_rvc : _GEN_145 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_2_fu_code = _GEN_681 ? _slots_39_io_uop_fu_code : _GEN_673 ? _slots_38_io_uop_fu_code : _GEN_660 ? _slots_37_io_uop_fu_code : _GEN_646 ? _slots_36_io_uop_fu_code : _GEN_632 ? _slots_35_io_uop_fu_code : _GEN_618 ? _slots_34_io_uop_fu_code : _GEN_604 ? _slots_33_io_uop_fu_code : _GEN_590 ? _slots_32_io_uop_fu_code : _GEN_576 ? _slots_31_io_uop_fu_code : _GEN_562 ? _slots_30_io_uop_fu_code : _GEN_548 ? _slots_29_io_uop_fu_code : _GEN_534 ? _slots_28_io_uop_fu_code : _GEN_520 ? _slots_27_io_uop_fu_code : _GEN_506 ? _slots_26_io_uop_fu_code : _GEN_492 ? _slots_25_io_uop_fu_code : _GEN_478 ? _slots_24_io_uop_fu_code : _GEN_464 ? _slots_23_io_uop_fu_code : _GEN_450 ? _slots_22_io_uop_fu_code : _GEN_436 ? _slots_21_io_uop_fu_code : _GEN_422 ? _slots_20_io_uop_fu_code : _GEN_408 ? _slots_19_io_uop_fu_code : _GEN_394 ? _slots_18_io_uop_fu_code : _GEN_380 ? _slots_17_io_uop_fu_code : _GEN_366 ? _slots_16_io_uop_fu_code : _GEN_352 ? _slots_15_io_uop_fu_code : _GEN_338 ? _slots_14_io_uop_fu_code : _GEN_324 ? _slots_13_io_uop_fu_code : _GEN_310 ? _slots_12_io_uop_fu_code : _GEN_296 ? _slots_11_io_uop_fu_code : _GEN_282 ? _slots_10_io_uop_fu_code : _GEN_268 ? _slots_9_io_uop_fu_code : _GEN_254 ? _slots_8_io_uop_fu_code : _GEN_240 ? _slots_7_io_uop_fu_code : _GEN_226 ? _slots_6_io_uop_fu_code : _GEN_212 ? _slots_5_io_uop_fu_code : _GEN_198 ? _slots_4_io_uop_fu_code : _GEN_184 ? _slots_3_io_uop_fu_code : _GEN_170 ? _slots_2_io_uop_fu_code : _GEN_156 ? _slots_1_io_uop_fu_code : _GEN_145 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_2_iw_p1_poisoned = _GEN_681 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_673 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_660 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_646 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_632 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_618 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_604 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_590 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_576 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_562 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_548 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_534 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_520 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_506 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_492 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_478 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_464 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_450 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_436 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_422 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_408 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_394 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_380 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_366 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_352 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_338 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_324 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_310 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_296 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_282 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_268 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_254 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_240 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_226 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_212 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_198 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_184 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_170 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_156 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_145 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_2_iw_p2_poisoned = _GEN_681 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_673 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_660 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_646 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_632 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_618 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_604 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_590 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_576 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_562 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_548 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_534 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_520 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_506 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_492 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_478 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_464 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_450 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_436 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_422 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_408 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_394 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_380 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_366 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_352 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_338 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_324 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_310 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_296 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_282 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_268 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_254 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_240 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_226 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_212 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_198 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_184 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_170 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_156 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_145 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_2_is_br = _GEN_681 ? _slots_39_io_uop_is_br : _GEN_673 ? _slots_38_io_uop_is_br : _GEN_660 ? _slots_37_io_uop_is_br : _GEN_646 ? _slots_36_io_uop_is_br : _GEN_632 ? _slots_35_io_uop_is_br : _GEN_618 ? _slots_34_io_uop_is_br : _GEN_604 ? _slots_33_io_uop_is_br : _GEN_590 ? _slots_32_io_uop_is_br : _GEN_576 ? _slots_31_io_uop_is_br : _GEN_562 ? _slots_30_io_uop_is_br : _GEN_548 ? _slots_29_io_uop_is_br : _GEN_534 ? _slots_28_io_uop_is_br : _GEN_520 ? _slots_27_io_uop_is_br : _GEN_506 ? _slots_26_io_uop_is_br : _GEN_492 ? _slots_25_io_uop_is_br : _GEN_478 ? _slots_24_io_uop_is_br : _GEN_464 ? _slots_23_io_uop_is_br : _GEN_450 ? _slots_22_io_uop_is_br : _GEN_436 ? _slots_21_io_uop_is_br : _GEN_422 ? _slots_20_io_uop_is_br : _GEN_408 ? _slots_19_io_uop_is_br : _GEN_394 ? _slots_18_io_uop_is_br : _GEN_380 ? _slots_17_io_uop_is_br : _GEN_366 ? _slots_16_io_uop_is_br : _GEN_352 ? _slots_15_io_uop_is_br : _GEN_338 ? _slots_14_io_uop_is_br : _GEN_324 ? _slots_13_io_uop_is_br : _GEN_310 ? _slots_12_io_uop_is_br : _GEN_296 ? _slots_11_io_uop_is_br : _GEN_282 ? _slots_10_io_uop_is_br : _GEN_268 ? _slots_9_io_uop_is_br : _GEN_254 ? _slots_8_io_uop_is_br : _GEN_240 ? _slots_7_io_uop_is_br : _GEN_226 ? _slots_6_io_uop_is_br : _GEN_212 ? _slots_5_io_uop_is_br : _GEN_198 ? _slots_4_io_uop_is_br : _GEN_184 ? _slots_3_io_uop_is_br : _GEN_170 ? _slots_2_io_uop_is_br : _GEN_156 ? _slots_1_io_uop_is_br : _GEN_145 & _slots_0_io_uop_is_br;
  assign io_iss_uops_2_is_jalr = _GEN_681 ? _slots_39_io_uop_is_jalr : _GEN_673 ? _slots_38_io_uop_is_jalr : _GEN_660 ? _slots_37_io_uop_is_jalr : _GEN_646 ? _slots_36_io_uop_is_jalr : _GEN_632 ? _slots_35_io_uop_is_jalr : _GEN_618 ? _slots_34_io_uop_is_jalr : _GEN_604 ? _slots_33_io_uop_is_jalr : _GEN_590 ? _slots_32_io_uop_is_jalr : _GEN_576 ? _slots_31_io_uop_is_jalr : _GEN_562 ? _slots_30_io_uop_is_jalr : _GEN_548 ? _slots_29_io_uop_is_jalr : _GEN_534 ? _slots_28_io_uop_is_jalr : _GEN_520 ? _slots_27_io_uop_is_jalr : _GEN_506 ? _slots_26_io_uop_is_jalr : _GEN_492 ? _slots_25_io_uop_is_jalr : _GEN_478 ? _slots_24_io_uop_is_jalr : _GEN_464 ? _slots_23_io_uop_is_jalr : _GEN_450 ? _slots_22_io_uop_is_jalr : _GEN_436 ? _slots_21_io_uop_is_jalr : _GEN_422 ? _slots_20_io_uop_is_jalr : _GEN_408 ? _slots_19_io_uop_is_jalr : _GEN_394 ? _slots_18_io_uop_is_jalr : _GEN_380 ? _slots_17_io_uop_is_jalr : _GEN_366 ? _slots_16_io_uop_is_jalr : _GEN_352 ? _slots_15_io_uop_is_jalr : _GEN_338 ? _slots_14_io_uop_is_jalr : _GEN_324 ? _slots_13_io_uop_is_jalr : _GEN_310 ? _slots_12_io_uop_is_jalr : _GEN_296 ? _slots_11_io_uop_is_jalr : _GEN_282 ? _slots_10_io_uop_is_jalr : _GEN_268 ? _slots_9_io_uop_is_jalr : _GEN_254 ? _slots_8_io_uop_is_jalr : _GEN_240 ? _slots_7_io_uop_is_jalr : _GEN_226 ? _slots_6_io_uop_is_jalr : _GEN_212 ? _slots_5_io_uop_is_jalr : _GEN_198 ? _slots_4_io_uop_is_jalr : _GEN_184 ? _slots_3_io_uop_is_jalr : _GEN_170 ? _slots_2_io_uop_is_jalr : _GEN_156 ? _slots_1_io_uop_is_jalr : _GEN_145 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_2_is_jal = _GEN_681 ? _slots_39_io_uop_is_jal : _GEN_673 ? _slots_38_io_uop_is_jal : _GEN_660 ? _slots_37_io_uop_is_jal : _GEN_646 ? _slots_36_io_uop_is_jal : _GEN_632 ? _slots_35_io_uop_is_jal : _GEN_618 ? _slots_34_io_uop_is_jal : _GEN_604 ? _slots_33_io_uop_is_jal : _GEN_590 ? _slots_32_io_uop_is_jal : _GEN_576 ? _slots_31_io_uop_is_jal : _GEN_562 ? _slots_30_io_uop_is_jal : _GEN_548 ? _slots_29_io_uop_is_jal : _GEN_534 ? _slots_28_io_uop_is_jal : _GEN_520 ? _slots_27_io_uop_is_jal : _GEN_506 ? _slots_26_io_uop_is_jal : _GEN_492 ? _slots_25_io_uop_is_jal : _GEN_478 ? _slots_24_io_uop_is_jal : _GEN_464 ? _slots_23_io_uop_is_jal : _GEN_450 ? _slots_22_io_uop_is_jal : _GEN_436 ? _slots_21_io_uop_is_jal : _GEN_422 ? _slots_20_io_uop_is_jal : _GEN_408 ? _slots_19_io_uop_is_jal : _GEN_394 ? _slots_18_io_uop_is_jal : _GEN_380 ? _slots_17_io_uop_is_jal : _GEN_366 ? _slots_16_io_uop_is_jal : _GEN_352 ? _slots_15_io_uop_is_jal : _GEN_338 ? _slots_14_io_uop_is_jal : _GEN_324 ? _slots_13_io_uop_is_jal : _GEN_310 ? _slots_12_io_uop_is_jal : _GEN_296 ? _slots_11_io_uop_is_jal : _GEN_282 ? _slots_10_io_uop_is_jal : _GEN_268 ? _slots_9_io_uop_is_jal : _GEN_254 ? _slots_8_io_uop_is_jal : _GEN_240 ? _slots_7_io_uop_is_jal : _GEN_226 ? _slots_6_io_uop_is_jal : _GEN_212 ? _slots_5_io_uop_is_jal : _GEN_198 ? _slots_4_io_uop_is_jal : _GEN_184 ? _slots_3_io_uop_is_jal : _GEN_170 ? _slots_2_io_uop_is_jal : _GEN_156 ? _slots_1_io_uop_is_jal : _GEN_145 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_2_is_sfb = _GEN_681 ? _slots_39_io_uop_is_sfb : _GEN_673 ? _slots_38_io_uop_is_sfb : _GEN_660 ? _slots_37_io_uop_is_sfb : _GEN_646 ? _slots_36_io_uop_is_sfb : _GEN_632 ? _slots_35_io_uop_is_sfb : _GEN_618 ? _slots_34_io_uop_is_sfb : _GEN_604 ? _slots_33_io_uop_is_sfb : _GEN_590 ? _slots_32_io_uop_is_sfb : _GEN_576 ? _slots_31_io_uop_is_sfb : _GEN_562 ? _slots_30_io_uop_is_sfb : _GEN_548 ? _slots_29_io_uop_is_sfb : _GEN_534 ? _slots_28_io_uop_is_sfb : _GEN_520 ? _slots_27_io_uop_is_sfb : _GEN_506 ? _slots_26_io_uop_is_sfb : _GEN_492 ? _slots_25_io_uop_is_sfb : _GEN_478 ? _slots_24_io_uop_is_sfb : _GEN_464 ? _slots_23_io_uop_is_sfb : _GEN_450 ? _slots_22_io_uop_is_sfb : _GEN_436 ? _slots_21_io_uop_is_sfb : _GEN_422 ? _slots_20_io_uop_is_sfb : _GEN_408 ? _slots_19_io_uop_is_sfb : _GEN_394 ? _slots_18_io_uop_is_sfb : _GEN_380 ? _slots_17_io_uop_is_sfb : _GEN_366 ? _slots_16_io_uop_is_sfb : _GEN_352 ? _slots_15_io_uop_is_sfb : _GEN_338 ? _slots_14_io_uop_is_sfb : _GEN_324 ? _slots_13_io_uop_is_sfb : _GEN_310 ? _slots_12_io_uop_is_sfb : _GEN_296 ? _slots_11_io_uop_is_sfb : _GEN_282 ? _slots_10_io_uop_is_sfb : _GEN_268 ? _slots_9_io_uop_is_sfb : _GEN_254 ? _slots_8_io_uop_is_sfb : _GEN_240 ? _slots_7_io_uop_is_sfb : _GEN_226 ? _slots_6_io_uop_is_sfb : _GEN_212 ? _slots_5_io_uop_is_sfb : _GEN_198 ? _slots_4_io_uop_is_sfb : _GEN_184 ? _slots_3_io_uop_is_sfb : _GEN_170 ? _slots_2_io_uop_is_sfb : _GEN_156 ? _slots_1_io_uop_is_sfb : _GEN_145 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_2_br_mask = _GEN_681 ? _slots_39_io_uop_br_mask : _GEN_673 ? _slots_38_io_uop_br_mask : _GEN_660 ? _slots_37_io_uop_br_mask : _GEN_646 ? _slots_36_io_uop_br_mask : _GEN_632 ? _slots_35_io_uop_br_mask : _GEN_618 ? _slots_34_io_uop_br_mask : _GEN_604 ? _slots_33_io_uop_br_mask : _GEN_590 ? _slots_32_io_uop_br_mask : _GEN_576 ? _slots_31_io_uop_br_mask : _GEN_562 ? _slots_30_io_uop_br_mask : _GEN_548 ? _slots_29_io_uop_br_mask : _GEN_534 ? _slots_28_io_uop_br_mask : _GEN_520 ? _slots_27_io_uop_br_mask : _GEN_506 ? _slots_26_io_uop_br_mask : _GEN_492 ? _slots_25_io_uop_br_mask : _GEN_478 ? _slots_24_io_uop_br_mask : _GEN_464 ? _slots_23_io_uop_br_mask : _GEN_450 ? _slots_22_io_uop_br_mask : _GEN_436 ? _slots_21_io_uop_br_mask : _GEN_422 ? _slots_20_io_uop_br_mask : _GEN_408 ? _slots_19_io_uop_br_mask : _GEN_394 ? _slots_18_io_uop_br_mask : _GEN_380 ? _slots_17_io_uop_br_mask : _GEN_366 ? _slots_16_io_uop_br_mask : _GEN_352 ? _slots_15_io_uop_br_mask : _GEN_338 ? _slots_14_io_uop_br_mask : _GEN_324 ? _slots_13_io_uop_br_mask : _GEN_310 ? _slots_12_io_uop_br_mask : _GEN_296 ? _slots_11_io_uop_br_mask : _GEN_282 ? _slots_10_io_uop_br_mask : _GEN_268 ? _slots_9_io_uop_br_mask : _GEN_254 ? _slots_8_io_uop_br_mask : _GEN_240 ? _slots_7_io_uop_br_mask : _GEN_226 ? _slots_6_io_uop_br_mask : _GEN_212 ? _slots_5_io_uop_br_mask : _GEN_198 ? _slots_4_io_uop_br_mask : _GEN_184 ? _slots_3_io_uop_br_mask : _GEN_170 ? _slots_2_io_uop_br_mask : _GEN_156 ? _slots_1_io_uop_br_mask : _GEN_145 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_2_br_tag = _GEN_681 ? _slots_39_io_uop_br_tag : _GEN_673 ? _slots_38_io_uop_br_tag : _GEN_660 ? _slots_37_io_uop_br_tag : _GEN_646 ? _slots_36_io_uop_br_tag : _GEN_632 ? _slots_35_io_uop_br_tag : _GEN_618 ? _slots_34_io_uop_br_tag : _GEN_604 ? _slots_33_io_uop_br_tag : _GEN_590 ? _slots_32_io_uop_br_tag : _GEN_576 ? _slots_31_io_uop_br_tag : _GEN_562 ? _slots_30_io_uop_br_tag : _GEN_548 ? _slots_29_io_uop_br_tag : _GEN_534 ? _slots_28_io_uop_br_tag : _GEN_520 ? _slots_27_io_uop_br_tag : _GEN_506 ? _slots_26_io_uop_br_tag : _GEN_492 ? _slots_25_io_uop_br_tag : _GEN_478 ? _slots_24_io_uop_br_tag : _GEN_464 ? _slots_23_io_uop_br_tag : _GEN_450 ? _slots_22_io_uop_br_tag : _GEN_436 ? _slots_21_io_uop_br_tag : _GEN_422 ? _slots_20_io_uop_br_tag : _GEN_408 ? _slots_19_io_uop_br_tag : _GEN_394 ? _slots_18_io_uop_br_tag : _GEN_380 ? _slots_17_io_uop_br_tag : _GEN_366 ? _slots_16_io_uop_br_tag : _GEN_352 ? _slots_15_io_uop_br_tag : _GEN_338 ? _slots_14_io_uop_br_tag : _GEN_324 ? _slots_13_io_uop_br_tag : _GEN_310 ? _slots_12_io_uop_br_tag : _GEN_296 ? _slots_11_io_uop_br_tag : _GEN_282 ? _slots_10_io_uop_br_tag : _GEN_268 ? _slots_9_io_uop_br_tag : _GEN_254 ? _slots_8_io_uop_br_tag : _GEN_240 ? _slots_7_io_uop_br_tag : _GEN_226 ? _slots_6_io_uop_br_tag : _GEN_212 ? _slots_5_io_uop_br_tag : _GEN_198 ? _slots_4_io_uop_br_tag : _GEN_184 ? _slots_3_io_uop_br_tag : _GEN_170 ? _slots_2_io_uop_br_tag : _GEN_156 ? _slots_1_io_uop_br_tag : _GEN_145 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_2_ftq_idx = _GEN_681 ? _slots_39_io_uop_ftq_idx : _GEN_673 ? _slots_38_io_uop_ftq_idx : _GEN_660 ? _slots_37_io_uop_ftq_idx : _GEN_646 ? _slots_36_io_uop_ftq_idx : _GEN_632 ? _slots_35_io_uop_ftq_idx : _GEN_618 ? _slots_34_io_uop_ftq_idx : _GEN_604 ? _slots_33_io_uop_ftq_idx : _GEN_590 ? _slots_32_io_uop_ftq_idx : _GEN_576 ? _slots_31_io_uop_ftq_idx : _GEN_562 ? _slots_30_io_uop_ftq_idx : _GEN_548 ? _slots_29_io_uop_ftq_idx : _GEN_534 ? _slots_28_io_uop_ftq_idx : _GEN_520 ? _slots_27_io_uop_ftq_idx : _GEN_506 ? _slots_26_io_uop_ftq_idx : _GEN_492 ? _slots_25_io_uop_ftq_idx : _GEN_478 ? _slots_24_io_uop_ftq_idx : _GEN_464 ? _slots_23_io_uop_ftq_idx : _GEN_450 ? _slots_22_io_uop_ftq_idx : _GEN_436 ? _slots_21_io_uop_ftq_idx : _GEN_422 ? _slots_20_io_uop_ftq_idx : _GEN_408 ? _slots_19_io_uop_ftq_idx : _GEN_394 ? _slots_18_io_uop_ftq_idx : _GEN_380 ? _slots_17_io_uop_ftq_idx : _GEN_366 ? _slots_16_io_uop_ftq_idx : _GEN_352 ? _slots_15_io_uop_ftq_idx : _GEN_338 ? _slots_14_io_uop_ftq_idx : _GEN_324 ? _slots_13_io_uop_ftq_idx : _GEN_310 ? _slots_12_io_uop_ftq_idx : _GEN_296 ? _slots_11_io_uop_ftq_idx : _GEN_282 ? _slots_10_io_uop_ftq_idx : _GEN_268 ? _slots_9_io_uop_ftq_idx : _GEN_254 ? _slots_8_io_uop_ftq_idx : _GEN_240 ? _slots_7_io_uop_ftq_idx : _GEN_226 ? _slots_6_io_uop_ftq_idx : _GEN_212 ? _slots_5_io_uop_ftq_idx : _GEN_198 ? _slots_4_io_uop_ftq_idx : _GEN_184 ? _slots_3_io_uop_ftq_idx : _GEN_170 ? _slots_2_io_uop_ftq_idx : _GEN_156 ? _slots_1_io_uop_ftq_idx : _GEN_145 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_2_edge_inst = _GEN_681 ? _slots_39_io_uop_edge_inst : _GEN_673 ? _slots_38_io_uop_edge_inst : _GEN_660 ? _slots_37_io_uop_edge_inst : _GEN_646 ? _slots_36_io_uop_edge_inst : _GEN_632 ? _slots_35_io_uop_edge_inst : _GEN_618 ? _slots_34_io_uop_edge_inst : _GEN_604 ? _slots_33_io_uop_edge_inst : _GEN_590 ? _slots_32_io_uop_edge_inst : _GEN_576 ? _slots_31_io_uop_edge_inst : _GEN_562 ? _slots_30_io_uop_edge_inst : _GEN_548 ? _slots_29_io_uop_edge_inst : _GEN_534 ? _slots_28_io_uop_edge_inst : _GEN_520 ? _slots_27_io_uop_edge_inst : _GEN_506 ? _slots_26_io_uop_edge_inst : _GEN_492 ? _slots_25_io_uop_edge_inst : _GEN_478 ? _slots_24_io_uop_edge_inst : _GEN_464 ? _slots_23_io_uop_edge_inst : _GEN_450 ? _slots_22_io_uop_edge_inst : _GEN_436 ? _slots_21_io_uop_edge_inst : _GEN_422 ? _slots_20_io_uop_edge_inst : _GEN_408 ? _slots_19_io_uop_edge_inst : _GEN_394 ? _slots_18_io_uop_edge_inst : _GEN_380 ? _slots_17_io_uop_edge_inst : _GEN_366 ? _slots_16_io_uop_edge_inst : _GEN_352 ? _slots_15_io_uop_edge_inst : _GEN_338 ? _slots_14_io_uop_edge_inst : _GEN_324 ? _slots_13_io_uop_edge_inst : _GEN_310 ? _slots_12_io_uop_edge_inst : _GEN_296 ? _slots_11_io_uop_edge_inst : _GEN_282 ? _slots_10_io_uop_edge_inst : _GEN_268 ? _slots_9_io_uop_edge_inst : _GEN_254 ? _slots_8_io_uop_edge_inst : _GEN_240 ? _slots_7_io_uop_edge_inst : _GEN_226 ? _slots_6_io_uop_edge_inst : _GEN_212 ? _slots_5_io_uop_edge_inst : _GEN_198 ? _slots_4_io_uop_edge_inst : _GEN_184 ? _slots_3_io_uop_edge_inst : _GEN_170 ? _slots_2_io_uop_edge_inst : _GEN_156 ? _slots_1_io_uop_edge_inst : _GEN_145 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_2_pc_lob = _GEN_681 ? _slots_39_io_uop_pc_lob : _GEN_673 ? _slots_38_io_uop_pc_lob : _GEN_660 ? _slots_37_io_uop_pc_lob : _GEN_646 ? _slots_36_io_uop_pc_lob : _GEN_632 ? _slots_35_io_uop_pc_lob : _GEN_618 ? _slots_34_io_uop_pc_lob : _GEN_604 ? _slots_33_io_uop_pc_lob : _GEN_590 ? _slots_32_io_uop_pc_lob : _GEN_576 ? _slots_31_io_uop_pc_lob : _GEN_562 ? _slots_30_io_uop_pc_lob : _GEN_548 ? _slots_29_io_uop_pc_lob : _GEN_534 ? _slots_28_io_uop_pc_lob : _GEN_520 ? _slots_27_io_uop_pc_lob : _GEN_506 ? _slots_26_io_uop_pc_lob : _GEN_492 ? _slots_25_io_uop_pc_lob : _GEN_478 ? _slots_24_io_uop_pc_lob : _GEN_464 ? _slots_23_io_uop_pc_lob : _GEN_450 ? _slots_22_io_uop_pc_lob : _GEN_436 ? _slots_21_io_uop_pc_lob : _GEN_422 ? _slots_20_io_uop_pc_lob : _GEN_408 ? _slots_19_io_uop_pc_lob : _GEN_394 ? _slots_18_io_uop_pc_lob : _GEN_380 ? _slots_17_io_uop_pc_lob : _GEN_366 ? _slots_16_io_uop_pc_lob : _GEN_352 ? _slots_15_io_uop_pc_lob : _GEN_338 ? _slots_14_io_uop_pc_lob : _GEN_324 ? _slots_13_io_uop_pc_lob : _GEN_310 ? _slots_12_io_uop_pc_lob : _GEN_296 ? _slots_11_io_uop_pc_lob : _GEN_282 ? _slots_10_io_uop_pc_lob : _GEN_268 ? _slots_9_io_uop_pc_lob : _GEN_254 ? _slots_8_io_uop_pc_lob : _GEN_240 ? _slots_7_io_uop_pc_lob : _GEN_226 ? _slots_6_io_uop_pc_lob : _GEN_212 ? _slots_5_io_uop_pc_lob : _GEN_198 ? _slots_4_io_uop_pc_lob : _GEN_184 ? _slots_3_io_uop_pc_lob : _GEN_170 ? _slots_2_io_uop_pc_lob : _GEN_156 ? _slots_1_io_uop_pc_lob : _GEN_145 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_2_taken = _GEN_681 ? _slots_39_io_uop_taken : _GEN_673 ? _slots_38_io_uop_taken : _GEN_660 ? _slots_37_io_uop_taken : _GEN_646 ? _slots_36_io_uop_taken : _GEN_632 ? _slots_35_io_uop_taken : _GEN_618 ? _slots_34_io_uop_taken : _GEN_604 ? _slots_33_io_uop_taken : _GEN_590 ? _slots_32_io_uop_taken : _GEN_576 ? _slots_31_io_uop_taken : _GEN_562 ? _slots_30_io_uop_taken : _GEN_548 ? _slots_29_io_uop_taken : _GEN_534 ? _slots_28_io_uop_taken : _GEN_520 ? _slots_27_io_uop_taken : _GEN_506 ? _slots_26_io_uop_taken : _GEN_492 ? _slots_25_io_uop_taken : _GEN_478 ? _slots_24_io_uop_taken : _GEN_464 ? _slots_23_io_uop_taken : _GEN_450 ? _slots_22_io_uop_taken : _GEN_436 ? _slots_21_io_uop_taken : _GEN_422 ? _slots_20_io_uop_taken : _GEN_408 ? _slots_19_io_uop_taken : _GEN_394 ? _slots_18_io_uop_taken : _GEN_380 ? _slots_17_io_uop_taken : _GEN_366 ? _slots_16_io_uop_taken : _GEN_352 ? _slots_15_io_uop_taken : _GEN_338 ? _slots_14_io_uop_taken : _GEN_324 ? _slots_13_io_uop_taken : _GEN_310 ? _slots_12_io_uop_taken : _GEN_296 ? _slots_11_io_uop_taken : _GEN_282 ? _slots_10_io_uop_taken : _GEN_268 ? _slots_9_io_uop_taken : _GEN_254 ? _slots_8_io_uop_taken : _GEN_240 ? _slots_7_io_uop_taken : _GEN_226 ? _slots_6_io_uop_taken : _GEN_212 ? _slots_5_io_uop_taken : _GEN_198 ? _slots_4_io_uop_taken : _GEN_184 ? _slots_3_io_uop_taken : _GEN_170 ? _slots_2_io_uop_taken : _GEN_156 ? _slots_1_io_uop_taken : _GEN_145 & _slots_0_io_uop_taken;
  assign io_iss_uops_2_imm_packed = _GEN_681 ? _slots_39_io_uop_imm_packed : _GEN_673 ? _slots_38_io_uop_imm_packed : _GEN_660 ? _slots_37_io_uop_imm_packed : _GEN_646 ? _slots_36_io_uop_imm_packed : _GEN_632 ? _slots_35_io_uop_imm_packed : _GEN_618 ? _slots_34_io_uop_imm_packed : _GEN_604 ? _slots_33_io_uop_imm_packed : _GEN_590 ? _slots_32_io_uop_imm_packed : _GEN_576 ? _slots_31_io_uop_imm_packed : _GEN_562 ? _slots_30_io_uop_imm_packed : _GEN_548 ? _slots_29_io_uop_imm_packed : _GEN_534 ? _slots_28_io_uop_imm_packed : _GEN_520 ? _slots_27_io_uop_imm_packed : _GEN_506 ? _slots_26_io_uop_imm_packed : _GEN_492 ? _slots_25_io_uop_imm_packed : _GEN_478 ? _slots_24_io_uop_imm_packed : _GEN_464 ? _slots_23_io_uop_imm_packed : _GEN_450 ? _slots_22_io_uop_imm_packed : _GEN_436 ? _slots_21_io_uop_imm_packed : _GEN_422 ? _slots_20_io_uop_imm_packed : _GEN_408 ? _slots_19_io_uop_imm_packed : _GEN_394 ? _slots_18_io_uop_imm_packed : _GEN_380 ? _slots_17_io_uop_imm_packed : _GEN_366 ? _slots_16_io_uop_imm_packed : _GEN_352 ? _slots_15_io_uop_imm_packed : _GEN_338 ? _slots_14_io_uop_imm_packed : _GEN_324 ? _slots_13_io_uop_imm_packed : _GEN_310 ? _slots_12_io_uop_imm_packed : _GEN_296 ? _slots_11_io_uop_imm_packed : _GEN_282 ? _slots_10_io_uop_imm_packed : _GEN_268 ? _slots_9_io_uop_imm_packed : _GEN_254 ? _slots_8_io_uop_imm_packed : _GEN_240 ? _slots_7_io_uop_imm_packed : _GEN_226 ? _slots_6_io_uop_imm_packed : _GEN_212 ? _slots_5_io_uop_imm_packed : _GEN_198 ? _slots_4_io_uop_imm_packed : _GEN_184 ? _slots_3_io_uop_imm_packed : _GEN_170 ? _slots_2_io_uop_imm_packed : _GEN_156 ? _slots_1_io_uop_imm_packed : _GEN_145 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_2_rob_idx = _GEN_681 ? _slots_39_io_uop_rob_idx : _GEN_673 ? _slots_38_io_uop_rob_idx : _GEN_660 ? _slots_37_io_uop_rob_idx : _GEN_646 ? _slots_36_io_uop_rob_idx : _GEN_632 ? _slots_35_io_uop_rob_idx : _GEN_618 ? _slots_34_io_uop_rob_idx : _GEN_604 ? _slots_33_io_uop_rob_idx : _GEN_590 ? _slots_32_io_uop_rob_idx : _GEN_576 ? _slots_31_io_uop_rob_idx : _GEN_562 ? _slots_30_io_uop_rob_idx : _GEN_548 ? _slots_29_io_uop_rob_idx : _GEN_534 ? _slots_28_io_uop_rob_idx : _GEN_520 ? _slots_27_io_uop_rob_idx : _GEN_506 ? _slots_26_io_uop_rob_idx : _GEN_492 ? _slots_25_io_uop_rob_idx : _GEN_478 ? _slots_24_io_uop_rob_idx : _GEN_464 ? _slots_23_io_uop_rob_idx : _GEN_450 ? _slots_22_io_uop_rob_idx : _GEN_436 ? _slots_21_io_uop_rob_idx : _GEN_422 ? _slots_20_io_uop_rob_idx : _GEN_408 ? _slots_19_io_uop_rob_idx : _GEN_394 ? _slots_18_io_uop_rob_idx : _GEN_380 ? _slots_17_io_uop_rob_idx : _GEN_366 ? _slots_16_io_uop_rob_idx : _GEN_352 ? _slots_15_io_uop_rob_idx : _GEN_338 ? _slots_14_io_uop_rob_idx : _GEN_324 ? _slots_13_io_uop_rob_idx : _GEN_310 ? _slots_12_io_uop_rob_idx : _GEN_296 ? _slots_11_io_uop_rob_idx : _GEN_282 ? _slots_10_io_uop_rob_idx : _GEN_268 ? _slots_9_io_uop_rob_idx : _GEN_254 ? _slots_8_io_uop_rob_idx : _GEN_240 ? _slots_7_io_uop_rob_idx : _GEN_226 ? _slots_6_io_uop_rob_idx : _GEN_212 ? _slots_5_io_uop_rob_idx : _GEN_198 ? _slots_4_io_uop_rob_idx : _GEN_184 ? _slots_3_io_uop_rob_idx : _GEN_170 ? _slots_2_io_uop_rob_idx : _GEN_156 ? _slots_1_io_uop_rob_idx : _GEN_145 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_2_ldq_idx = _GEN_681 ? _slots_39_io_uop_ldq_idx : _GEN_673 ? _slots_38_io_uop_ldq_idx : _GEN_660 ? _slots_37_io_uop_ldq_idx : _GEN_646 ? _slots_36_io_uop_ldq_idx : _GEN_632 ? _slots_35_io_uop_ldq_idx : _GEN_618 ? _slots_34_io_uop_ldq_idx : _GEN_604 ? _slots_33_io_uop_ldq_idx : _GEN_590 ? _slots_32_io_uop_ldq_idx : _GEN_576 ? _slots_31_io_uop_ldq_idx : _GEN_562 ? _slots_30_io_uop_ldq_idx : _GEN_548 ? _slots_29_io_uop_ldq_idx : _GEN_534 ? _slots_28_io_uop_ldq_idx : _GEN_520 ? _slots_27_io_uop_ldq_idx : _GEN_506 ? _slots_26_io_uop_ldq_idx : _GEN_492 ? _slots_25_io_uop_ldq_idx : _GEN_478 ? _slots_24_io_uop_ldq_idx : _GEN_464 ? _slots_23_io_uop_ldq_idx : _GEN_450 ? _slots_22_io_uop_ldq_idx : _GEN_436 ? _slots_21_io_uop_ldq_idx : _GEN_422 ? _slots_20_io_uop_ldq_idx : _GEN_408 ? _slots_19_io_uop_ldq_idx : _GEN_394 ? _slots_18_io_uop_ldq_idx : _GEN_380 ? _slots_17_io_uop_ldq_idx : _GEN_366 ? _slots_16_io_uop_ldq_idx : _GEN_352 ? _slots_15_io_uop_ldq_idx : _GEN_338 ? _slots_14_io_uop_ldq_idx : _GEN_324 ? _slots_13_io_uop_ldq_idx : _GEN_310 ? _slots_12_io_uop_ldq_idx : _GEN_296 ? _slots_11_io_uop_ldq_idx : _GEN_282 ? _slots_10_io_uop_ldq_idx : _GEN_268 ? _slots_9_io_uop_ldq_idx : _GEN_254 ? _slots_8_io_uop_ldq_idx : _GEN_240 ? _slots_7_io_uop_ldq_idx : _GEN_226 ? _slots_6_io_uop_ldq_idx : _GEN_212 ? _slots_5_io_uop_ldq_idx : _GEN_198 ? _slots_4_io_uop_ldq_idx : _GEN_184 ? _slots_3_io_uop_ldq_idx : _GEN_170 ? _slots_2_io_uop_ldq_idx : _GEN_156 ? _slots_1_io_uop_ldq_idx : _GEN_145 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_2_stq_idx = _GEN_681 ? _slots_39_io_uop_stq_idx : _GEN_673 ? _slots_38_io_uop_stq_idx : _GEN_660 ? _slots_37_io_uop_stq_idx : _GEN_646 ? _slots_36_io_uop_stq_idx : _GEN_632 ? _slots_35_io_uop_stq_idx : _GEN_618 ? _slots_34_io_uop_stq_idx : _GEN_604 ? _slots_33_io_uop_stq_idx : _GEN_590 ? _slots_32_io_uop_stq_idx : _GEN_576 ? _slots_31_io_uop_stq_idx : _GEN_562 ? _slots_30_io_uop_stq_idx : _GEN_548 ? _slots_29_io_uop_stq_idx : _GEN_534 ? _slots_28_io_uop_stq_idx : _GEN_520 ? _slots_27_io_uop_stq_idx : _GEN_506 ? _slots_26_io_uop_stq_idx : _GEN_492 ? _slots_25_io_uop_stq_idx : _GEN_478 ? _slots_24_io_uop_stq_idx : _GEN_464 ? _slots_23_io_uop_stq_idx : _GEN_450 ? _slots_22_io_uop_stq_idx : _GEN_436 ? _slots_21_io_uop_stq_idx : _GEN_422 ? _slots_20_io_uop_stq_idx : _GEN_408 ? _slots_19_io_uop_stq_idx : _GEN_394 ? _slots_18_io_uop_stq_idx : _GEN_380 ? _slots_17_io_uop_stq_idx : _GEN_366 ? _slots_16_io_uop_stq_idx : _GEN_352 ? _slots_15_io_uop_stq_idx : _GEN_338 ? _slots_14_io_uop_stq_idx : _GEN_324 ? _slots_13_io_uop_stq_idx : _GEN_310 ? _slots_12_io_uop_stq_idx : _GEN_296 ? _slots_11_io_uop_stq_idx : _GEN_282 ? _slots_10_io_uop_stq_idx : _GEN_268 ? _slots_9_io_uop_stq_idx : _GEN_254 ? _slots_8_io_uop_stq_idx : _GEN_240 ? _slots_7_io_uop_stq_idx : _GEN_226 ? _slots_6_io_uop_stq_idx : _GEN_212 ? _slots_5_io_uop_stq_idx : _GEN_198 ? _slots_4_io_uop_stq_idx : _GEN_184 ? _slots_3_io_uop_stq_idx : _GEN_170 ? _slots_2_io_uop_stq_idx : _GEN_156 ? _slots_1_io_uop_stq_idx : _GEN_145 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_2_pdst = _GEN_681 ? _slots_39_io_uop_pdst : _GEN_673 ? _slots_38_io_uop_pdst : _GEN_660 ? _slots_37_io_uop_pdst : _GEN_646 ? _slots_36_io_uop_pdst : _GEN_632 ? _slots_35_io_uop_pdst : _GEN_618 ? _slots_34_io_uop_pdst : _GEN_604 ? _slots_33_io_uop_pdst : _GEN_590 ? _slots_32_io_uop_pdst : _GEN_576 ? _slots_31_io_uop_pdst : _GEN_562 ? _slots_30_io_uop_pdst : _GEN_548 ? _slots_29_io_uop_pdst : _GEN_534 ? _slots_28_io_uop_pdst : _GEN_520 ? _slots_27_io_uop_pdst : _GEN_506 ? _slots_26_io_uop_pdst : _GEN_492 ? _slots_25_io_uop_pdst : _GEN_478 ? _slots_24_io_uop_pdst : _GEN_464 ? _slots_23_io_uop_pdst : _GEN_450 ? _slots_22_io_uop_pdst : _GEN_436 ? _slots_21_io_uop_pdst : _GEN_422 ? _slots_20_io_uop_pdst : _GEN_408 ? _slots_19_io_uop_pdst : _GEN_394 ? _slots_18_io_uop_pdst : _GEN_380 ? _slots_17_io_uop_pdst : _GEN_366 ? _slots_16_io_uop_pdst : _GEN_352 ? _slots_15_io_uop_pdst : _GEN_338 ? _slots_14_io_uop_pdst : _GEN_324 ? _slots_13_io_uop_pdst : _GEN_310 ? _slots_12_io_uop_pdst : _GEN_296 ? _slots_11_io_uop_pdst : _GEN_282 ? _slots_10_io_uop_pdst : _GEN_268 ? _slots_9_io_uop_pdst : _GEN_254 ? _slots_8_io_uop_pdst : _GEN_240 ? _slots_7_io_uop_pdst : _GEN_226 ? _slots_6_io_uop_pdst : _GEN_212 ? _slots_5_io_uop_pdst : _GEN_198 ? _slots_4_io_uop_pdst : _GEN_184 ? _slots_3_io_uop_pdst : _GEN_170 ? _slots_2_io_uop_pdst : _GEN_156 ? _slots_1_io_uop_pdst : _GEN_145 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_2_prs1 = _GEN_681 ? _slots_39_io_uop_prs1 : _GEN_673 ? _slots_38_io_uop_prs1 : _GEN_660 ? _slots_37_io_uop_prs1 : _GEN_646 ? _slots_36_io_uop_prs1 : _GEN_632 ? _slots_35_io_uop_prs1 : _GEN_618 ? _slots_34_io_uop_prs1 : _GEN_604 ? _slots_33_io_uop_prs1 : _GEN_590 ? _slots_32_io_uop_prs1 : _GEN_576 ? _slots_31_io_uop_prs1 : _GEN_562 ? _slots_30_io_uop_prs1 : _GEN_548 ? _slots_29_io_uop_prs1 : _GEN_534 ? _slots_28_io_uop_prs1 : _GEN_520 ? _slots_27_io_uop_prs1 : _GEN_506 ? _slots_26_io_uop_prs1 : _GEN_492 ? _slots_25_io_uop_prs1 : _GEN_478 ? _slots_24_io_uop_prs1 : _GEN_464 ? _slots_23_io_uop_prs1 : _GEN_450 ? _slots_22_io_uop_prs1 : _GEN_436 ? _slots_21_io_uop_prs1 : _GEN_422 ? _slots_20_io_uop_prs1 : _GEN_408 ? _slots_19_io_uop_prs1 : _GEN_394 ? _slots_18_io_uop_prs1 : _GEN_380 ? _slots_17_io_uop_prs1 : _GEN_366 ? _slots_16_io_uop_prs1 : _GEN_352 ? _slots_15_io_uop_prs1 : _GEN_338 ? _slots_14_io_uop_prs1 : _GEN_324 ? _slots_13_io_uop_prs1 : _GEN_310 ? _slots_12_io_uop_prs1 : _GEN_296 ? _slots_11_io_uop_prs1 : _GEN_282 ? _slots_10_io_uop_prs1 : _GEN_268 ? _slots_9_io_uop_prs1 : _GEN_254 ? _slots_8_io_uop_prs1 : _GEN_240 ? _slots_7_io_uop_prs1 : _GEN_226 ? _slots_6_io_uop_prs1 : _GEN_212 ? _slots_5_io_uop_prs1 : _GEN_198 ? _slots_4_io_uop_prs1 : _GEN_184 ? _slots_3_io_uop_prs1 : _GEN_170 ? _slots_2_io_uop_prs1 : _GEN_156 ? _slots_1_io_uop_prs1 : _GEN_145 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_2_prs2 = _GEN_681 ? _slots_39_io_uop_prs2 : _GEN_673 ? _slots_38_io_uop_prs2 : _GEN_660 ? _slots_37_io_uop_prs2 : _GEN_646 ? _slots_36_io_uop_prs2 : _GEN_632 ? _slots_35_io_uop_prs2 : _GEN_618 ? _slots_34_io_uop_prs2 : _GEN_604 ? _slots_33_io_uop_prs2 : _GEN_590 ? _slots_32_io_uop_prs2 : _GEN_576 ? _slots_31_io_uop_prs2 : _GEN_562 ? _slots_30_io_uop_prs2 : _GEN_548 ? _slots_29_io_uop_prs2 : _GEN_534 ? _slots_28_io_uop_prs2 : _GEN_520 ? _slots_27_io_uop_prs2 : _GEN_506 ? _slots_26_io_uop_prs2 : _GEN_492 ? _slots_25_io_uop_prs2 : _GEN_478 ? _slots_24_io_uop_prs2 : _GEN_464 ? _slots_23_io_uop_prs2 : _GEN_450 ? _slots_22_io_uop_prs2 : _GEN_436 ? _slots_21_io_uop_prs2 : _GEN_422 ? _slots_20_io_uop_prs2 : _GEN_408 ? _slots_19_io_uop_prs2 : _GEN_394 ? _slots_18_io_uop_prs2 : _GEN_380 ? _slots_17_io_uop_prs2 : _GEN_366 ? _slots_16_io_uop_prs2 : _GEN_352 ? _slots_15_io_uop_prs2 : _GEN_338 ? _slots_14_io_uop_prs2 : _GEN_324 ? _slots_13_io_uop_prs2 : _GEN_310 ? _slots_12_io_uop_prs2 : _GEN_296 ? _slots_11_io_uop_prs2 : _GEN_282 ? _slots_10_io_uop_prs2 : _GEN_268 ? _slots_9_io_uop_prs2 : _GEN_254 ? _slots_8_io_uop_prs2 : _GEN_240 ? _slots_7_io_uop_prs2 : _GEN_226 ? _slots_6_io_uop_prs2 : _GEN_212 ? _slots_5_io_uop_prs2 : _GEN_198 ? _slots_4_io_uop_prs2 : _GEN_184 ? _slots_3_io_uop_prs2 : _GEN_170 ? _slots_2_io_uop_prs2 : _GEN_156 ? _slots_1_io_uop_prs2 : _GEN_145 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_2_bypassable = _GEN_681 ? _slots_39_io_uop_bypassable : _GEN_673 ? _slots_38_io_uop_bypassable : _GEN_660 ? _slots_37_io_uop_bypassable : _GEN_646 ? _slots_36_io_uop_bypassable : _GEN_632 ? _slots_35_io_uop_bypassable : _GEN_618 ? _slots_34_io_uop_bypassable : _GEN_604 ? _slots_33_io_uop_bypassable : _GEN_590 ? _slots_32_io_uop_bypassable : _GEN_576 ? _slots_31_io_uop_bypassable : _GEN_562 ? _slots_30_io_uop_bypassable : _GEN_548 ? _slots_29_io_uop_bypassable : _GEN_534 ? _slots_28_io_uop_bypassable : _GEN_520 ? _slots_27_io_uop_bypassable : _GEN_506 ? _slots_26_io_uop_bypassable : _GEN_492 ? _slots_25_io_uop_bypassable : _GEN_478 ? _slots_24_io_uop_bypassable : _GEN_464 ? _slots_23_io_uop_bypassable : _GEN_450 ? _slots_22_io_uop_bypassable : _GEN_436 ? _slots_21_io_uop_bypassable : _GEN_422 ? _slots_20_io_uop_bypassable : _GEN_408 ? _slots_19_io_uop_bypassable : _GEN_394 ? _slots_18_io_uop_bypassable : _GEN_380 ? _slots_17_io_uop_bypassable : _GEN_366 ? _slots_16_io_uop_bypassable : _GEN_352 ? _slots_15_io_uop_bypassable : _GEN_338 ? _slots_14_io_uop_bypassable : _GEN_324 ? _slots_13_io_uop_bypassable : _GEN_310 ? _slots_12_io_uop_bypassable : _GEN_296 ? _slots_11_io_uop_bypassable : _GEN_282 ? _slots_10_io_uop_bypassable : _GEN_268 ? _slots_9_io_uop_bypassable : _GEN_254 ? _slots_8_io_uop_bypassable : _GEN_240 ? _slots_7_io_uop_bypassable : _GEN_226 ? _slots_6_io_uop_bypassable : _GEN_212 ? _slots_5_io_uop_bypassable : _GEN_198 ? _slots_4_io_uop_bypassable : _GEN_184 ? _slots_3_io_uop_bypassable : _GEN_170 ? _slots_2_io_uop_bypassable : _GEN_156 ? _slots_1_io_uop_bypassable : _GEN_145 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_2_mem_cmd = _GEN_681 ? _slots_39_io_uop_mem_cmd : _GEN_673 ? _slots_38_io_uop_mem_cmd : _GEN_660 ? _slots_37_io_uop_mem_cmd : _GEN_646 ? _slots_36_io_uop_mem_cmd : _GEN_632 ? _slots_35_io_uop_mem_cmd : _GEN_618 ? _slots_34_io_uop_mem_cmd : _GEN_604 ? _slots_33_io_uop_mem_cmd : _GEN_590 ? _slots_32_io_uop_mem_cmd : _GEN_576 ? _slots_31_io_uop_mem_cmd : _GEN_562 ? _slots_30_io_uop_mem_cmd : _GEN_548 ? _slots_29_io_uop_mem_cmd : _GEN_534 ? _slots_28_io_uop_mem_cmd : _GEN_520 ? _slots_27_io_uop_mem_cmd : _GEN_506 ? _slots_26_io_uop_mem_cmd : _GEN_492 ? _slots_25_io_uop_mem_cmd : _GEN_478 ? _slots_24_io_uop_mem_cmd : _GEN_464 ? _slots_23_io_uop_mem_cmd : _GEN_450 ? _slots_22_io_uop_mem_cmd : _GEN_436 ? _slots_21_io_uop_mem_cmd : _GEN_422 ? _slots_20_io_uop_mem_cmd : _GEN_408 ? _slots_19_io_uop_mem_cmd : _GEN_394 ? _slots_18_io_uop_mem_cmd : _GEN_380 ? _slots_17_io_uop_mem_cmd : _GEN_366 ? _slots_16_io_uop_mem_cmd : _GEN_352 ? _slots_15_io_uop_mem_cmd : _GEN_338 ? _slots_14_io_uop_mem_cmd : _GEN_324 ? _slots_13_io_uop_mem_cmd : _GEN_310 ? _slots_12_io_uop_mem_cmd : _GEN_296 ? _slots_11_io_uop_mem_cmd : _GEN_282 ? _slots_10_io_uop_mem_cmd : _GEN_268 ? _slots_9_io_uop_mem_cmd : _GEN_254 ? _slots_8_io_uop_mem_cmd : _GEN_240 ? _slots_7_io_uop_mem_cmd : _GEN_226 ? _slots_6_io_uop_mem_cmd : _GEN_212 ? _slots_5_io_uop_mem_cmd : _GEN_198 ? _slots_4_io_uop_mem_cmd : _GEN_184 ? _slots_3_io_uop_mem_cmd : _GEN_170 ? _slots_2_io_uop_mem_cmd : _GEN_156 ? _slots_1_io_uop_mem_cmd : _GEN_145 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_2_is_amo = _GEN_681 ? _slots_39_io_uop_is_amo : _GEN_673 ? _slots_38_io_uop_is_amo : _GEN_660 ? _slots_37_io_uop_is_amo : _GEN_646 ? _slots_36_io_uop_is_amo : _GEN_632 ? _slots_35_io_uop_is_amo : _GEN_618 ? _slots_34_io_uop_is_amo : _GEN_604 ? _slots_33_io_uop_is_amo : _GEN_590 ? _slots_32_io_uop_is_amo : _GEN_576 ? _slots_31_io_uop_is_amo : _GEN_562 ? _slots_30_io_uop_is_amo : _GEN_548 ? _slots_29_io_uop_is_amo : _GEN_534 ? _slots_28_io_uop_is_amo : _GEN_520 ? _slots_27_io_uop_is_amo : _GEN_506 ? _slots_26_io_uop_is_amo : _GEN_492 ? _slots_25_io_uop_is_amo : _GEN_478 ? _slots_24_io_uop_is_amo : _GEN_464 ? _slots_23_io_uop_is_amo : _GEN_450 ? _slots_22_io_uop_is_amo : _GEN_436 ? _slots_21_io_uop_is_amo : _GEN_422 ? _slots_20_io_uop_is_amo : _GEN_408 ? _slots_19_io_uop_is_amo : _GEN_394 ? _slots_18_io_uop_is_amo : _GEN_380 ? _slots_17_io_uop_is_amo : _GEN_366 ? _slots_16_io_uop_is_amo : _GEN_352 ? _slots_15_io_uop_is_amo : _GEN_338 ? _slots_14_io_uop_is_amo : _GEN_324 ? _slots_13_io_uop_is_amo : _GEN_310 ? _slots_12_io_uop_is_amo : _GEN_296 ? _slots_11_io_uop_is_amo : _GEN_282 ? _slots_10_io_uop_is_amo : _GEN_268 ? _slots_9_io_uop_is_amo : _GEN_254 ? _slots_8_io_uop_is_amo : _GEN_240 ? _slots_7_io_uop_is_amo : _GEN_226 ? _slots_6_io_uop_is_amo : _GEN_212 ? _slots_5_io_uop_is_amo : _GEN_198 ? _slots_4_io_uop_is_amo : _GEN_184 ? _slots_3_io_uop_is_amo : _GEN_170 ? _slots_2_io_uop_is_amo : _GEN_156 ? _slots_1_io_uop_is_amo : _GEN_145 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_2_uses_stq = _GEN_681 ? _slots_39_io_uop_uses_stq : _GEN_673 ? _slots_38_io_uop_uses_stq : _GEN_660 ? _slots_37_io_uop_uses_stq : _GEN_646 ? _slots_36_io_uop_uses_stq : _GEN_632 ? _slots_35_io_uop_uses_stq : _GEN_618 ? _slots_34_io_uop_uses_stq : _GEN_604 ? _slots_33_io_uop_uses_stq : _GEN_590 ? _slots_32_io_uop_uses_stq : _GEN_576 ? _slots_31_io_uop_uses_stq : _GEN_562 ? _slots_30_io_uop_uses_stq : _GEN_548 ? _slots_29_io_uop_uses_stq : _GEN_534 ? _slots_28_io_uop_uses_stq : _GEN_520 ? _slots_27_io_uop_uses_stq : _GEN_506 ? _slots_26_io_uop_uses_stq : _GEN_492 ? _slots_25_io_uop_uses_stq : _GEN_478 ? _slots_24_io_uop_uses_stq : _GEN_464 ? _slots_23_io_uop_uses_stq : _GEN_450 ? _slots_22_io_uop_uses_stq : _GEN_436 ? _slots_21_io_uop_uses_stq : _GEN_422 ? _slots_20_io_uop_uses_stq : _GEN_408 ? _slots_19_io_uop_uses_stq : _GEN_394 ? _slots_18_io_uop_uses_stq : _GEN_380 ? _slots_17_io_uop_uses_stq : _GEN_366 ? _slots_16_io_uop_uses_stq : _GEN_352 ? _slots_15_io_uop_uses_stq : _GEN_338 ? _slots_14_io_uop_uses_stq : _GEN_324 ? _slots_13_io_uop_uses_stq : _GEN_310 ? _slots_12_io_uop_uses_stq : _GEN_296 ? _slots_11_io_uop_uses_stq : _GEN_282 ? _slots_10_io_uop_uses_stq : _GEN_268 ? _slots_9_io_uop_uses_stq : _GEN_254 ? _slots_8_io_uop_uses_stq : _GEN_240 ? _slots_7_io_uop_uses_stq : _GEN_226 ? _slots_6_io_uop_uses_stq : _GEN_212 ? _slots_5_io_uop_uses_stq : _GEN_198 ? _slots_4_io_uop_uses_stq : _GEN_184 ? _slots_3_io_uop_uses_stq : _GEN_170 ? _slots_2_io_uop_uses_stq : _GEN_156 ? _slots_1_io_uop_uses_stq : _GEN_145 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_2_ldst_val = _GEN_681 ? _slots_39_io_uop_ldst_val : _GEN_673 ? _slots_38_io_uop_ldst_val : _GEN_660 ? _slots_37_io_uop_ldst_val : _GEN_646 ? _slots_36_io_uop_ldst_val : _GEN_632 ? _slots_35_io_uop_ldst_val : _GEN_618 ? _slots_34_io_uop_ldst_val : _GEN_604 ? _slots_33_io_uop_ldst_val : _GEN_590 ? _slots_32_io_uop_ldst_val : _GEN_576 ? _slots_31_io_uop_ldst_val : _GEN_562 ? _slots_30_io_uop_ldst_val : _GEN_548 ? _slots_29_io_uop_ldst_val : _GEN_534 ? _slots_28_io_uop_ldst_val : _GEN_520 ? _slots_27_io_uop_ldst_val : _GEN_506 ? _slots_26_io_uop_ldst_val : _GEN_492 ? _slots_25_io_uop_ldst_val : _GEN_478 ? _slots_24_io_uop_ldst_val : _GEN_464 ? _slots_23_io_uop_ldst_val : _GEN_450 ? _slots_22_io_uop_ldst_val : _GEN_436 ? _slots_21_io_uop_ldst_val : _GEN_422 ? _slots_20_io_uop_ldst_val : _GEN_408 ? _slots_19_io_uop_ldst_val : _GEN_394 ? _slots_18_io_uop_ldst_val : _GEN_380 ? _slots_17_io_uop_ldst_val : _GEN_366 ? _slots_16_io_uop_ldst_val : _GEN_352 ? _slots_15_io_uop_ldst_val : _GEN_338 ? _slots_14_io_uop_ldst_val : _GEN_324 ? _slots_13_io_uop_ldst_val : _GEN_310 ? _slots_12_io_uop_ldst_val : _GEN_296 ? _slots_11_io_uop_ldst_val : _GEN_282 ? _slots_10_io_uop_ldst_val : _GEN_268 ? _slots_9_io_uop_ldst_val : _GEN_254 ? _slots_8_io_uop_ldst_val : _GEN_240 ? _slots_7_io_uop_ldst_val : _GEN_226 ? _slots_6_io_uop_ldst_val : _GEN_212 ? _slots_5_io_uop_ldst_val : _GEN_198 ? _slots_4_io_uop_ldst_val : _GEN_184 ? _slots_3_io_uop_ldst_val : _GEN_170 ? _slots_2_io_uop_ldst_val : _GEN_156 ? _slots_1_io_uop_ldst_val : _GEN_145 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_2_dst_rtype = _GEN_681 ? _slots_39_io_uop_dst_rtype : _GEN_673 ? _slots_38_io_uop_dst_rtype : _GEN_660 ? _slots_37_io_uop_dst_rtype : _GEN_646 ? _slots_36_io_uop_dst_rtype : _GEN_632 ? _slots_35_io_uop_dst_rtype : _GEN_618 ? _slots_34_io_uop_dst_rtype : _GEN_604 ? _slots_33_io_uop_dst_rtype : _GEN_590 ? _slots_32_io_uop_dst_rtype : _GEN_576 ? _slots_31_io_uop_dst_rtype : _GEN_562 ? _slots_30_io_uop_dst_rtype : _GEN_548 ? _slots_29_io_uop_dst_rtype : _GEN_534 ? _slots_28_io_uop_dst_rtype : _GEN_520 ? _slots_27_io_uop_dst_rtype : _GEN_506 ? _slots_26_io_uop_dst_rtype : _GEN_492 ? _slots_25_io_uop_dst_rtype : _GEN_478 ? _slots_24_io_uop_dst_rtype : _GEN_464 ? _slots_23_io_uop_dst_rtype : _GEN_450 ? _slots_22_io_uop_dst_rtype : _GEN_436 ? _slots_21_io_uop_dst_rtype : _GEN_422 ? _slots_20_io_uop_dst_rtype : _GEN_408 ? _slots_19_io_uop_dst_rtype : _GEN_394 ? _slots_18_io_uop_dst_rtype : _GEN_380 ? _slots_17_io_uop_dst_rtype : _GEN_366 ? _slots_16_io_uop_dst_rtype : _GEN_352 ? _slots_15_io_uop_dst_rtype : _GEN_338 ? _slots_14_io_uop_dst_rtype : _GEN_324 ? _slots_13_io_uop_dst_rtype : _GEN_310 ? _slots_12_io_uop_dst_rtype : _GEN_296 ? _slots_11_io_uop_dst_rtype : _GEN_282 ? _slots_10_io_uop_dst_rtype : _GEN_268 ? _slots_9_io_uop_dst_rtype : _GEN_254 ? _slots_8_io_uop_dst_rtype : _GEN_240 ? _slots_7_io_uop_dst_rtype : _GEN_226 ? _slots_6_io_uop_dst_rtype : _GEN_212 ? _slots_5_io_uop_dst_rtype : _GEN_198 ? _slots_4_io_uop_dst_rtype : _GEN_184 ? _slots_3_io_uop_dst_rtype : _GEN_170 ? _slots_2_io_uop_dst_rtype : _GEN_156 ? _slots_1_io_uop_dst_rtype : _GEN_145 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_2_lrs1_rtype = _GEN_681 ? _slots_39_io_uop_lrs1_rtype : _GEN_673 ? _slots_38_io_uop_lrs1_rtype : _GEN_660 ? _slots_37_io_uop_lrs1_rtype : _GEN_646 ? _slots_36_io_uop_lrs1_rtype : _GEN_632 ? _slots_35_io_uop_lrs1_rtype : _GEN_618 ? _slots_34_io_uop_lrs1_rtype : _GEN_604 ? _slots_33_io_uop_lrs1_rtype : _GEN_590 ? _slots_32_io_uop_lrs1_rtype : _GEN_576 ? _slots_31_io_uop_lrs1_rtype : _GEN_562 ? _slots_30_io_uop_lrs1_rtype : _GEN_548 ? _slots_29_io_uop_lrs1_rtype : _GEN_534 ? _slots_28_io_uop_lrs1_rtype : _GEN_520 ? _slots_27_io_uop_lrs1_rtype : _GEN_506 ? _slots_26_io_uop_lrs1_rtype : _GEN_492 ? _slots_25_io_uop_lrs1_rtype : _GEN_478 ? _slots_24_io_uop_lrs1_rtype : _GEN_464 ? _slots_23_io_uop_lrs1_rtype : _GEN_450 ? _slots_22_io_uop_lrs1_rtype : _GEN_436 ? _slots_21_io_uop_lrs1_rtype : _GEN_422 ? _slots_20_io_uop_lrs1_rtype : _GEN_408 ? _slots_19_io_uop_lrs1_rtype : _GEN_394 ? _slots_18_io_uop_lrs1_rtype : _GEN_380 ? _slots_17_io_uop_lrs1_rtype : _GEN_366 ? _slots_16_io_uop_lrs1_rtype : _GEN_352 ? _slots_15_io_uop_lrs1_rtype : _GEN_338 ? _slots_14_io_uop_lrs1_rtype : _GEN_324 ? _slots_13_io_uop_lrs1_rtype : _GEN_310 ? _slots_12_io_uop_lrs1_rtype : _GEN_296 ? _slots_11_io_uop_lrs1_rtype : _GEN_282 ? _slots_10_io_uop_lrs1_rtype : _GEN_268 ? _slots_9_io_uop_lrs1_rtype : _GEN_254 ? _slots_8_io_uop_lrs1_rtype : _GEN_240 ? _slots_7_io_uop_lrs1_rtype : _GEN_226 ? _slots_6_io_uop_lrs1_rtype : _GEN_212 ? _slots_5_io_uop_lrs1_rtype : _GEN_198 ? _slots_4_io_uop_lrs1_rtype : _GEN_184 ? _slots_3_io_uop_lrs1_rtype : _GEN_170 ? _slots_2_io_uop_lrs1_rtype : _GEN_156 ? _slots_1_io_uop_lrs1_rtype : _GEN_145 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_2_lrs2_rtype = _GEN_681 ? _slots_39_io_uop_lrs2_rtype : _GEN_673 ? _slots_38_io_uop_lrs2_rtype : _GEN_660 ? _slots_37_io_uop_lrs2_rtype : _GEN_646 ? _slots_36_io_uop_lrs2_rtype : _GEN_632 ? _slots_35_io_uop_lrs2_rtype : _GEN_618 ? _slots_34_io_uop_lrs2_rtype : _GEN_604 ? _slots_33_io_uop_lrs2_rtype : _GEN_590 ? _slots_32_io_uop_lrs2_rtype : _GEN_576 ? _slots_31_io_uop_lrs2_rtype : _GEN_562 ? _slots_30_io_uop_lrs2_rtype : _GEN_548 ? _slots_29_io_uop_lrs2_rtype : _GEN_534 ? _slots_28_io_uop_lrs2_rtype : _GEN_520 ? _slots_27_io_uop_lrs2_rtype : _GEN_506 ? _slots_26_io_uop_lrs2_rtype : _GEN_492 ? _slots_25_io_uop_lrs2_rtype : _GEN_478 ? _slots_24_io_uop_lrs2_rtype : _GEN_464 ? _slots_23_io_uop_lrs2_rtype : _GEN_450 ? _slots_22_io_uop_lrs2_rtype : _GEN_436 ? _slots_21_io_uop_lrs2_rtype : _GEN_422 ? _slots_20_io_uop_lrs2_rtype : _GEN_408 ? _slots_19_io_uop_lrs2_rtype : _GEN_394 ? _slots_18_io_uop_lrs2_rtype : _GEN_380 ? _slots_17_io_uop_lrs2_rtype : _GEN_366 ? _slots_16_io_uop_lrs2_rtype : _GEN_352 ? _slots_15_io_uop_lrs2_rtype : _GEN_338 ? _slots_14_io_uop_lrs2_rtype : _GEN_324 ? _slots_13_io_uop_lrs2_rtype : _GEN_310 ? _slots_12_io_uop_lrs2_rtype : _GEN_296 ? _slots_11_io_uop_lrs2_rtype : _GEN_282 ? _slots_10_io_uop_lrs2_rtype : _GEN_268 ? _slots_9_io_uop_lrs2_rtype : _GEN_254 ? _slots_8_io_uop_lrs2_rtype : _GEN_240 ? _slots_7_io_uop_lrs2_rtype : _GEN_226 ? _slots_6_io_uop_lrs2_rtype : _GEN_212 ? _slots_5_io_uop_lrs2_rtype : _GEN_198 ? _slots_4_io_uop_lrs2_rtype : _GEN_184 ? _slots_3_io_uop_lrs2_rtype : _GEN_170 ? _slots_2_io_uop_lrs2_rtype : _GEN_156 ? _slots_1_io_uop_lrs2_rtype : _GEN_145 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_3_uopc = _GEN_682 ? _slots_39_io_uop_uopc : _GEN_676 ? _slots_38_io_uop_uopc : _GEN_663 ? _slots_37_io_uop_uopc : _GEN_649 ? _slots_36_io_uop_uopc : _GEN_635 ? _slots_35_io_uop_uopc : _GEN_621 ? _slots_34_io_uop_uopc : _GEN_607 ? _slots_33_io_uop_uopc : _GEN_593 ? _slots_32_io_uop_uopc : _GEN_579 ? _slots_31_io_uop_uopc : _GEN_565 ? _slots_30_io_uop_uopc : _GEN_551 ? _slots_29_io_uop_uopc : _GEN_537 ? _slots_28_io_uop_uopc : _GEN_523 ? _slots_27_io_uop_uopc : _GEN_509 ? _slots_26_io_uop_uopc : _GEN_495 ? _slots_25_io_uop_uopc : _GEN_481 ? _slots_24_io_uop_uopc : _GEN_467 ? _slots_23_io_uop_uopc : _GEN_453 ? _slots_22_io_uop_uopc : _GEN_439 ? _slots_21_io_uop_uopc : _GEN_425 ? _slots_20_io_uop_uopc : _GEN_411 ? _slots_19_io_uop_uopc : _GEN_397 ? _slots_18_io_uop_uopc : _GEN_383 ? _slots_17_io_uop_uopc : _GEN_369 ? _slots_16_io_uop_uopc : _GEN_355 ? _slots_15_io_uop_uopc : _GEN_341 ? _slots_14_io_uop_uopc : _GEN_327 ? _slots_13_io_uop_uopc : _GEN_313 ? _slots_12_io_uop_uopc : _GEN_299 ? _slots_11_io_uop_uopc : _GEN_285 ? _slots_10_io_uop_uopc : _GEN_271 ? _slots_9_io_uop_uopc : _GEN_257 ? _slots_8_io_uop_uopc : _GEN_243 ? _slots_7_io_uop_uopc : _GEN_229 ? _slots_6_io_uop_uopc : _GEN_215 ? _slots_5_io_uop_uopc : _GEN_201 ? _slots_4_io_uop_uopc : _GEN_187 ? _slots_3_io_uop_uopc : _GEN_173 ? _slots_2_io_uop_uopc : _GEN_159 ? _slots_1_io_uop_uopc : _GEN_146 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_3_is_rvc = _GEN_682 ? _slots_39_io_uop_is_rvc : _GEN_676 ? _slots_38_io_uop_is_rvc : _GEN_663 ? _slots_37_io_uop_is_rvc : _GEN_649 ? _slots_36_io_uop_is_rvc : _GEN_635 ? _slots_35_io_uop_is_rvc : _GEN_621 ? _slots_34_io_uop_is_rvc : _GEN_607 ? _slots_33_io_uop_is_rvc : _GEN_593 ? _slots_32_io_uop_is_rvc : _GEN_579 ? _slots_31_io_uop_is_rvc : _GEN_565 ? _slots_30_io_uop_is_rvc : _GEN_551 ? _slots_29_io_uop_is_rvc : _GEN_537 ? _slots_28_io_uop_is_rvc : _GEN_523 ? _slots_27_io_uop_is_rvc : _GEN_509 ? _slots_26_io_uop_is_rvc : _GEN_495 ? _slots_25_io_uop_is_rvc : _GEN_481 ? _slots_24_io_uop_is_rvc : _GEN_467 ? _slots_23_io_uop_is_rvc : _GEN_453 ? _slots_22_io_uop_is_rvc : _GEN_439 ? _slots_21_io_uop_is_rvc : _GEN_425 ? _slots_20_io_uop_is_rvc : _GEN_411 ? _slots_19_io_uop_is_rvc : _GEN_397 ? _slots_18_io_uop_is_rvc : _GEN_383 ? _slots_17_io_uop_is_rvc : _GEN_369 ? _slots_16_io_uop_is_rvc : _GEN_355 ? _slots_15_io_uop_is_rvc : _GEN_341 ? _slots_14_io_uop_is_rvc : _GEN_327 ? _slots_13_io_uop_is_rvc : _GEN_313 ? _slots_12_io_uop_is_rvc : _GEN_299 ? _slots_11_io_uop_is_rvc : _GEN_285 ? _slots_10_io_uop_is_rvc : _GEN_271 ? _slots_9_io_uop_is_rvc : _GEN_257 ? _slots_8_io_uop_is_rvc : _GEN_243 ? _slots_7_io_uop_is_rvc : _GEN_229 ? _slots_6_io_uop_is_rvc : _GEN_215 ? _slots_5_io_uop_is_rvc : _GEN_201 ? _slots_4_io_uop_is_rvc : _GEN_187 ? _slots_3_io_uop_is_rvc : _GEN_173 ? _slots_2_io_uop_is_rvc : _GEN_159 ? _slots_1_io_uop_is_rvc : _GEN_146 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_3_fu_code = _GEN_682 ? _slots_39_io_uop_fu_code : _GEN_676 ? _slots_38_io_uop_fu_code : _GEN_663 ? _slots_37_io_uop_fu_code : _GEN_649 ? _slots_36_io_uop_fu_code : _GEN_635 ? _slots_35_io_uop_fu_code : _GEN_621 ? _slots_34_io_uop_fu_code : _GEN_607 ? _slots_33_io_uop_fu_code : _GEN_593 ? _slots_32_io_uop_fu_code : _GEN_579 ? _slots_31_io_uop_fu_code : _GEN_565 ? _slots_30_io_uop_fu_code : _GEN_551 ? _slots_29_io_uop_fu_code : _GEN_537 ? _slots_28_io_uop_fu_code : _GEN_523 ? _slots_27_io_uop_fu_code : _GEN_509 ? _slots_26_io_uop_fu_code : _GEN_495 ? _slots_25_io_uop_fu_code : _GEN_481 ? _slots_24_io_uop_fu_code : _GEN_467 ? _slots_23_io_uop_fu_code : _GEN_453 ? _slots_22_io_uop_fu_code : _GEN_439 ? _slots_21_io_uop_fu_code : _GEN_425 ? _slots_20_io_uop_fu_code : _GEN_411 ? _slots_19_io_uop_fu_code : _GEN_397 ? _slots_18_io_uop_fu_code : _GEN_383 ? _slots_17_io_uop_fu_code : _GEN_369 ? _slots_16_io_uop_fu_code : _GEN_355 ? _slots_15_io_uop_fu_code : _GEN_341 ? _slots_14_io_uop_fu_code : _GEN_327 ? _slots_13_io_uop_fu_code : _GEN_313 ? _slots_12_io_uop_fu_code : _GEN_299 ? _slots_11_io_uop_fu_code : _GEN_285 ? _slots_10_io_uop_fu_code : _GEN_271 ? _slots_9_io_uop_fu_code : _GEN_257 ? _slots_8_io_uop_fu_code : _GEN_243 ? _slots_7_io_uop_fu_code : _GEN_229 ? _slots_6_io_uop_fu_code : _GEN_215 ? _slots_5_io_uop_fu_code : _GEN_201 ? _slots_4_io_uop_fu_code : _GEN_187 ? _slots_3_io_uop_fu_code : _GEN_173 ? _slots_2_io_uop_fu_code : _GEN_159 ? _slots_1_io_uop_fu_code : _GEN_146 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_3_iw_p1_poisoned = _GEN_682 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_676 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_663 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_649 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_635 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_621 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_607 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_593 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_579 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_565 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_551 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_537 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_523 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_509 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_495 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_481 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_467 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_453 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_439 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_425 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_411 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_397 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_383 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_369 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_355 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_341 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_327 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_313 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_299 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_285 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_271 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_257 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_243 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_229 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_215 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_201 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_187 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_173 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_159 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_146 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_3_iw_p2_poisoned = _GEN_682 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_676 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_663 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_649 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_635 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_621 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_607 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_593 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_579 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_565 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_551 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_537 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_523 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_509 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_495 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_481 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_467 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_453 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_439 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_425 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_411 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_397 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_383 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_369 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_355 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_341 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_327 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_313 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_299 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_285 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_271 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_257 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_243 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_229 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_215 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_201 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_187 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_173 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_159 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_146 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_3_is_br = _GEN_682 ? _slots_39_io_uop_is_br : _GEN_676 ? _slots_38_io_uop_is_br : _GEN_663 ? _slots_37_io_uop_is_br : _GEN_649 ? _slots_36_io_uop_is_br : _GEN_635 ? _slots_35_io_uop_is_br : _GEN_621 ? _slots_34_io_uop_is_br : _GEN_607 ? _slots_33_io_uop_is_br : _GEN_593 ? _slots_32_io_uop_is_br : _GEN_579 ? _slots_31_io_uop_is_br : _GEN_565 ? _slots_30_io_uop_is_br : _GEN_551 ? _slots_29_io_uop_is_br : _GEN_537 ? _slots_28_io_uop_is_br : _GEN_523 ? _slots_27_io_uop_is_br : _GEN_509 ? _slots_26_io_uop_is_br : _GEN_495 ? _slots_25_io_uop_is_br : _GEN_481 ? _slots_24_io_uop_is_br : _GEN_467 ? _slots_23_io_uop_is_br : _GEN_453 ? _slots_22_io_uop_is_br : _GEN_439 ? _slots_21_io_uop_is_br : _GEN_425 ? _slots_20_io_uop_is_br : _GEN_411 ? _slots_19_io_uop_is_br : _GEN_397 ? _slots_18_io_uop_is_br : _GEN_383 ? _slots_17_io_uop_is_br : _GEN_369 ? _slots_16_io_uop_is_br : _GEN_355 ? _slots_15_io_uop_is_br : _GEN_341 ? _slots_14_io_uop_is_br : _GEN_327 ? _slots_13_io_uop_is_br : _GEN_313 ? _slots_12_io_uop_is_br : _GEN_299 ? _slots_11_io_uop_is_br : _GEN_285 ? _slots_10_io_uop_is_br : _GEN_271 ? _slots_9_io_uop_is_br : _GEN_257 ? _slots_8_io_uop_is_br : _GEN_243 ? _slots_7_io_uop_is_br : _GEN_229 ? _slots_6_io_uop_is_br : _GEN_215 ? _slots_5_io_uop_is_br : _GEN_201 ? _slots_4_io_uop_is_br : _GEN_187 ? _slots_3_io_uop_is_br : _GEN_173 ? _slots_2_io_uop_is_br : _GEN_159 ? _slots_1_io_uop_is_br : _GEN_146 & _slots_0_io_uop_is_br;
  assign io_iss_uops_3_is_jalr = _GEN_682 ? _slots_39_io_uop_is_jalr : _GEN_676 ? _slots_38_io_uop_is_jalr : _GEN_663 ? _slots_37_io_uop_is_jalr : _GEN_649 ? _slots_36_io_uop_is_jalr : _GEN_635 ? _slots_35_io_uop_is_jalr : _GEN_621 ? _slots_34_io_uop_is_jalr : _GEN_607 ? _slots_33_io_uop_is_jalr : _GEN_593 ? _slots_32_io_uop_is_jalr : _GEN_579 ? _slots_31_io_uop_is_jalr : _GEN_565 ? _slots_30_io_uop_is_jalr : _GEN_551 ? _slots_29_io_uop_is_jalr : _GEN_537 ? _slots_28_io_uop_is_jalr : _GEN_523 ? _slots_27_io_uop_is_jalr : _GEN_509 ? _slots_26_io_uop_is_jalr : _GEN_495 ? _slots_25_io_uop_is_jalr : _GEN_481 ? _slots_24_io_uop_is_jalr : _GEN_467 ? _slots_23_io_uop_is_jalr : _GEN_453 ? _slots_22_io_uop_is_jalr : _GEN_439 ? _slots_21_io_uop_is_jalr : _GEN_425 ? _slots_20_io_uop_is_jalr : _GEN_411 ? _slots_19_io_uop_is_jalr : _GEN_397 ? _slots_18_io_uop_is_jalr : _GEN_383 ? _slots_17_io_uop_is_jalr : _GEN_369 ? _slots_16_io_uop_is_jalr : _GEN_355 ? _slots_15_io_uop_is_jalr : _GEN_341 ? _slots_14_io_uop_is_jalr : _GEN_327 ? _slots_13_io_uop_is_jalr : _GEN_313 ? _slots_12_io_uop_is_jalr : _GEN_299 ? _slots_11_io_uop_is_jalr : _GEN_285 ? _slots_10_io_uop_is_jalr : _GEN_271 ? _slots_9_io_uop_is_jalr : _GEN_257 ? _slots_8_io_uop_is_jalr : _GEN_243 ? _slots_7_io_uop_is_jalr : _GEN_229 ? _slots_6_io_uop_is_jalr : _GEN_215 ? _slots_5_io_uop_is_jalr : _GEN_201 ? _slots_4_io_uop_is_jalr : _GEN_187 ? _slots_3_io_uop_is_jalr : _GEN_173 ? _slots_2_io_uop_is_jalr : _GEN_159 ? _slots_1_io_uop_is_jalr : _GEN_146 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_3_is_jal = _GEN_682 ? _slots_39_io_uop_is_jal : _GEN_676 ? _slots_38_io_uop_is_jal : _GEN_663 ? _slots_37_io_uop_is_jal : _GEN_649 ? _slots_36_io_uop_is_jal : _GEN_635 ? _slots_35_io_uop_is_jal : _GEN_621 ? _slots_34_io_uop_is_jal : _GEN_607 ? _slots_33_io_uop_is_jal : _GEN_593 ? _slots_32_io_uop_is_jal : _GEN_579 ? _slots_31_io_uop_is_jal : _GEN_565 ? _slots_30_io_uop_is_jal : _GEN_551 ? _slots_29_io_uop_is_jal : _GEN_537 ? _slots_28_io_uop_is_jal : _GEN_523 ? _slots_27_io_uop_is_jal : _GEN_509 ? _slots_26_io_uop_is_jal : _GEN_495 ? _slots_25_io_uop_is_jal : _GEN_481 ? _slots_24_io_uop_is_jal : _GEN_467 ? _slots_23_io_uop_is_jal : _GEN_453 ? _slots_22_io_uop_is_jal : _GEN_439 ? _slots_21_io_uop_is_jal : _GEN_425 ? _slots_20_io_uop_is_jal : _GEN_411 ? _slots_19_io_uop_is_jal : _GEN_397 ? _slots_18_io_uop_is_jal : _GEN_383 ? _slots_17_io_uop_is_jal : _GEN_369 ? _slots_16_io_uop_is_jal : _GEN_355 ? _slots_15_io_uop_is_jal : _GEN_341 ? _slots_14_io_uop_is_jal : _GEN_327 ? _slots_13_io_uop_is_jal : _GEN_313 ? _slots_12_io_uop_is_jal : _GEN_299 ? _slots_11_io_uop_is_jal : _GEN_285 ? _slots_10_io_uop_is_jal : _GEN_271 ? _slots_9_io_uop_is_jal : _GEN_257 ? _slots_8_io_uop_is_jal : _GEN_243 ? _slots_7_io_uop_is_jal : _GEN_229 ? _slots_6_io_uop_is_jal : _GEN_215 ? _slots_5_io_uop_is_jal : _GEN_201 ? _slots_4_io_uop_is_jal : _GEN_187 ? _slots_3_io_uop_is_jal : _GEN_173 ? _slots_2_io_uop_is_jal : _GEN_159 ? _slots_1_io_uop_is_jal : _GEN_146 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_3_is_sfb = _GEN_682 ? _slots_39_io_uop_is_sfb : _GEN_676 ? _slots_38_io_uop_is_sfb : _GEN_663 ? _slots_37_io_uop_is_sfb : _GEN_649 ? _slots_36_io_uop_is_sfb : _GEN_635 ? _slots_35_io_uop_is_sfb : _GEN_621 ? _slots_34_io_uop_is_sfb : _GEN_607 ? _slots_33_io_uop_is_sfb : _GEN_593 ? _slots_32_io_uop_is_sfb : _GEN_579 ? _slots_31_io_uop_is_sfb : _GEN_565 ? _slots_30_io_uop_is_sfb : _GEN_551 ? _slots_29_io_uop_is_sfb : _GEN_537 ? _slots_28_io_uop_is_sfb : _GEN_523 ? _slots_27_io_uop_is_sfb : _GEN_509 ? _slots_26_io_uop_is_sfb : _GEN_495 ? _slots_25_io_uop_is_sfb : _GEN_481 ? _slots_24_io_uop_is_sfb : _GEN_467 ? _slots_23_io_uop_is_sfb : _GEN_453 ? _slots_22_io_uop_is_sfb : _GEN_439 ? _slots_21_io_uop_is_sfb : _GEN_425 ? _slots_20_io_uop_is_sfb : _GEN_411 ? _slots_19_io_uop_is_sfb : _GEN_397 ? _slots_18_io_uop_is_sfb : _GEN_383 ? _slots_17_io_uop_is_sfb : _GEN_369 ? _slots_16_io_uop_is_sfb : _GEN_355 ? _slots_15_io_uop_is_sfb : _GEN_341 ? _slots_14_io_uop_is_sfb : _GEN_327 ? _slots_13_io_uop_is_sfb : _GEN_313 ? _slots_12_io_uop_is_sfb : _GEN_299 ? _slots_11_io_uop_is_sfb : _GEN_285 ? _slots_10_io_uop_is_sfb : _GEN_271 ? _slots_9_io_uop_is_sfb : _GEN_257 ? _slots_8_io_uop_is_sfb : _GEN_243 ? _slots_7_io_uop_is_sfb : _GEN_229 ? _slots_6_io_uop_is_sfb : _GEN_215 ? _slots_5_io_uop_is_sfb : _GEN_201 ? _slots_4_io_uop_is_sfb : _GEN_187 ? _slots_3_io_uop_is_sfb : _GEN_173 ? _slots_2_io_uop_is_sfb : _GEN_159 ? _slots_1_io_uop_is_sfb : _GEN_146 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_3_br_mask = _GEN_682 ? _slots_39_io_uop_br_mask : _GEN_676 ? _slots_38_io_uop_br_mask : _GEN_663 ? _slots_37_io_uop_br_mask : _GEN_649 ? _slots_36_io_uop_br_mask : _GEN_635 ? _slots_35_io_uop_br_mask : _GEN_621 ? _slots_34_io_uop_br_mask : _GEN_607 ? _slots_33_io_uop_br_mask : _GEN_593 ? _slots_32_io_uop_br_mask : _GEN_579 ? _slots_31_io_uop_br_mask : _GEN_565 ? _slots_30_io_uop_br_mask : _GEN_551 ? _slots_29_io_uop_br_mask : _GEN_537 ? _slots_28_io_uop_br_mask : _GEN_523 ? _slots_27_io_uop_br_mask : _GEN_509 ? _slots_26_io_uop_br_mask : _GEN_495 ? _slots_25_io_uop_br_mask : _GEN_481 ? _slots_24_io_uop_br_mask : _GEN_467 ? _slots_23_io_uop_br_mask : _GEN_453 ? _slots_22_io_uop_br_mask : _GEN_439 ? _slots_21_io_uop_br_mask : _GEN_425 ? _slots_20_io_uop_br_mask : _GEN_411 ? _slots_19_io_uop_br_mask : _GEN_397 ? _slots_18_io_uop_br_mask : _GEN_383 ? _slots_17_io_uop_br_mask : _GEN_369 ? _slots_16_io_uop_br_mask : _GEN_355 ? _slots_15_io_uop_br_mask : _GEN_341 ? _slots_14_io_uop_br_mask : _GEN_327 ? _slots_13_io_uop_br_mask : _GEN_313 ? _slots_12_io_uop_br_mask : _GEN_299 ? _slots_11_io_uop_br_mask : _GEN_285 ? _slots_10_io_uop_br_mask : _GEN_271 ? _slots_9_io_uop_br_mask : _GEN_257 ? _slots_8_io_uop_br_mask : _GEN_243 ? _slots_7_io_uop_br_mask : _GEN_229 ? _slots_6_io_uop_br_mask : _GEN_215 ? _slots_5_io_uop_br_mask : _GEN_201 ? _slots_4_io_uop_br_mask : _GEN_187 ? _slots_3_io_uop_br_mask : _GEN_173 ? _slots_2_io_uop_br_mask : _GEN_159 ? _slots_1_io_uop_br_mask : _GEN_146 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_3_br_tag = _GEN_682 ? _slots_39_io_uop_br_tag : _GEN_676 ? _slots_38_io_uop_br_tag : _GEN_663 ? _slots_37_io_uop_br_tag : _GEN_649 ? _slots_36_io_uop_br_tag : _GEN_635 ? _slots_35_io_uop_br_tag : _GEN_621 ? _slots_34_io_uop_br_tag : _GEN_607 ? _slots_33_io_uop_br_tag : _GEN_593 ? _slots_32_io_uop_br_tag : _GEN_579 ? _slots_31_io_uop_br_tag : _GEN_565 ? _slots_30_io_uop_br_tag : _GEN_551 ? _slots_29_io_uop_br_tag : _GEN_537 ? _slots_28_io_uop_br_tag : _GEN_523 ? _slots_27_io_uop_br_tag : _GEN_509 ? _slots_26_io_uop_br_tag : _GEN_495 ? _slots_25_io_uop_br_tag : _GEN_481 ? _slots_24_io_uop_br_tag : _GEN_467 ? _slots_23_io_uop_br_tag : _GEN_453 ? _slots_22_io_uop_br_tag : _GEN_439 ? _slots_21_io_uop_br_tag : _GEN_425 ? _slots_20_io_uop_br_tag : _GEN_411 ? _slots_19_io_uop_br_tag : _GEN_397 ? _slots_18_io_uop_br_tag : _GEN_383 ? _slots_17_io_uop_br_tag : _GEN_369 ? _slots_16_io_uop_br_tag : _GEN_355 ? _slots_15_io_uop_br_tag : _GEN_341 ? _slots_14_io_uop_br_tag : _GEN_327 ? _slots_13_io_uop_br_tag : _GEN_313 ? _slots_12_io_uop_br_tag : _GEN_299 ? _slots_11_io_uop_br_tag : _GEN_285 ? _slots_10_io_uop_br_tag : _GEN_271 ? _slots_9_io_uop_br_tag : _GEN_257 ? _slots_8_io_uop_br_tag : _GEN_243 ? _slots_7_io_uop_br_tag : _GEN_229 ? _slots_6_io_uop_br_tag : _GEN_215 ? _slots_5_io_uop_br_tag : _GEN_201 ? _slots_4_io_uop_br_tag : _GEN_187 ? _slots_3_io_uop_br_tag : _GEN_173 ? _slots_2_io_uop_br_tag : _GEN_159 ? _slots_1_io_uop_br_tag : _GEN_146 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_3_ftq_idx = _GEN_682 ? _slots_39_io_uop_ftq_idx : _GEN_676 ? _slots_38_io_uop_ftq_idx : _GEN_663 ? _slots_37_io_uop_ftq_idx : _GEN_649 ? _slots_36_io_uop_ftq_idx : _GEN_635 ? _slots_35_io_uop_ftq_idx : _GEN_621 ? _slots_34_io_uop_ftq_idx : _GEN_607 ? _slots_33_io_uop_ftq_idx : _GEN_593 ? _slots_32_io_uop_ftq_idx : _GEN_579 ? _slots_31_io_uop_ftq_idx : _GEN_565 ? _slots_30_io_uop_ftq_idx : _GEN_551 ? _slots_29_io_uop_ftq_idx : _GEN_537 ? _slots_28_io_uop_ftq_idx : _GEN_523 ? _slots_27_io_uop_ftq_idx : _GEN_509 ? _slots_26_io_uop_ftq_idx : _GEN_495 ? _slots_25_io_uop_ftq_idx : _GEN_481 ? _slots_24_io_uop_ftq_idx : _GEN_467 ? _slots_23_io_uop_ftq_idx : _GEN_453 ? _slots_22_io_uop_ftq_idx : _GEN_439 ? _slots_21_io_uop_ftq_idx : _GEN_425 ? _slots_20_io_uop_ftq_idx : _GEN_411 ? _slots_19_io_uop_ftq_idx : _GEN_397 ? _slots_18_io_uop_ftq_idx : _GEN_383 ? _slots_17_io_uop_ftq_idx : _GEN_369 ? _slots_16_io_uop_ftq_idx : _GEN_355 ? _slots_15_io_uop_ftq_idx : _GEN_341 ? _slots_14_io_uop_ftq_idx : _GEN_327 ? _slots_13_io_uop_ftq_idx : _GEN_313 ? _slots_12_io_uop_ftq_idx : _GEN_299 ? _slots_11_io_uop_ftq_idx : _GEN_285 ? _slots_10_io_uop_ftq_idx : _GEN_271 ? _slots_9_io_uop_ftq_idx : _GEN_257 ? _slots_8_io_uop_ftq_idx : _GEN_243 ? _slots_7_io_uop_ftq_idx : _GEN_229 ? _slots_6_io_uop_ftq_idx : _GEN_215 ? _slots_5_io_uop_ftq_idx : _GEN_201 ? _slots_4_io_uop_ftq_idx : _GEN_187 ? _slots_3_io_uop_ftq_idx : _GEN_173 ? _slots_2_io_uop_ftq_idx : _GEN_159 ? _slots_1_io_uop_ftq_idx : _GEN_146 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_3_edge_inst = _GEN_682 ? _slots_39_io_uop_edge_inst : _GEN_676 ? _slots_38_io_uop_edge_inst : _GEN_663 ? _slots_37_io_uop_edge_inst : _GEN_649 ? _slots_36_io_uop_edge_inst : _GEN_635 ? _slots_35_io_uop_edge_inst : _GEN_621 ? _slots_34_io_uop_edge_inst : _GEN_607 ? _slots_33_io_uop_edge_inst : _GEN_593 ? _slots_32_io_uop_edge_inst : _GEN_579 ? _slots_31_io_uop_edge_inst : _GEN_565 ? _slots_30_io_uop_edge_inst : _GEN_551 ? _slots_29_io_uop_edge_inst : _GEN_537 ? _slots_28_io_uop_edge_inst : _GEN_523 ? _slots_27_io_uop_edge_inst : _GEN_509 ? _slots_26_io_uop_edge_inst : _GEN_495 ? _slots_25_io_uop_edge_inst : _GEN_481 ? _slots_24_io_uop_edge_inst : _GEN_467 ? _slots_23_io_uop_edge_inst : _GEN_453 ? _slots_22_io_uop_edge_inst : _GEN_439 ? _slots_21_io_uop_edge_inst : _GEN_425 ? _slots_20_io_uop_edge_inst : _GEN_411 ? _slots_19_io_uop_edge_inst : _GEN_397 ? _slots_18_io_uop_edge_inst : _GEN_383 ? _slots_17_io_uop_edge_inst : _GEN_369 ? _slots_16_io_uop_edge_inst : _GEN_355 ? _slots_15_io_uop_edge_inst : _GEN_341 ? _slots_14_io_uop_edge_inst : _GEN_327 ? _slots_13_io_uop_edge_inst : _GEN_313 ? _slots_12_io_uop_edge_inst : _GEN_299 ? _slots_11_io_uop_edge_inst : _GEN_285 ? _slots_10_io_uop_edge_inst : _GEN_271 ? _slots_9_io_uop_edge_inst : _GEN_257 ? _slots_8_io_uop_edge_inst : _GEN_243 ? _slots_7_io_uop_edge_inst : _GEN_229 ? _slots_6_io_uop_edge_inst : _GEN_215 ? _slots_5_io_uop_edge_inst : _GEN_201 ? _slots_4_io_uop_edge_inst : _GEN_187 ? _slots_3_io_uop_edge_inst : _GEN_173 ? _slots_2_io_uop_edge_inst : _GEN_159 ? _slots_1_io_uop_edge_inst : _GEN_146 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_3_pc_lob = _GEN_682 ? _slots_39_io_uop_pc_lob : _GEN_676 ? _slots_38_io_uop_pc_lob : _GEN_663 ? _slots_37_io_uop_pc_lob : _GEN_649 ? _slots_36_io_uop_pc_lob : _GEN_635 ? _slots_35_io_uop_pc_lob : _GEN_621 ? _slots_34_io_uop_pc_lob : _GEN_607 ? _slots_33_io_uop_pc_lob : _GEN_593 ? _slots_32_io_uop_pc_lob : _GEN_579 ? _slots_31_io_uop_pc_lob : _GEN_565 ? _slots_30_io_uop_pc_lob : _GEN_551 ? _slots_29_io_uop_pc_lob : _GEN_537 ? _slots_28_io_uop_pc_lob : _GEN_523 ? _slots_27_io_uop_pc_lob : _GEN_509 ? _slots_26_io_uop_pc_lob : _GEN_495 ? _slots_25_io_uop_pc_lob : _GEN_481 ? _slots_24_io_uop_pc_lob : _GEN_467 ? _slots_23_io_uop_pc_lob : _GEN_453 ? _slots_22_io_uop_pc_lob : _GEN_439 ? _slots_21_io_uop_pc_lob : _GEN_425 ? _slots_20_io_uop_pc_lob : _GEN_411 ? _slots_19_io_uop_pc_lob : _GEN_397 ? _slots_18_io_uop_pc_lob : _GEN_383 ? _slots_17_io_uop_pc_lob : _GEN_369 ? _slots_16_io_uop_pc_lob : _GEN_355 ? _slots_15_io_uop_pc_lob : _GEN_341 ? _slots_14_io_uop_pc_lob : _GEN_327 ? _slots_13_io_uop_pc_lob : _GEN_313 ? _slots_12_io_uop_pc_lob : _GEN_299 ? _slots_11_io_uop_pc_lob : _GEN_285 ? _slots_10_io_uop_pc_lob : _GEN_271 ? _slots_9_io_uop_pc_lob : _GEN_257 ? _slots_8_io_uop_pc_lob : _GEN_243 ? _slots_7_io_uop_pc_lob : _GEN_229 ? _slots_6_io_uop_pc_lob : _GEN_215 ? _slots_5_io_uop_pc_lob : _GEN_201 ? _slots_4_io_uop_pc_lob : _GEN_187 ? _slots_3_io_uop_pc_lob : _GEN_173 ? _slots_2_io_uop_pc_lob : _GEN_159 ? _slots_1_io_uop_pc_lob : _GEN_146 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_3_taken = _GEN_682 ? _slots_39_io_uop_taken : _GEN_676 ? _slots_38_io_uop_taken : _GEN_663 ? _slots_37_io_uop_taken : _GEN_649 ? _slots_36_io_uop_taken : _GEN_635 ? _slots_35_io_uop_taken : _GEN_621 ? _slots_34_io_uop_taken : _GEN_607 ? _slots_33_io_uop_taken : _GEN_593 ? _slots_32_io_uop_taken : _GEN_579 ? _slots_31_io_uop_taken : _GEN_565 ? _slots_30_io_uop_taken : _GEN_551 ? _slots_29_io_uop_taken : _GEN_537 ? _slots_28_io_uop_taken : _GEN_523 ? _slots_27_io_uop_taken : _GEN_509 ? _slots_26_io_uop_taken : _GEN_495 ? _slots_25_io_uop_taken : _GEN_481 ? _slots_24_io_uop_taken : _GEN_467 ? _slots_23_io_uop_taken : _GEN_453 ? _slots_22_io_uop_taken : _GEN_439 ? _slots_21_io_uop_taken : _GEN_425 ? _slots_20_io_uop_taken : _GEN_411 ? _slots_19_io_uop_taken : _GEN_397 ? _slots_18_io_uop_taken : _GEN_383 ? _slots_17_io_uop_taken : _GEN_369 ? _slots_16_io_uop_taken : _GEN_355 ? _slots_15_io_uop_taken : _GEN_341 ? _slots_14_io_uop_taken : _GEN_327 ? _slots_13_io_uop_taken : _GEN_313 ? _slots_12_io_uop_taken : _GEN_299 ? _slots_11_io_uop_taken : _GEN_285 ? _slots_10_io_uop_taken : _GEN_271 ? _slots_9_io_uop_taken : _GEN_257 ? _slots_8_io_uop_taken : _GEN_243 ? _slots_7_io_uop_taken : _GEN_229 ? _slots_6_io_uop_taken : _GEN_215 ? _slots_5_io_uop_taken : _GEN_201 ? _slots_4_io_uop_taken : _GEN_187 ? _slots_3_io_uop_taken : _GEN_173 ? _slots_2_io_uop_taken : _GEN_159 ? _slots_1_io_uop_taken : _GEN_146 & _slots_0_io_uop_taken;
  assign io_iss_uops_3_imm_packed = _GEN_682 ? _slots_39_io_uop_imm_packed : _GEN_676 ? _slots_38_io_uop_imm_packed : _GEN_663 ? _slots_37_io_uop_imm_packed : _GEN_649 ? _slots_36_io_uop_imm_packed : _GEN_635 ? _slots_35_io_uop_imm_packed : _GEN_621 ? _slots_34_io_uop_imm_packed : _GEN_607 ? _slots_33_io_uop_imm_packed : _GEN_593 ? _slots_32_io_uop_imm_packed : _GEN_579 ? _slots_31_io_uop_imm_packed : _GEN_565 ? _slots_30_io_uop_imm_packed : _GEN_551 ? _slots_29_io_uop_imm_packed : _GEN_537 ? _slots_28_io_uop_imm_packed : _GEN_523 ? _slots_27_io_uop_imm_packed : _GEN_509 ? _slots_26_io_uop_imm_packed : _GEN_495 ? _slots_25_io_uop_imm_packed : _GEN_481 ? _slots_24_io_uop_imm_packed : _GEN_467 ? _slots_23_io_uop_imm_packed : _GEN_453 ? _slots_22_io_uop_imm_packed : _GEN_439 ? _slots_21_io_uop_imm_packed : _GEN_425 ? _slots_20_io_uop_imm_packed : _GEN_411 ? _slots_19_io_uop_imm_packed : _GEN_397 ? _slots_18_io_uop_imm_packed : _GEN_383 ? _slots_17_io_uop_imm_packed : _GEN_369 ? _slots_16_io_uop_imm_packed : _GEN_355 ? _slots_15_io_uop_imm_packed : _GEN_341 ? _slots_14_io_uop_imm_packed : _GEN_327 ? _slots_13_io_uop_imm_packed : _GEN_313 ? _slots_12_io_uop_imm_packed : _GEN_299 ? _slots_11_io_uop_imm_packed : _GEN_285 ? _slots_10_io_uop_imm_packed : _GEN_271 ? _slots_9_io_uop_imm_packed : _GEN_257 ? _slots_8_io_uop_imm_packed : _GEN_243 ? _slots_7_io_uop_imm_packed : _GEN_229 ? _slots_6_io_uop_imm_packed : _GEN_215 ? _slots_5_io_uop_imm_packed : _GEN_201 ? _slots_4_io_uop_imm_packed : _GEN_187 ? _slots_3_io_uop_imm_packed : _GEN_173 ? _slots_2_io_uop_imm_packed : _GEN_159 ? _slots_1_io_uop_imm_packed : _GEN_146 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_3_rob_idx = _GEN_682 ? _slots_39_io_uop_rob_idx : _GEN_676 ? _slots_38_io_uop_rob_idx : _GEN_663 ? _slots_37_io_uop_rob_idx : _GEN_649 ? _slots_36_io_uop_rob_idx : _GEN_635 ? _slots_35_io_uop_rob_idx : _GEN_621 ? _slots_34_io_uop_rob_idx : _GEN_607 ? _slots_33_io_uop_rob_idx : _GEN_593 ? _slots_32_io_uop_rob_idx : _GEN_579 ? _slots_31_io_uop_rob_idx : _GEN_565 ? _slots_30_io_uop_rob_idx : _GEN_551 ? _slots_29_io_uop_rob_idx : _GEN_537 ? _slots_28_io_uop_rob_idx : _GEN_523 ? _slots_27_io_uop_rob_idx : _GEN_509 ? _slots_26_io_uop_rob_idx : _GEN_495 ? _slots_25_io_uop_rob_idx : _GEN_481 ? _slots_24_io_uop_rob_idx : _GEN_467 ? _slots_23_io_uop_rob_idx : _GEN_453 ? _slots_22_io_uop_rob_idx : _GEN_439 ? _slots_21_io_uop_rob_idx : _GEN_425 ? _slots_20_io_uop_rob_idx : _GEN_411 ? _slots_19_io_uop_rob_idx : _GEN_397 ? _slots_18_io_uop_rob_idx : _GEN_383 ? _slots_17_io_uop_rob_idx : _GEN_369 ? _slots_16_io_uop_rob_idx : _GEN_355 ? _slots_15_io_uop_rob_idx : _GEN_341 ? _slots_14_io_uop_rob_idx : _GEN_327 ? _slots_13_io_uop_rob_idx : _GEN_313 ? _slots_12_io_uop_rob_idx : _GEN_299 ? _slots_11_io_uop_rob_idx : _GEN_285 ? _slots_10_io_uop_rob_idx : _GEN_271 ? _slots_9_io_uop_rob_idx : _GEN_257 ? _slots_8_io_uop_rob_idx : _GEN_243 ? _slots_7_io_uop_rob_idx : _GEN_229 ? _slots_6_io_uop_rob_idx : _GEN_215 ? _slots_5_io_uop_rob_idx : _GEN_201 ? _slots_4_io_uop_rob_idx : _GEN_187 ? _slots_3_io_uop_rob_idx : _GEN_173 ? _slots_2_io_uop_rob_idx : _GEN_159 ? _slots_1_io_uop_rob_idx : _GEN_146 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_3_ldq_idx = _GEN_682 ? _slots_39_io_uop_ldq_idx : _GEN_676 ? _slots_38_io_uop_ldq_idx : _GEN_663 ? _slots_37_io_uop_ldq_idx : _GEN_649 ? _slots_36_io_uop_ldq_idx : _GEN_635 ? _slots_35_io_uop_ldq_idx : _GEN_621 ? _slots_34_io_uop_ldq_idx : _GEN_607 ? _slots_33_io_uop_ldq_idx : _GEN_593 ? _slots_32_io_uop_ldq_idx : _GEN_579 ? _slots_31_io_uop_ldq_idx : _GEN_565 ? _slots_30_io_uop_ldq_idx : _GEN_551 ? _slots_29_io_uop_ldq_idx : _GEN_537 ? _slots_28_io_uop_ldq_idx : _GEN_523 ? _slots_27_io_uop_ldq_idx : _GEN_509 ? _slots_26_io_uop_ldq_idx : _GEN_495 ? _slots_25_io_uop_ldq_idx : _GEN_481 ? _slots_24_io_uop_ldq_idx : _GEN_467 ? _slots_23_io_uop_ldq_idx : _GEN_453 ? _slots_22_io_uop_ldq_idx : _GEN_439 ? _slots_21_io_uop_ldq_idx : _GEN_425 ? _slots_20_io_uop_ldq_idx : _GEN_411 ? _slots_19_io_uop_ldq_idx : _GEN_397 ? _slots_18_io_uop_ldq_idx : _GEN_383 ? _slots_17_io_uop_ldq_idx : _GEN_369 ? _slots_16_io_uop_ldq_idx : _GEN_355 ? _slots_15_io_uop_ldq_idx : _GEN_341 ? _slots_14_io_uop_ldq_idx : _GEN_327 ? _slots_13_io_uop_ldq_idx : _GEN_313 ? _slots_12_io_uop_ldq_idx : _GEN_299 ? _slots_11_io_uop_ldq_idx : _GEN_285 ? _slots_10_io_uop_ldq_idx : _GEN_271 ? _slots_9_io_uop_ldq_idx : _GEN_257 ? _slots_8_io_uop_ldq_idx : _GEN_243 ? _slots_7_io_uop_ldq_idx : _GEN_229 ? _slots_6_io_uop_ldq_idx : _GEN_215 ? _slots_5_io_uop_ldq_idx : _GEN_201 ? _slots_4_io_uop_ldq_idx : _GEN_187 ? _slots_3_io_uop_ldq_idx : _GEN_173 ? _slots_2_io_uop_ldq_idx : _GEN_159 ? _slots_1_io_uop_ldq_idx : _GEN_146 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_3_stq_idx = _GEN_682 ? _slots_39_io_uop_stq_idx : _GEN_676 ? _slots_38_io_uop_stq_idx : _GEN_663 ? _slots_37_io_uop_stq_idx : _GEN_649 ? _slots_36_io_uop_stq_idx : _GEN_635 ? _slots_35_io_uop_stq_idx : _GEN_621 ? _slots_34_io_uop_stq_idx : _GEN_607 ? _slots_33_io_uop_stq_idx : _GEN_593 ? _slots_32_io_uop_stq_idx : _GEN_579 ? _slots_31_io_uop_stq_idx : _GEN_565 ? _slots_30_io_uop_stq_idx : _GEN_551 ? _slots_29_io_uop_stq_idx : _GEN_537 ? _slots_28_io_uop_stq_idx : _GEN_523 ? _slots_27_io_uop_stq_idx : _GEN_509 ? _slots_26_io_uop_stq_idx : _GEN_495 ? _slots_25_io_uop_stq_idx : _GEN_481 ? _slots_24_io_uop_stq_idx : _GEN_467 ? _slots_23_io_uop_stq_idx : _GEN_453 ? _slots_22_io_uop_stq_idx : _GEN_439 ? _slots_21_io_uop_stq_idx : _GEN_425 ? _slots_20_io_uop_stq_idx : _GEN_411 ? _slots_19_io_uop_stq_idx : _GEN_397 ? _slots_18_io_uop_stq_idx : _GEN_383 ? _slots_17_io_uop_stq_idx : _GEN_369 ? _slots_16_io_uop_stq_idx : _GEN_355 ? _slots_15_io_uop_stq_idx : _GEN_341 ? _slots_14_io_uop_stq_idx : _GEN_327 ? _slots_13_io_uop_stq_idx : _GEN_313 ? _slots_12_io_uop_stq_idx : _GEN_299 ? _slots_11_io_uop_stq_idx : _GEN_285 ? _slots_10_io_uop_stq_idx : _GEN_271 ? _slots_9_io_uop_stq_idx : _GEN_257 ? _slots_8_io_uop_stq_idx : _GEN_243 ? _slots_7_io_uop_stq_idx : _GEN_229 ? _slots_6_io_uop_stq_idx : _GEN_215 ? _slots_5_io_uop_stq_idx : _GEN_201 ? _slots_4_io_uop_stq_idx : _GEN_187 ? _slots_3_io_uop_stq_idx : _GEN_173 ? _slots_2_io_uop_stq_idx : _GEN_159 ? _slots_1_io_uop_stq_idx : _GEN_146 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_3_pdst = _GEN_682 ? _slots_39_io_uop_pdst : _GEN_676 ? _slots_38_io_uop_pdst : _GEN_663 ? _slots_37_io_uop_pdst : _GEN_649 ? _slots_36_io_uop_pdst : _GEN_635 ? _slots_35_io_uop_pdst : _GEN_621 ? _slots_34_io_uop_pdst : _GEN_607 ? _slots_33_io_uop_pdst : _GEN_593 ? _slots_32_io_uop_pdst : _GEN_579 ? _slots_31_io_uop_pdst : _GEN_565 ? _slots_30_io_uop_pdst : _GEN_551 ? _slots_29_io_uop_pdst : _GEN_537 ? _slots_28_io_uop_pdst : _GEN_523 ? _slots_27_io_uop_pdst : _GEN_509 ? _slots_26_io_uop_pdst : _GEN_495 ? _slots_25_io_uop_pdst : _GEN_481 ? _slots_24_io_uop_pdst : _GEN_467 ? _slots_23_io_uop_pdst : _GEN_453 ? _slots_22_io_uop_pdst : _GEN_439 ? _slots_21_io_uop_pdst : _GEN_425 ? _slots_20_io_uop_pdst : _GEN_411 ? _slots_19_io_uop_pdst : _GEN_397 ? _slots_18_io_uop_pdst : _GEN_383 ? _slots_17_io_uop_pdst : _GEN_369 ? _slots_16_io_uop_pdst : _GEN_355 ? _slots_15_io_uop_pdst : _GEN_341 ? _slots_14_io_uop_pdst : _GEN_327 ? _slots_13_io_uop_pdst : _GEN_313 ? _slots_12_io_uop_pdst : _GEN_299 ? _slots_11_io_uop_pdst : _GEN_285 ? _slots_10_io_uop_pdst : _GEN_271 ? _slots_9_io_uop_pdst : _GEN_257 ? _slots_8_io_uop_pdst : _GEN_243 ? _slots_7_io_uop_pdst : _GEN_229 ? _slots_6_io_uop_pdst : _GEN_215 ? _slots_5_io_uop_pdst : _GEN_201 ? _slots_4_io_uop_pdst : _GEN_187 ? _slots_3_io_uop_pdst : _GEN_173 ? _slots_2_io_uop_pdst : _GEN_159 ? _slots_1_io_uop_pdst : _GEN_146 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_3_prs1 = _GEN_682 ? _slots_39_io_uop_prs1 : _GEN_676 ? _slots_38_io_uop_prs1 : _GEN_663 ? _slots_37_io_uop_prs1 : _GEN_649 ? _slots_36_io_uop_prs1 : _GEN_635 ? _slots_35_io_uop_prs1 : _GEN_621 ? _slots_34_io_uop_prs1 : _GEN_607 ? _slots_33_io_uop_prs1 : _GEN_593 ? _slots_32_io_uop_prs1 : _GEN_579 ? _slots_31_io_uop_prs1 : _GEN_565 ? _slots_30_io_uop_prs1 : _GEN_551 ? _slots_29_io_uop_prs1 : _GEN_537 ? _slots_28_io_uop_prs1 : _GEN_523 ? _slots_27_io_uop_prs1 : _GEN_509 ? _slots_26_io_uop_prs1 : _GEN_495 ? _slots_25_io_uop_prs1 : _GEN_481 ? _slots_24_io_uop_prs1 : _GEN_467 ? _slots_23_io_uop_prs1 : _GEN_453 ? _slots_22_io_uop_prs1 : _GEN_439 ? _slots_21_io_uop_prs1 : _GEN_425 ? _slots_20_io_uop_prs1 : _GEN_411 ? _slots_19_io_uop_prs1 : _GEN_397 ? _slots_18_io_uop_prs1 : _GEN_383 ? _slots_17_io_uop_prs1 : _GEN_369 ? _slots_16_io_uop_prs1 : _GEN_355 ? _slots_15_io_uop_prs1 : _GEN_341 ? _slots_14_io_uop_prs1 : _GEN_327 ? _slots_13_io_uop_prs1 : _GEN_313 ? _slots_12_io_uop_prs1 : _GEN_299 ? _slots_11_io_uop_prs1 : _GEN_285 ? _slots_10_io_uop_prs1 : _GEN_271 ? _slots_9_io_uop_prs1 : _GEN_257 ? _slots_8_io_uop_prs1 : _GEN_243 ? _slots_7_io_uop_prs1 : _GEN_229 ? _slots_6_io_uop_prs1 : _GEN_215 ? _slots_5_io_uop_prs1 : _GEN_201 ? _slots_4_io_uop_prs1 : _GEN_187 ? _slots_3_io_uop_prs1 : _GEN_173 ? _slots_2_io_uop_prs1 : _GEN_159 ? _slots_1_io_uop_prs1 : _GEN_146 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_3_prs2 = _GEN_682 ? _slots_39_io_uop_prs2 : _GEN_676 ? _slots_38_io_uop_prs2 : _GEN_663 ? _slots_37_io_uop_prs2 : _GEN_649 ? _slots_36_io_uop_prs2 : _GEN_635 ? _slots_35_io_uop_prs2 : _GEN_621 ? _slots_34_io_uop_prs2 : _GEN_607 ? _slots_33_io_uop_prs2 : _GEN_593 ? _slots_32_io_uop_prs2 : _GEN_579 ? _slots_31_io_uop_prs2 : _GEN_565 ? _slots_30_io_uop_prs2 : _GEN_551 ? _slots_29_io_uop_prs2 : _GEN_537 ? _slots_28_io_uop_prs2 : _GEN_523 ? _slots_27_io_uop_prs2 : _GEN_509 ? _slots_26_io_uop_prs2 : _GEN_495 ? _slots_25_io_uop_prs2 : _GEN_481 ? _slots_24_io_uop_prs2 : _GEN_467 ? _slots_23_io_uop_prs2 : _GEN_453 ? _slots_22_io_uop_prs2 : _GEN_439 ? _slots_21_io_uop_prs2 : _GEN_425 ? _slots_20_io_uop_prs2 : _GEN_411 ? _slots_19_io_uop_prs2 : _GEN_397 ? _slots_18_io_uop_prs2 : _GEN_383 ? _slots_17_io_uop_prs2 : _GEN_369 ? _slots_16_io_uop_prs2 : _GEN_355 ? _slots_15_io_uop_prs2 : _GEN_341 ? _slots_14_io_uop_prs2 : _GEN_327 ? _slots_13_io_uop_prs2 : _GEN_313 ? _slots_12_io_uop_prs2 : _GEN_299 ? _slots_11_io_uop_prs2 : _GEN_285 ? _slots_10_io_uop_prs2 : _GEN_271 ? _slots_9_io_uop_prs2 : _GEN_257 ? _slots_8_io_uop_prs2 : _GEN_243 ? _slots_7_io_uop_prs2 : _GEN_229 ? _slots_6_io_uop_prs2 : _GEN_215 ? _slots_5_io_uop_prs2 : _GEN_201 ? _slots_4_io_uop_prs2 : _GEN_187 ? _slots_3_io_uop_prs2 : _GEN_173 ? _slots_2_io_uop_prs2 : _GEN_159 ? _slots_1_io_uop_prs2 : _GEN_146 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_3_bypassable = _GEN_682 ? _slots_39_io_uop_bypassable : _GEN_676 ? _slots_38_io_uop_bypassable : _GEN_663 ? _slots_37_io_uop_bypassable : _GEN_649 ? _slots_36_io_uop_bypassable : _GEN_635 ? _slots_35_io_uop_bypassable : _GEN_621 ? _slots_34_io_uop_bypassable : _GEN_607 ? _slots_33_io_uop_bypassable : _GEN_593 ? _slots_32_io_uop_bypassable : _GEN_579 ? _slots_31_io_uop_bypassable : _GEN_565 ? _slots_30_io_uop_bypassable : _GEN_551 ? _slots_29_io_uop_bypassable : _GEN_537 ? _slots_28_io_uop_bypassable : _GEN_523 ? _slots_27_io_uop_bypassable : _GEN_509 ? _slots_26_io_uop_bypassable : _GEN_495 ? _slots_25_io_uop_bypassable : _GEN_481 ? _slots_24_io_uop_bypassable : _GEN_467 ? _slots_23_io_uop_bypassable : _GEN_453 ? _slots_22_io_uop_bypassable : _GEN_439 ? _slots_21_io_uop_bypassable : _GEN_425 ? _slots_20_io_uop_bypassable : _GEN_411 ? _slots_19_io_uop_bypassable : _GEN_397 ? _slots_18_io_uop_bypassable : _GEN_383 ? _slots_17_io_uop_bypassable : _GEN_369 ? _slots_16_io_uop_bypassable : _GEN_355 ? _slots_15_io_uop_bypassable : _GEN_341 ? _slots_14_io_uop_bypassable : _GEN_327 ? _slots_13_io_uop_bypassable : _GEN_313 ? _slots_12_io_uop_bypassable : _GEN_299 ? _slots_11_io_uop_bypassable : _GEN_285 ? _slots_10_io_uop_bypassable : _GEN_271 ? _slots_9_io_uop_bypassable : _GEN_257 ? _slots_8_io_uop_bypassable : _GEN_243 ? _slots_7_io_uop_bypassable : _GEN_229 ? _slots_6_io_uop_bypassable : _GEN_215 ? _slots_5_io_uop_bypassable : _GEN_201 ? _slots_4_io_uop_bypassable : _GEN_187 ? _slots_3_io_uop_bypassable : _GEN_173 ? _slots_2_io_uop_bypassable : _GEN_159 ? _slots_1_io_uop_bypassable : _GEN_146 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_3_mem_cmd = _GEN_682 ? _slots_39_io_uop_mem_cmd : _GEN_676 ? _slots_38_io_uop_mem_cmd : _GEN_663 ? _slots_37_io_uop_mem_cmd : _GEN_649 ? _slots_36_io_uop_mem_cmd : _GEN_635 ? _slots_35_io_uop_mem_cmd : _GEN_621 ? _slots_34_io_uop_mem_cmd : _GEN_607 ? _slots_33_io_uop_mem_cmd : _GEN_593 ? _slots_32_io_uop_mem_cmd : _GEN_579 ? _slots_31_io_uop_mem_cmd : _GEN_565 ? _slots_30_io_uop_mem_cmd : _GEN_551 ? _slots_29_io_uop_mem_cmd : _GEN_537 ? _slots_28_io_uop_mem_cmd : _GEN_523 ? _slots_27_io_uop_mem_cmd : _GEN_509 ? _slots_26_io_uop_mem_cmd : _GEN_495 ? _slots_25_io_uop_mem_cmd : _GEN_481 ? _slots_24_io_uop_mem_cmd : _GEN_467 ? _slots_23_io_uop_mem_cmd : _GEN_453 ? _slots_22_io_uop_mem_cmd : _GEN_439 ? _slots_21_io_uop_mem_cmd : _GEN_425 ? _slots_20_io_uop_mem_cmd : _GEN_411 ? _slots_19_io_uop_mem_cmd : _GEN_397 ? _slots_18_io_uop_mem_cmd : _GEN_383 ? _slots_17_io_uop_mem_cmd : _GEN_369 ? _slots_16_io_uop_mem_cmd : _GEN_355 ? _slots_15_io_uop_mem_cmd : _GEN_341 ? _slots_14_io_uop_mem_cmd : _GEN_327 ? _slots_13_io_uop_mem_cmd : _GEN_313 ? _slots_12_io_uop_mem_cmd : _GEN_299 ? _slots_11_io_uop_mem_cmd : _GEN_285 ? _slots_10_io_uop_mem_cmd : _GEN_271 ? _slots_9_io_uop_mem_cmd : _GEN_257 ? _slots_8_io_uop_mem_cmd : _GEN_243 ? _slots_7_io_uop_mem_cmd : _GEN_229 ? _slots_6_io_uop_mem_cmd : _GEN_215 ? _slots_5_io_uop_mem_cmd : _GEN_201 ? _slots_4_io_uop_mem_cmd : _GEN_187 ? _slots_3_io_uop_mem_cmd : _GEN_173 ? _slots_2_io_uop_mem_cmd : _GEN_159 ? _slots_1_io_uop_mem_cmd : _GEN_146 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_3_is_amo = _GEN_682 ? _slots_39_io_uop_is_amo : _GEN_676 ? _slots_38_io_uop_is_amo : _GEN_663 ? _slots_37_io_uop_is_amo : _GEN_649 ? _slots_36_io_uop_is_amo : _GEN_635 ? _slots_35_io_uop_is_amo : _GEN_621 ? _slots_34_io_uop_is_amo : _GEN_607 ? _slots_33_io_uop_is_amo : _GEN_593 ? _slots_32_io_uop_is_amo : _GEN_579 ? _slots_31_io_uop_is_amo : _GEN_565 ? _slots_30_io_uop_is_amo : _GEN_551 ? _slots_29_io_uop_is_amo : _GEN_537 ? _slots_28_io_uop_is_amo : _GEN_523 ? _slots_27_io_uop_is_amo : _GEN_509 ? _slots_26_io_uop_is_amo : _GEN_495 ? _slots_25_io_uop_is_amo : _GEN_481 ? _slots_24_io_uop_is_amo : _GEN_467 ? _slots_23_io_uop_is_amo : _GEN_453 ? _slots_22_io_uop_is_amo : _GEN_439 ? _slots_21_io_uop_is_amo : _GEN_425 ? _slots_20_io_uop_is_amo : _GEN_411 ? _slots_19_io_uop_is_amo : _GEN_397 ? _slots_18_io_uop_is_amo : _GEN_383 ? _slots_17_io_uop_is_amo : _GEN_369 ? _slots_16_io_uop_is_amo : _GEN_355 ? _slots_15_io_uop_is_amo : _GEN_341 ? _slots_14_io_uop_is_amo : _GEN_327 ? _slots_13_io_uop_is_amo : _GEN_313 ? _slots_12_io_uop_is_amo : _GEN_299 ? _slots_11_io_uop_is_amo : _GEN_285 ? _slots_10_io_uop_is_amo : _GEN_271 ? _slots_9_io_uop_is_amo : _GEN_257 ? _slots_8_io_uop_is_amo : _GEN_243 ? _slots_7_io_uop_is_amo : _GEN_229 ? _slots_6_io_uop_is_amo : _GEN_215 ? _slots_5_io_uop_is_amo : _GEN_201 ? _slots_4_io_uop_is_amo : _GEN_187 ? _slots_3_io_uop_is_amo : _GEN_173 ? _slots_2_io_uop_is_amo : _GEN_159 ? _slots_1_io_uop_is_amo : _GEN_146 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_3_uses_stq = _GEN_682 ? _slots_39_io_uop_uses_stq : _GEN_676 ? _slots_38_io_uop_uses_stq : _GEN_663 ? _slots_37_io_uop_uses_stq : _GEN_649 ? _slots_36_io_uop_uses_stq : _GEN_635 ? _slots_35_io_uop_uses_stq : _GEN_621 ? _slots_34_io_uop_uses_stq : _GEN_607 ? _slots_33_io_uop_uses_stq : _GEN_593 ? _slots_32_io_uop_uses_stq : _GEN_579 ? _slots_31_io_uop_uses_stq : _GEN_565 ? _slots_30_io_uop_uses_stq : _GEN_551 ? _slots_29_io_uop_uses_stq : _GEN_537 ? _slots_28_io_uop_uses_stq : _GEN_523 ? _slots_27_io_uop_uses_stq : _GEN_509 ? _slots_26_io_uop_uses_stq : _GEN_495 ? _slots_25_io_uop_uses_stq : _GEN_481 ? _slots_24_io_uop_uses_stq : _GEN_467 ? _slots_23_io_uop_uses_stq : _GEN_453 ? _slots_22_io_uop_uses_stq : _GEN_439 ? _slots_21_io_uop_uses_stq : _GEN_425 ? _slots_20_io_uop_uses_stq : _GEN_411 ? _slots_19_io_uop_uses_stq : _GEN_397 ? _slots_18_io_uop_uses_stq : _GEN_383 ? _slots_17_io_uop_uses_stq : _GEN_369 ? _slots_16_io_uop_uses_stq : _GEN_355 ? _slots_15_io_uop_uses_stq : _GEN_341 ? _slots_14_io_uop_uses_stq : _GEN_327 ? _slots_13_io_uop_uses_stq : _GEN_313 ? _slots_12_io_uop_uses_stq : _GEN_299 ? _slots_11_io_uop_uses_stq : _GEN_285 ? _slots_10_io_uop_uses_stq : _GEN_271 ? _slots_9_io_uop_uses_stq : _GEN_257 ? _slots_8_io_uop_uses_stq : _GEN_243 ? _slots_7_io_uop_uses_stq : _GEN_229 ? _slots_6_io_uop_uses_stq : _GEN_215 ? _slots_5_io_uop_uses_stq : _GEN_201 ? _slots_4_io_uop_uses_stq : _GEN_187 ? _slots_3_io_uop_uses_stq : _GEN_173 ? _slots_2_io_uop_uses_stq : _GEN_159 ? _slots_1_io_uop_uses_stq : _GEN_146 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_3_ldst_val = _GEN_682 ? _slots_39_io_uop_ldst_val : _GEN_676 ? _slots_38_io_uop_ldst_val : _GEN_663 ? _slots_37_io_uop_ldst_val : _GEN_649 ? _slots_36_io_uop_ldst_val : _GEN_635 ? _slots_35_io_uop_ldst_val : _GEN_621 ? _slots_34_io_uop_ldst_val : _GEN_607 ? _slots_33_io_uop_ldst_val : _GEN_593 ? _slots_32_io_uop_ldst_val : _GEN_579 ? _slots_31_io_uop_ldst_val : _GEN_565 ? _slots_30_io_uop_ldst_val : _GEN_551 ? _slots_29_io_uop_ldst_val : _GEN_537 ? _slots_28_io_uop_ldst_val : _GEN_523 ? _slots_27_io_uop_ldst_val : _GEN_509 ? _slots_26_io_uop_ldst_val : _GEN_495 ? _slots_25_io_uop_ldst_val : _GEN_481 ? _slots_24_io_uop_ldst_val : _GEN_467 ? _slots_23_io_uop_ldst_val : _GEN_453 ? _slots_22_io_uop_ldst_val : _GEN_439 ? _slots_21_io_uop_ldst_val : _GEN_425 ? _slots_20_io_uop_ldst_val : _GEN_411 ? _slots_19_io_uop_ldst_val : _GEN_397 ? _slots_18_io_uop_ldst_val : _GEN_383 ? _slots_17_io_uop_ldst_val : _GEN_369 ? _slots_16_io_uop_ldst_val : _GEN_355 ? _slots_15_io_uop_ldst_val : _GEN_341 ? _slots_14_io_uop_ldst_val : _GEN_327 ? _slots_13_io_uop_ldst_val : _GEN_313 ? _slots_12_io_uop_ldst_val : _GEN_299 ? _slots_11_io_uop_ldst_val : _GEN_285 ? _slots_10_io_uop_ldst_val : _GEN_271 ? _slots_9_io_uop_ldst_val : _GEN_257 ? _slots_8_io_uop_ldst_val : _GEN_243 ? _slots_7_io_uop_ldst_val : _GEN_229 ? _slots_6_io_uop_ldst_val : _GEN_215 ? _slots_5_io_uop_ldst_val : _GEN_201 ? _slots_4_io_uop_ldst_val : _GEN_187 ? _slots_3_io_uop_ldst_val : _GEN_173 ? _slots_2_io_uop_ldst_val : _GEN_159 ? _slots_1_io_uop_ldst_val : _GEN_146 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_3_dst_rtype = _GEN_682 ? _slots_39_io_uop_dst_rtype : _GEN_676 ? _slots_38_io_uop_dst_rtype : _GEN_663 ? _slots_37_io_uop_dst_rtype : _GEN_649 ? _slots_36_io_uop_dst_rtype : _GEN_635 ? _slots_35_io_uop_dst_rtype : _GEN_621 ? _slots_34_io_uop_dst_rtype : _GEN_607 ? _slots_33_io_uop_dst_rtype : _GEN_593 ? _slots_32_io_uop_dst_rtype : _GEN_579 ? _slots_31_io_uop_dst_rtype : _GEN_565 ? _slots_30_io_uop_dst_rtype : _GEN_551 ? _slots_29_io_uop_dst_rtype : _GEN_537 ? _slots_28_io_uop_dst_rtype : _GEN_523 ? _slots_27_io_uop_dst_rtype : _GEN_509 ? _slots_26_io_uop_dst_rtype : _GEN_495 ? _slots_25_io_uop_dst_rtype : _GEN_481 ? _slots_24_io_uop_dst_rtype : _GEN_467 ? _slots_23_io_uop_dst_rtype : _GEN_453 ? _slots_22_io_uop_dst_rtype : _GEN_439 ? _slots_21_io_uop_dst_rtype : _GEN_425 ? _slots_20_io_uop_dst_rtype : _GEN_411 ? _slots_19_io_uop_dst_rtype : _GEN_397 ? _slots_18_io_uop_dst_rtype : _GEN_383 ? _slots_17_io_uop_dst_rtype : _GEN_369 ? _slots_16_io_uop_dst_rtype : _GEN_355 ? _slots_15_io_uop_dst_rtype : _GEN_341 ? _slots_14_io_uop_dst_rtype : _GEN_327 ? _slots_13_io_uop_dst_rtype : _GEN_313 ? _slots_12_io_uop_dst_rtype : _GEN_299 ? _slots_11_io_uop_dst_rtype : _GEN_285 ? _slots_10_io_uop_dst_rtype : _GEN_271 ? _slots_9_io_uop_dst_rtype : _GEN_257 ? _slots_8_io_uop_dst_rtype : _GEN_243 ? _slots_7_io_uop_dst_rtype : _GEN_229 ? _slots_6_io_uop_dst_rtype : _GEN_215 ? _slots_5_io_uop_dst_rtype : _GEN_201 ? _slots_4_io_uop_dst_rtype : _GEN_187 ? _slots_3_io_uop_dst_rtype : _GEN_173 ? _slots_2_io_uop_dst_rtype : _GEN_159 ? _slots_1_io_uop_dst_rtype : _GEN_146 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_3_lrs1_rtype = _GEN_682 ? _slots_39_io_uop_lrs1_rtype : _GEN_676 ? _slots_38_io_uop_lrs1_rtype : _GEN_663 ? _slots_37_io_uop_lrs1_rtype : _GEN_649 ? _slots_36_io_uop_lrs1_rtype : _GEN_635 ? _slots_35_io_uop_lrs1_rtype : _GEN_621 ? _slots_34_io_uop_lrs1_rtype : _GEN_607 ? _slots_33_io_uop_lrs1_rtype : _GEN_593 ? _slots_32_io_uop_lrs1_rtype : _GEN_579 ? _slots_31_io_uop_lrs1_rtype : _GEN_565 ? _slots_30_io_uop_lrs1_rtype : _GEN_551 ? _slots_29_io_uop_lrs1_rtype : _GEN_537 ? _slots_28_io_uop_lrs1_rtype : _GEN_523 ? _slots_27_io_uop_lrs1_rtype : _GEN_509 ? _slots_26_io_uop_lrs1_rtype : _GEN_495 ? _slots_25_io_uop_lrs1_rtype : _GEN_481 ? _slots_24_io_uop_lrs1_rtype : _GEN_467 ? _slots_23_io_uop_lrs1_rtype : _GEN_453 ? _slots_22_io_uop_lrs1_rtype : _GEN_439 ? _slots_21_io_uop_lrs1_rtype : _GEN_425 ? _slots_20_io_uop_lrs1_rtype : _GEN_411 ? _slots_19_io_uop_lrs1_rtype : _GEN_397 ? _slots_18_io_uop_lrs1_rtype : _GEN_383 ? _slots_17_io_uop_lrs1_rtype : _GEN_369 ? _slots_16_io_uop_lrs1_rtype : _GEN_355 ? _slots_15_io_uop_lrs1_rtype : _GEN_341 ? _slots_14_io_uop_lrs1_rtype : _GEN_327 ? _slots_13_io_uop_lrs1_rtype : _GEN_313 ? _slots_12_io_uop_lrs1_rtype : _GEN_299 ? _slots_11_io_uop_lrs1_rtype : _GEN_285 ? _slots_10_io_uop_lrs1_rtype : _GEN_271 ? _slots_9_io_uop_lrs1_rtype : _GEN_257 ? _slots_8_io_uop_lrs1_rtype : _GEN_243 ? _slots_7_io_uop_lrs1_rtype : _GEN_229 ? _slots_6_io_uop_lrs1_rtype : _GEN_215 ? _slots_5_io_uop_lrs1_rtype : _GEN_201 ? _slots_4_io_uop_lrs1_rtype : _GEN_187 ? _slots_3_io_uop_lrs1_rtype : _GEN_173 ? _slots_2_io_uop_lrs1_rtype : _GEN_159 ? _slots_1_io_uop_lrs1_rtype : _GEN_146 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_3_lrs2_rtype = _GEN_682 ? _slots_39_io_uop_lrs2_rtype : _GEN_676 ? _slots_38_io_uop_lrs2_rtype : _GEN_663 ? _slots_37_io_uop_lrs2_rtype : _GEN_649 ? _slots_36_io_uop_lrs2_rtype : _GEN_635 ? _slots_35_io_uop_lrs2_rtype : _GEN_621 ? _slots_34_io_uop_lrs2_rtype : _GEN_607 ? _slots_33_io_uop_lrs2_rtype : _GEN_593 ? _slots_32_io_uop_lrs2_rtype : _GEN_579 ? _slots_31_io_uop_lrs2_rtype : _GEN_565 ? _slots_30_io_uop_lrs2_rtype : _GEN_551 ? _slots_29_io_uop_lrs2_rtype : _GEN_537 ? _slots_28_io_uop_lrs2_rtype : _GEN_523 ? _slots_27_io_uop_lrs2_rtype : _GEN_509 ? _slots_26_io_uop_lrs2_rtype : _GEN_495 ? _slots_25_io_uop_lrs2_rtype : _GEN_481 ? _slots_24_io_uop_lrs2_rtype : _GEN_467 ? _slots_23_io_uop_lrs2_rtype : _GEN_453 ? _slots_22_io_uop_lrs2_rtype : _GEN_439 ? _slots_21_io_uop_lrs2_rtype : _GEN_425 ? _slots_20_io_uop_lrs2_rtype : _GEN_411 ? _slots_19_io_uop_lrs2_rtype : _GEN_397 ? _slots_18_io_uop_lrs2_rtype : _GEN_383 ? _slots_17_io_uop_lrs2_rtype : _GEN_369 ? _slots_16_io_uop_lrs2_rtype : _GEN_355 ? _slots_15_io_uop_lrs2_rtype : _GEN_341 ? _slots_14_io_uop_lrs2_rtype : _GEN_327 ? _slots_13_io_uop_lrs2_rtype : _GEN_313 ? _slots_12_io_uop_lrs2_rtype : _GEN_299 ? _slots_11_io_uop_lrs2_rtype : _GEN_285 ? _slots_10_io_uop_lrs2_rtype : _GEN_271 ? _slots_9_io_uop_lrs2_rtype : _GEN_257 ? _slots_8_io_uop_lrs2_rtype : _GEN_243 ? _slots_7_io_uop_lrs2_rtype : _GEN_229 ? _slots_6_io_uop_lrs2_rtype : _GEN_215 ? _slots_5_io_uop_lrs2_rtype : _GEN_201 ? _slots_4_io_uop_lrs2_rtype : _GEN_187 ? _slots_3_io_uop_lrs2_rtype : _GEN_173 ? _slots_2_io_uop_lrs2_rtype : _GEN_159 ? _slots_1_io_uop_lrs2_rtype : _GEN_146 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
endmodule

