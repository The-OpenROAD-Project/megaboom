// Standard header to adapt well known macros for prints and assertions.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module LSU(
  input         clock,
                reset,
                io_ptw_req_ready,
  output        io_ptw_req_valid,
                io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
                io_ptw_resp_bits_ae_final,
  input  [43:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
                io_ptw_resp_bits_pte_a,
                io_ptw_resp_bits_pte_g,
                io_ptw_resp_bits_pte_u,
                io_ptw_resp_bits_pte_x,
                io_ptw_resp_bits_pte_w,
                io_ptw_resp_bits_pte_r,
                io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
                io_ptw_status_sum,
                io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
                io_ptw_pmp_0_cfg_w,
                io_ptw_pmp_0_cfg_r,
  input  [30:0] io_ptw_pmp_0_addr,
  input  [32:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
                io_ptw_pmp_1_cfg_w,
                io_ptw_pmp_1_cfg_r,
  input  [30:0] io_ptw_pmp_1_addr,
  input  [32:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
                io_ptw_pmp_2_cfg_w,
                io_ptw_pmp_2_cfg_r,
  input  [30:0] io_ptw_pmp_2_addr,
  input  [32:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
                io_ptw_pmp_3_cfg_w,
                io_ptw_pmp_3_cfg_r,
  input  [30:0] io_ptw_pmp_3_addr,
  input  [32:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
                io_ptw_pmp_4_cfg_w,
                io_ptw_pmp_4_cfg_r,
  input  [30:0] io_ptw_pmp_4_addr,
  input  [32:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
                io_ptw_pmp_5_cfg_w,
                io_ptw_pmp_5_cfg_r,
  input  [30:0] io_ptw_pmp_5_addr,
  input  [32:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
                io_ptw_pmp_6_cfg_w,
                io_ptw_pmp_6_cfg_r,
  input  [30:0] io_ptw_pmp_6_addr,
  input  [32:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
                io_ptw_pmp_7_cfg_w,
                io_ptw_pmp_7_cfg_r,
  input  [30:0] io_ptw_pmp_7_addr,
  input  [32:0] io_ptw_pmp_7_mask,
  input         io_core_exe_0_req_valid,
  input  [6:0]  io_core_exe_0_req_bits_uop_uopc,
  input  [31:0] io_core_exe_0_req_bits_uop_inst,
                io_core_exe_0_req_bits_uop_debug_inst,
  input         io_core_exe_0_req_bits_uop_is_rvc,
  input  [39:0] io_core_exe_0_req_bits_uop_debug_pc,
  input  [2:0]  io_core_exe_0_req_bits_uop_iq_type,
  input  [9:0]  io_core_exe_0_req_bits_uop_fu_code,
  input  [3:0]  io_core_exe_0_req_bits_uop_ctrl_br_type,
  input  [1:0]  io_core_exe_0_req_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_core_exe_0_req_bits_uop_ctrl_op2_sel,
                io_core_exe_0_req_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_core_exe_0_req_bits_uop_ctrl_op_fcn,
  input         io_core_exe_0_req_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_core_exe_0_req_bits_uop_ctrl_csr_cmd,
  input         io_core_exe_0_req_bits_uop_ctrl_is_load,
                io_core_exe_0_req_bits_uop_ctrl_is_sta,
                io_core_exe_0_req_bits_uop_ctrl_is_std,
  input  [1:0]  io_core_exe_0_req_bits_uop_iw_state,
  input         io_core_exe_0_req_bits_uop_is_br,
                io_core_exe_0_req_bits_uop_is_jalr,
                io_core_exe_0_req_bits_uop_is_jal,
                io_core_exe_0_req_bits_uop_is_sfb,
  input  [19:0] io_core_exe_0_req_bits_uop_br_mask,
  input  [4:0]  io_core_exe_0_req_bits_uop_br_tag,
  input  [5:0]  io_core_exe_0_req_bits_uop_ftq_idx,
  input         io_core_exe_0_req_bits_uop_edge_inst,
  input  [5:0]  io_core_exe_0_req_bits_uop_pc_lob,
  input         io_core_exe_0_req_bits_uop_taken,
  input  [19:0] io_core_exe_0_req_bits_uop_imm_packed,
  input  [11:0] io_core_exe_0_req_bits_uop_csr_addr,
  input  [6:0]  io_core_exe_0_req_bits_uop_rob_idx,
  input  [4:0]  io_core_exe_0_req_bits_uop_ldq_idx,
                io_core_exe_0_req_bits_uop_stq_idx,
  input  [1:0]  io_core_exe_0_req_bits_uop_rxq_idx,
  input  [6:0]  io_core_exe_0_req_bits_uop_pdst,
                io_core_exe_0_req_bits_uop_prs1,
                io_core_exe_0_req_bits_uop_prs2,
                io_core_exe_0_req_bits_uop_prs3,
  input  [5:0]  io_core_exe_0_req_bits_uop_ppred,
  input         io_core_exe_0_req_bits_uop_prs1_busy,
                io_core_exe_0_req_bits_uop_prs2_busy,
                io_core_exe_0_req_bits_uop_prs3_busy,
                io_core_exe_0_req_bits_uop_ppred_busy,
  input  [6:0]  io_core_exe_0_req_bits_uop_stale_pdst,
  input         io_core_exe_0_req_bits_uop_exception,
  input  [63:0] io_core_exe_0_req_bits_uop_exc_cause,
  input         io_core_exe_0_req_bits_uop_bypassable,
  input  [4:0]  io_core_exe_0_req_bits_uop_mem_cmd,
  input  [1:0]  io_core_exe_0_req_bits_uop_mem_size,
  input         io_core_exe_0_req_bits_uop_mem_signed,
                io_core_exe_0_req_bits_uop_is_fence,
                io_core_exe_0_req_bits_uop_is_fencei,
                io_core_exe_0_req_bits_uop_is_amo,
                io_core_exe_0_req_bits_uop_uses_ldq,
                io_core_exe_0_req_bits_uop_uses_stq,
                io_core_exe_0_req_bits_uop_is_sys_pc2epc,
                io_core_exe_0_req_bits_uop_is_unique,
                io_core_exe_0_req_bits_uop_flush_on_commit,
                io_core_exe_0_req_bits_uop_ldst_is_rs1,
  input  [5:0]  io_core_exe_0_req_bits_uop_ldst,
                io_core_exe_0_req_bits_uop_lrs1,
                io_core_exe_0_req_bits_uop_lrs2,
                io_core_exe_0_req_bits_uop_lrs3,
  input         io_core_exe_0_req_bits_uop_ldst_val,
  input  [1:0]  io_core_exe_0_req_bits_uop_dst_rtype,
                io_core_exe_0_req_bits_uop_lrs1_rtype,
                io_core_exe_0_req_bits_uop_lrs2_rtype,
  input         io_core_exe_0_req_bits_uop_frs3_en,
                io_core_exe_0_req_bits_uop_fp_val,
                io_core_exe_0_req_bits_uop_fp_single,
                io_core_exe_0_req_bits_uop_xcpt_pf_if,
                io_core_exe_0_req_bits_uop_xcpt_ae_if,
                io_core_exe_0_req_bits_uop_xcpt_ma_if,
                io_core_exe_0_req_bits_uop_bp_debug_if,
                io_core_exe_0_req_bits_uop_bp_xcpt_if,
  input  [1:0]  io_core_exe_0_req_bits_uop_debug_fsrc,
                io_core_exe_0_req_bits_uop_debug_tsrc,
  input  [63:0] io_core_exe_0_req_bits_data,
  input  [39:0] io_core_exe_0_req_bits_addr,
  input         io_core_exe_0_req_bits_mxcpt_valid,
                io_core_exe_0_req_bits_sfence_valid,
                io_core_exe_0_req_bits_sfence_bits_rs1,
                io_core_exe_0_req_bits_sfence_bits_rs2,
  input  [38:0] io_core_exe_0_req_bits_sfence_bits_addr,
  output        io_core_exe_0_iresp_valid,
  output [6:0]  io_core_exe_0_iresp_bits_uop_rob_idx,
                io_core_exe_0_iresp_bits_uop_pdst,
  output        io_core_exe_0_iresp_bits_uop_is_amo,
                io_core_exe_0_iresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_iresp_bits_uop_dst_rtype,
  output [63:0] io_core_exe_0_iresp_bits_data,
  output        io_core_exe_0_fresp_valid,
  output [6:0]  io_core_exe_0_fresp_bits_uop_uopc,
  output [19:0] io_core_exe_0_fresp_bits_uop_br_mask,
  output [6:0]  io_core_exe_0_fresp_bits_uop_rob_idx,
  output [4:0]  io_core_exe_0_fresp_bits_uop_stq_idx,
  output [6:0]  io_core_exe_0_fresp_bits_uop_pdst,
  output [1:0]  io_core_exe_0_fresp_bits_uop_mem_size,
  output        io_core_exe_0_fresp_bits_uop_is_amo,
                io_core_exe_0_fresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_fresp_bits_uop_dst_rtype,
  output        io_core_exe_0_fresp_bits_uop_fp_val,
  output [64:0] io_core_exe_0_fresp_bits_data,
  input         io_core_exe_1_req_valid,
  input  [6:0]  io_core_exe_1_req_bits_uop_uopc,
  input  [31:0] io_core_exe_1_req_bits_uop_inst,
                io_core_exe_1_req_bits_uop_debug_inst,
  input         io_core_exe_1_req_bits_uop_is_rvc,
  input  [39:0] io_core_exe_1_req_bits_uop_debug_pc,
  input  [2:0]  io_core_exe_1_req_bits_uop_iq_type,
  input  [9:0]  io_core_exe_1_req_bits_uop_fu_code,
  input  [3:0]  io_core_exe_1_req_bits_uop_ctrl_br_type,
  input  [1:0]  io_core_exe_1_req_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_core_exe_1_req_bits_uop_ctrl_op2_sel,
                io_core_exe_1_req_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_core_exe_1_req_bits_uop_ctrl_op_fcn,
  input         io_core_exe_1_req_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_core_exe_1_req_bits_uop_ctrl_csr_cmd,
  input         io_core_exe_1_req_bits_uop_ctrl_is_load,
                io_core_exe_1_req_bits_uop_ctrl_is_sta,
                io_core_exe_1_req_bits_uop_ctrl_is_std,
  input  [1:0]  io_core_exe_1_req_bits_uop_iw_state,
  input         io_core_exe_1_req_bits_uop_is_br,
                io_core_exe_1_req_bits_uop_is_jalr,
                io_core_exe_1_req_bits_uop_is_jal,
                io_core_exe_1_req_bits_uop_is_sfb,
  input  [19:0] io_core_exe_1_req_bits_uop_br_mask,
  input  [4:0]  io_core_exe_1_req_bits_uop_br_tag,
  input  [5:0]  io_core_exe_1_req_bits_uop_ftq_idx,
  input         io_core_exe_1_req_bits_uop_edge_inst,
  input  [5:0]  io_core_exe_1_req_bits_uop_pc_lob,
  input         io_core_exe_1_req_bits_uop_taken,
  input  [19:0] io_core_exe_1_req_bits_uop_imm_packed,
  input  [11:0] io_core_exe_1_req_bits_uop_csr_addr,
  input  [6:0]  io_core_exe_1_req_bits_uop_rob_idx,
  input  [4:0]  io_core_exe_1_req_bits_uop_ldq_idx,
                io_core_exe_1_req_bits_uop_stq_idx,
  input  [1:0]  io_core_exe_1_req_bits_uop_rxq_idx,
  input  [6:0]  io_core_exe_1_req_bits_uop_pdst,
                io_core_exe_1_req_bits_uop_prs1,
                io_core_exe_1_req_bits_uop_prs2,
                io_core_exe_1_req_bits_uop_prs3,
  input  [5:0]  io_core_exe_1_req_bits_uop_ppred,
  input         io_core_exe_1_req_bits_uop_prs1_busy,
                io_core_exe_1_req_bits_uop_prs2_busy,
                io_core_exe_1_req_bits_uop_prs3_busy,
                io_core_exe_1_req_bits_uop_ppred_busy,
  input  [6:0]  io_core_exe_1_req_bits_uop_stale_pdst,
  input         io_core_exe_1_req_bits_uop_exception,
  input  [63:0] io_core_exe_1_req_bits_uop_exc_cause,
  input         io_core_exe_1_req_bits_uop_bypassable,
  input  [4:0]  io_core_exe_1_req_bits_uop_mem_cmd,
  input  [1:0]  io_core_exe_1_req_bits_uop_mem_size,
  input         io_core_exe_1_req_bits_uop_mem_signed,
                io_core_exe_1_req_bits_uop_is_fence,
                io_core_exe_1_req_bits_uop_is_fencei,
                io_core_exe_1_req_bits_uop_is_amo,
                io_core_exe_1_req_bits_uop_uses_ldq,
                io_core_exe_1_req_bits_uop_uses_stq,
                io_core_exe_1_req_bits_uop_is_sys_pc2epc,
                io_core_exe_1_req_bits_uop_is_unique,
                io_core_exe_1_req_bits_uop_flush_on_commit,
                io_core_exe_1_req_bits_uop_ldst_is_rs1,
  input  [5:0]  io_core_exe_1_req_bits_uop_ldst,
                io_core_exe_1_req_bits_uop_lrs1,
                io_core_exe_1_req_bits_uop_lrs2,
                io_core_exe_1_req_bits_uop_lrs3,
  input         io_core_exe_1_req_bits_uop_ldst_val,
  input  [1:0]  io_core_exe_1_req_bits_uop_dst_rtype,
                io_core_exe_1_req_bits_uop_lrs1_rtype,
                io_core_exe_1_req_bits_uop_lrs2_rtype,
  input         io_core_exe_1_req_bits_uop_frs3_en,
                io_core_exe_1_req_bits_uop_fp_val,
                io_core_exe_1_req_bits_uop_fp_single,
                io_core_exe_1_req_bits_uop_xcpt_pf_if,
                io_core_exe_1_req_bits_uop_xcpt_ae_if,
                io_core_exe_1_req_bits_uop_xcpt_ma_if,
                io_core_exe_1_req_bits_uop_bp_debug_if,
                io_core_exe_1_req_bits_uop_bp_xcpt_if,
  input  [1:0]  io_core_exe_1_req_bits_uop_debug_fsrc,
                io_core_exe_1_req_bits_uop_debug_tsrc,
  input  [63:0] io_core_exe_1_req_bits_data,
  input  [39:0] io_core_exe_1_req_bits_addr,
  input         io_core_exe_1_req_bits_mxcpt_valid,
                io_core_exe_1_req_bits_sfence_valid,
                io_core_exe_1_req_bits_sfence_bits_rs1,
                io_core_exe_1_req_bits_sfence_bits_rs2,
  input  [38:0] io_core_exe_1_req_bits_sfence_bits_addr,
  output        io_core_exe_1_iresp_valid,
  output [6:0]  io_core_exe_1_iresp_bits_uop_rob_idx,
                io_core_exe_1_iresp_bits_uop_pdst,
  output        io_core_exe_1_iresp_bits_uop_is_amo,
                io_core_exe_1_iresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_1_iresp_bits_uop_dst_rtype,
  output [63:0] io_core_exe_1_iresp_bits_data,
  output        io_core_exe_1_fresp_valid,
  output [6:0]  io_core_exe_1_fresp_bits_uop_uopc,
  output [19:0] io_core_exe_1_fresp_bits_uop_br_mask,
  output [6:0]  io_core_exe_1_fresp_bits_uop_rob_idx,
  output [4:0]  io_core_exe_1_fresp_bits_uop_stq_idx,
  output [6:0]  io_core_exe_1_fresp_bits_uop_pdst,
  output [1:0]  io_core_exe_1_fresp_bits_uop_mem_size,
  output        io_core_exe_1_fresp_bits_uop_is_amo,
                io_core_exe_1_fresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_1_fresp_bits_uop_dst_rtype,
  output        io_core_exe_1_fresp_bits_uop_fp_val,
  output [64:0] io_core_exe_1_fresp_bits_data,
  input         io_core_dis_uops_0_valid,
  input  [6:0]  io_core_dis_uops_0_bits_uopc,
  input  [31:0] io_core_dis_uops_0_bits_inst,
                io_core_dis_uops_0_bits_debug_inst,
  input         io_core_dis_uops_0_bits_is_rvc,
  input  [39:0] io_core_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_0_bits_iq_type,
  input  [9:0]  io_core_dis_uops_0_bits_fu_code,
  input  [3:0]  io_core_dis_uops_0_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_0_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_0_bits_ctrl_op2_sel,
                io_core_dis_uops_0_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_0_bits_ctrl_op_fcn,
  input         io_core_dis_uops_0_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_0_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_0_bits_ctrl_is_load,
                io_core_dis_uops_0_bits_ctrl_is_sta,
                io_core_dis_uops_0_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_0_bits_iw_state,
  input         io_core_dis_uops_0_bits_iw_p1_poisoned,
                io_core_dis_uops_0_bits_iw_p2_poisoned,
                io_core_dis_uops_0_bits_is_br,
                io_core_dis_uops_0_bits_is_jalr,
                io_core_dis_uops_0_bits_is_jal,
                io_core_dis_uops_0_bits_is_sfb,
  input  [19:0] io_core_dis_uops_0_bits_br_mask,
  input  [4:0]  io_core_dis_uops_0_bits_br_tag,
  input  [5:0]  io_core_dis_uops_0_bits_ftq_idx,
  input         io_core_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_0_bits_pc_lob,
  input         io_core_dis_uops_0_bits_taken,
  input  [19:0] io_core_dis_uops_0_bits_imm_packed,
  input  [11:0] io_core_dis_uops_0_bits_csr_addr,
  input  [6:0]  io_core_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_0_bits_ldq_idx,
                io_core_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_0_bits_pdst,
                io_core_dis_uops_0_bits_prs1,
                io_core_dis_uops_0_bits_prs2,
                io_core_dis_uops_0_bits_prs3,
  input         io_core_dis_uops_0_bits_prs1_busy,
                io_core_dis_uops_0_bits_prs2_busy,
                io_core_dis_uops_0_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_0_bits_stale_pdst,
  input         io_core_dis_uops_0_bits_exception,
  input  [63:0] io_core_dis_uops_0_bits_exc_cause,
  input         io_core_dis_uops_0_bits_bypassable,
  input  [4:0]  io_core_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_0_bits_mem_size,
  input         io_core_dis_uops_0_bits_mem_signed,
                io_core_dis_uops_0_bits_is_fence,
                io_core_dis_uops_0_bits_is_fencei,
                io_core_dis_uops_0_bits_is_amo,
                io_core_dis_uops_0_bits_uses_ldq,
                io_core_dis_uops_0_bits_uses_stq,
                io_core_dis_uops_0_bits_is_sys_pc2epc,
                io_core_dis_uops_0_bits_is_unique,
                io_core_dis_uops_0_bits_flush_on_commit,
                io_core_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_0_bits_ldst,
                io_core_dis_uops_0_bits_lrs1,
                io_core_dis_uops_0_bits_lrs2,
                io_core_dis_uops_0_bits_lrs3,
  input         io_core_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_0_bits_dst_rtype,
                io_core_dis_uops_0_bits_lrs1_rtype,
                io_core_dis_uops_0_bits_lrs2_rtype,
  input         io_core_dis_uops_0_bits_frs3_en,
                io_core_dis_uops_0_bits_fp_val,
                io_core_dis_uops_0_bits_fp_single,
                io_core_dis_uops_0_bits_xcpt_pf_if,
                io_core_dis_uops_0_bits_xcpt_ae_if,
                io_core_dis_uops_0_bits_xcpt_ma_if,
                io_core_dis_uops_0_bits_bp_debug_if,
                io_core_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_0_bits_debug_fsrc,
                io_core_dis_uops_0_bits_debug_tsrc,
  input         io_core_dis_uops_1_valid,
  input  [6:0]  io_core_dis_uops_1_bits_uopc,
  input  [31:0] io_core_dis_uops_1_bits_inst,
                io_core_dis_uops_1_bits_debug_inst,
  input         io_core_dis_uops_1_bits_is_rvc,
  input  [39:0] io_core_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_1_bits_iq_type,
  input  [9:0]  io_core_dis_uops_1_bits_fu_code,
  input  [3:0]  io_core_dis_uops_1_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_1_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_1_bits_ctrl_op2_sel,
                io_core_dis_uops_1_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_1_bits_ctrl_op_fcn,
  input         io_core_dis_uops_1_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_1_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_1_bits_ctrl_is_load,
                io_core_dis_uops_1_bits_ctrl_is_sta,
                io_core_dis_uops_1_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_1_bits_iw_state,
  input         io_core_dis_uops_1_bits_iw_p1_poisoned,
                io_core_dis_uops_1_bits_iw_p2_poisoned,
                io_core_dis_uops_1_bits_is_br,
                io_core_dis_uops_1_bits_is_jalr,
                io_core_dis_uops_1_bits_is_jal,
                io_core_dis_uops_1_bits_is_sfb,
  input  [19:0] io_core_dis_uops_1_bits_br_mask,
  input  [4:0]  io_core_dis_uops_1_bits_br_tag,
  input  [5:0]  io_core_dis_uops_1_bits_ftq_idx,
  input         io_core_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_1_bits_pc_lob,
  input         io_core_dis_uops_1_bits_taken,
  input  [19:0] io_core_dis_uops_1_bits_imm_packed,
  input  [11:0] io_core_dis_uops_1_bits_csr_addr,
  input  [6:0]  io_core_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_1_bits_ldq_idx,
                io_core_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_1_bits_pdst,
                io_core_dis_uops_1_bits_prs1,
                io_core_dis_uops_1_bits_prs2,
                io_core_dis_uops_1_bits_prs3,
  input         io_core_dis_uops_1_bits_prs1_busy,
                io_core_dis_uops_1_bits_prs2_busy,
                io_core_dis_uops_1_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_1_bits_stale_pdst,
  input         io_core_dis_uops_1_bits_exception,
  input  [63:0] io_core_dis_uops_1_bits_exc_cause,
  input         io_core_dis_uops_1_bits_bypassable,
  input  [4:0]  io_core_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_1_bits_mem_size,
  input         io_core_dis_uops_1_bits_mem_signed,
                io_core_dis_uops_1_bits_is_fence,
                io_core_dis_uops_1_bits_is_fencei,
                io_core_dis_uops_1_bits_is_amo,
                io_core_dis_uops_1_bits_uses_ldq,
                io_core_dis_uops_1_bits_uses_stq,
                io_core_dis_uops_1_bits_is_sys_pc2epc,
                io_core_dis_uops_1_bits_is_unique,
                io_core_dis_uops_1_bits_flush_on_commit,
                io_core_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_1_bits_ldst,
                io_core_dis_uops_1_bits_lrs1,
                io_core_dis_uops_1_bits_lrs2,
                io_core_dis_uops_1_bits_lrs3,
  input         io_core_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_1_bits_dst_rtype,
                io_core_dis_uops_1_bits_lrs1_rtype,
                io_core_dis_uops_1_bits_lrs2_rtype,
  input         io_core_dis_uops_1_bits_frs3_en,
                io_core_dis_uops_1_bits_fp_val,
                io_core_dis_uops_1_bits_fp_single,
                io_core_dis_uops_1_bits_xcpt_pf_if,
                io_core_dis_uops_1_bits_xcpt_ae_if,
                io_core_dis_uops_1_bits_xcpt_ma_if,
                io_core_dis_uops_1_bits_bp_debug_if,
                io_core_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_1_bits_debug_fsrc,
                io_core_dis_uops_1_bits_debug_tsrc,
  input         io_core_dis_uops_2_valid,
  input  [6:0]  io_core_dis_uops_2_bits_uopc,
  input  [31:0] io_core_dis_uops_2_bits_inst,
                io_core_dis_uops_2_bits_debug_inst,
  input         io_core_dis_uops_2_bits_is_rvc,
  input  [39:0] io_core_dis_uops_2_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_2_bits_iq_type,
  input  [9:0]  io_core_dis_uops_2_bits_fu_code,
  input  [3:0]  io_core_dis_uops_2_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_2_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_2_bits_ctrl_op2_sel,
                io_core_dis_uops_2_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_2_bits_ctrl_op_fcn,
  input         io_core_dis_uops_2_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_2_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_2_bits_ctrl_is_load,
                io_core_dis_uops_2_bits_ctrl_is_sta,
                io_core_dis_uops_2_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_2_bits_iw_state,
  input         io_core_dis_uops_2_bits_iw_p1_poisoned,
                io_core_dis_uops_2_bits_iw_p2_poisoned,
                io_core_dis_uops_2_bits_is_br,
                io_core_dis_uops_2_bits_is_jalr,
                io_core_dis_uops_2_bits_is_jal,
                io_core_dis_uops_2_bits_is_sfb,
  input  [19:0] io_core_dis_uops_2_bits_br_mask,
  input  [4:0]  io_core_dis_uops_2_bits_br_tag,
  input  [5:0]  io_core_dis_uops_2_bits_ftq_idx,
  input         io_core_dis_uops_2_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_2_bits_pc_lob,
  input         io_core_dis_uops_2_bits_taken,
  input  [19:0] io_core_dis_uops_2_bits_imm_packed,
  input  [11:0] io_core_dis_uops_2_bits_csr_addr,
  input  [6:0]  io_core_dis_uops_2_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_2_bits_ldq_idx,
                io_core_dis_uops_2_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_2_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_2_bits_pdst,
                io_core_dis_uops_2_bits_prs1,
                io_core_dis_uops_2_bits_prs2,
                io_core_dis_uops_2_bits_prs3,
  input         io_core_dis_uops_2_bits_prs1_busy,
                io_core_dis_uops_2_bits_prs2_busy,
                io_core_dis_uops_2_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_2_bits_stale_pdst,
  input         io_core_dis_uops_2_bits_exception,
  input  [63:0] io_core_dis_uops_2_bits_exc_cause,
  input         io_core_dis_uops_2_bits_bypassable,
  input  [4:0]  io_core_dis_uops_2_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_2_bits_mem_size,
  input         io_core_dis_uops_2_bits_mem_signed,
                io_core_dis_uops_2_bits_is_fence,
                io_core_dis_uops_2_bits_is_fencei,
                io_core_dis_uops_2_bits_is_amo,
                io_core_dis_uops_2_bits_uses_ldq,
                io_core_dis_uops_2_bits_uses_stq,
                io_core_dis_uops_2_bits_is_sys_pc2epc,
                io_core_dis_uops_2_bits_is_unique,
                io_core_dis_uops_2_bits_flush_on_commit,
                io_core_dis_uops_2_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_2_bits_ldst,
                io_core_dis_uops_2_bits_lrs1,
                io_core_dis_uops_2_bits_lrs2,
                io_core_dis_uops_2_bits_lrs3,
  input         io_core_dis_uops_2_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_2_bits_dst_rtype,
                io_core_dis_uops_2_bits_lrs1_rtype,
                io_core_dis_uops_2_bits_lrs2_rtype,
  input         io_core_dis_uops_2_bits_frs3_en,
                io_core_dis_uops_2_bits_fp_val,
                io_core_dis_uops_2_bits_fp_single,
                io_core_dis_uops_2_bits_xcpt_pf_if,
                io_core_dis_uops_2_bits_xcpt_ae_if,
                io_core_dis_uops_2_bits_xcpt_ma_if,
                io_core_dis_uops_2_bits_bp_debug_if,
                io_core_dis_uops_2_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_2_bits_debug_fsrc,
                io_core_dis_uops_2_bits_debug_tsrc,
  input         io_core_dis_uops_3_valid,
  input  [6:0]  io_core_dis_uops_3_bits_uopc,
  input  [31:0] io_core_dis_uops_3_bits_inst,
                io_core_dis_uops_3_bits_debug_inst,
  input         io_core_dis_uops_3_bits_is_rvc,
  input  [39:0] io_core_dis_uops_3_bits_debug_pc,
  input  [2:0]  io_core_dis_uops_3_bits_iq_type,
  input  [9:0]  io_core_dis_uops_3_bits_fu_code,
  input  [3:0]  io_core_dis_uops_3_bits_ctrl_br_type,
  input  [1:0]  io_core_dis_uops_3_bits_ctrl_op1_sel,
  input  [2:0]  io_core_dis_uops_3_bits_ctrl_op2_sel,
                io_core_dis_uops_3_bits_ctrl_imm_sel,
  input  [3:0]  io_core_dis_uops_3_bits_ctrl_op_fcn,
  input         io_core_dis_uops_3_bits_ctrl_fcn_dw,
  input  [2:0]  io_core_dis_uops_3_bits_ctrl_csr_cmd,
  input         io_core_dis_uops_3_bits_ctrl_is_load,
                io_core_dis_uops_3_bits_ctrl_is_sta,
                io_core_dis_uops_3_bits_ctrl_is_std,
  input  [1:0]  io_core_dis_uops_3_bits_iw_state,
  input         io_core_dis_uops_3_bits_iw_p1_poisoned,
                io_core_dis_uops_3_bits_iw_p2_poisoned,
                io_core_dis_uops_3_bits_is_br,
                io_core_dis_uops_3_bits_is_jalr,
                io_core_dis_uops_3_bits_is_jal,
                io_core_dis_uops_3_bits_is_sfb,
  input  [19:0] io_core_dis_uops_3_bits_br_mask,
  input  [4:0]  io_core_dis_uops_3_bits_br_tag,
  input  [5:0]  io_core_dis_uops_3_bits_ftq_idx,
  input         io_core_dis_uops_3_bits_edge_inst,
  input  [5:0]  io_core_dis_uops_3_bits_pc_lob,
  input         io_core_dis_uops_3_bits_taken,
  input  [19:0] io_core_dis_uops_3_bits_imm_packed,
  input  [11:0] io_core_dis_uops_3_bits_csr_addr,
  input  [6:0]  io_core_dis_uops_3_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_3_bits_ldq_idx,
                io_core_dis_uops_3_bits_stq_idx,
  input  [1:0]  io_core_dis_uops_3_bits_rxq_idx,
  input  [6:0]  io_core_dis_uops_3_bits_pdst,
                io_core_dis_uops_3_bits_prs1,
                io_core_dis_uops_3_bits_prs2,
                io_core_dis_uops_3_bits_prs3,
  input         io_core_dis_uops_3_bits_prs1_busy,
                io_core_dis_uops_3_bits_prs2_busy,
                io_core_dis_uops_3_bits_prs3_busy,
  input  [6:0]  io_core_dis_uops_3_bits_stale_pdst,
  input         io_core_dis_uops_3_bits_exception,
  input  [63:0] io_core_dis_uops_3_bits_exc_cause,
  input         io_core_dis_uops_3_bits_bypassable,
  input  [4:0]  io_core_dis_uops_3_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_3_bits_mem_size,
  input         io_core_dis_uops_3_bits_mem_signed,
                io_core_dis_uops_3_bits_is_fence,
                io_core_dis_uops_3_bits_is_fencei,
                io_core_dis_uops_3_bits_is_amo,
                io_core_dis_uops_3_bits_uses_ldq,
                io_core_dis_uops_3_bits_uses_stq,
                io_core_dis_uops_3_bits_is_sys_pc2epc,
                io_core_dis_uops_3_bits_is_unique,
                io_core_dis_uops_3_bits_flush_on_commit,
                io_core_dis_uops_3_bits_ldst_is_rs1,
  input  [5:0]  io_core_dis_uops_3_bits_ldst,
                io_core_dis_uops_3_bits_lrs1,
                io_core_dis_uops_3_bits_lrs2,
                io_core_dis_uops_3_bits_lrs3,
  input         io_core_dis_uops_3_bits_ldst_val,
  input  [1:0]  io_core_dis_uops_3_bits_dst_rtype,
                io_core_dis_uops_3_bits_lrs1_rtype,
                io_core_dis_uops_3_bits_lrs2_rtype,
  input         io_core_dis_uops_3_bits_frs3_en,
                io_core_dis_uops_3_bits_fp_val,
                io_core_dis_uops_3_bits_fp_single,
                io_core_dis_uops_3_bits_xcpt_pf_if,
                io_core_dis_uops_3_bits_xcpt_ae_if,
                io_core_dis_uops_3_bits_xcpt_ma_if,
                io_core_dis_uops_3_bits_bp_debug_if,
                io_core_dis_uops_3_bits_bp_xcpt_if,
  input  [1:0]  io_core_dis_uops_3_bits_debug_fsrc,
                io_core_dis_uops_3_bits_debug_tsrc,
  output [4:0]  io_core_dis_ldq_idx_0,
                io_core_dis_ldq_idx_1,
                io_core_dis_ldq_idx_2,
                io_core_dis_ldq_idx_3,
                io_core_dis_stq_idx_0,
                io_core_dis_stq_idx_1,
                io_core_dis_stq_idx_2,
                io_core_dis_stq_idx_3,
  output        io_core_ldq_full_0,
                io_core_ldq_full_1,
                io_core_ldq_full_2,
                io_core_ldq_full_3,
                io_core_stq_full_0,
                io_core_stq_full_1,
                io_core_stq_full_2,
                io_core_stq_full_3,
                io_core_fp_stdata_ready,
  input         io_core_fp_stdata_valid,
  input  [19:0] io_core_fp_stdata_bits_uop_br_mask,
  input  [6:0]  io_core_fp_stdata_bits_uop_rob_idx,
  input  [4:0]  io_core_fp_stdata_bits_uop_stq_idx,
  input  [63:0] io_core_fp_stdata_bits_data,
  input         io_core_commit_valids_0,
                io_core_commit_valids_1,
                io_core_commit_valids_2,
                io_core_commit_valids_3,
                io_core_commit_uops_0_uses_ldq,
                io_core_commit_uops_0_uses_stq,
                io_core_commit_uops_1_uses_ldq,
                io_core_commit_uops_1_uses_stq,
                io_core_commit_uops_2_uses_ldq,
                io_core_commit_uops_2_uses_stq,
                io_core_commit_uops_3_uses_ldq,
                io_core_commit_uops_3_uses_stq,
                io_core_commit_load_at_rob_head,
  output        io_core_clr_bsy_0_valid,
  output [6:0]  io_core_clr_bsy_0_bits,
  output        io_core_clr_bsy_1_valid,
  output [6:0]  io_core_clr_bsy_1_bits,
  output        io_core_clr_bsy_2_valid,
  output [6:0]  io_core_clr_bsy_2_bits,
  input         io_core_fence_dmem,
  output        io_core_spec_ld_wakeup_0_valid,
  output [6:0]  io_core_spec_ld_wakeup_0_bits,
  output        io_core_spec_ld_wakeup_1_valid,
  output [6:0]  io_core_spec_ld_wakeup_1_bits,
  output        io_core_ld_miss,
  input  [19:0] io_core_brupdate_b1_resolve_mask,
                io_core_brupdate_b1_mispredict_mask,
  input  [4:0]  io_core_brupdate_b2_uop_ldq_idx,
                io_core_brupdate_b2_uop_stq_idx,
  input         io_core_brupdate_b2_mispredict,
  input  [6:0]  io_core_rob_head_idx,
  input         io_core_exception,
  output        io_core_fencei_rdy,
                io_core_lxcpt_valid,
  output [19:0] io_core_lxcpt_bits_uop_br_mask,
  output [6:0]  io_core_lxcpt_bits_uop_rob_idx,
  output [4:0]  io_core_lxcpt_bits_cause,
  output [39:0] io_core_lxcpt_bits_badvaddr,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
                io_dmem_req_bits_0_valid,
  output [6:0]  io_dmem_req_bits_0_bits_uop_uopc,
  output [31:0] io_dmem_req_bits_0_bits_uop_inst,
                io_dmem_req_bits_0_bits_uop_debug_inst,
  output        io_dmem_req_bits_0_bits_uop_is_rvc,
  output [39:0] io_dmem_req_bits_0_bits_uop_debug_pc,
  output [2:0]  io_dmem_req_bits_0_bits_uop_iq_type,
  output [9:0]  io_dmem_req_bits_0_bits_uop_fu_code,
  output [3:0]  io_dmem_req_bits_0_bits_uop_ctrl_br_type,
  output [1:0]  io_dmem_req_bits_0_bits_uop_ctrl_op1_sel,
  output [2:0]  io_dmem_req_bits_0_bits_uop_ctrl_op2_sel,
                io_dmem_req_bits_0_bits_uop_ctrl_imm_sel,
  output [3:0]  io_dmem_req_bits_0_bits_uop_ctrl_op_fcn,
  output        io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd,
  output        io_dmem_req_bits_0_bits_uop_ctrl_is_load,
                io_dmem_req_bits_0_bits_uop_ctrl_is_sta,
                io_dmem_req_bits_0_bits_uop_ctrl_is_std,
  output [1:0]  io_dmem_req_bits_0_bits_uop_iw_state,
  output        io_dmem_req_bits_0_bits_uop_iw_p1_poisoned,
                io_dmem_req_bits_0_bits_uop_iw_p2_poisoned,
                io_dmem_req_bits_0_bits_uop_is_br,
                io_dmem_req_bits_0_bits_uop_is_jalr,
                io_dmem_req_bits_0_bits_uop_is_jal,
                io_dmem_req_bits_0_bits_uop_is_sfb,
  output [19:0] io_dmem_req_bits_0_bits_uop_br_mask,
  output [4:0]  io_dmem_req_bits_0_bits_uop_br_tag,
  output [5:0]  io_dmem_req_bits_0_bits_uop_ftq_idx,
  output        io_dmem_req_bits_0_bits_uop_edge_inst,
  output [5:0]  io_dmem_req_bits_0_bits_uop_pc_lob,
  output        io_dmem_req_bits_0_bits_uop_taken,
  output [19:0] io_dmem_req_bits_0_bits_uop_imm_packed,
  output [11:0] io_dmem_req_bits_0_bits_uop_csr_addr,
  output [6:0]  io_dmem_req_bits_0_bits_uop_rob_idx,
  output [4:0]  io_dmem_req_bits_0_bits_uop_ldq_idx,
                io_dmem_req_bits_0_bits_uop_stq_idx,
  output [1:0]  io_dmem_req_bits_0_bits_uop_rxq_idx,
  output [6:0]  io_dmem_req_bits_0_bits_uop_pdst,
                io_dmem_req_bits_0_bits_uop_prs1,
                io_dmem_req_bits_0_bits_uop_prs2,
                io_dmem_req_bits_0_bits_uop_prs3,
  output [5:0]  io_dmem_req_bits_0_bits_uop_ppred,
  output        io_dmem_req_bits_0_bits_uop_prs1_busy,
                io_dmem_req_bits_0_bits_uop_prs2_busy,
                io_dmem_req_bits_0_bits_uop_prs3_busy,
                io_dmem_req_bits_0_bits_uop_ppred_busy,
  output [6:0]  io_dmem_req_bits_0_bits_uop_stale_pdst,
  output        io_dmem_req_bits_0_bits_uop_exception,
  output [63:0] io_dmem_req_bits_0_bits_uop_exc_cause,
  output        io_dmem_req_bits_0_bits_uop_bypassable,
  output [4:0]  io_dmem_req_bits_0_bits_uop_mem_cmd,
  output [1:0]  io_dmem_req_bits_0_bits_uop_mem_size,
  output        io_dmem_req_bits_0_bits_uop_mem_signed,
                io_dmem_req_bits_0_bits_uop_is_fence,
                io_dmem_req_bits_0_bits_uop_is_fencei,
                io_dmem_req_bits_0_bits_uop_is_amo,
                io_dmem_req_bits_0_bits_uop_uses_ldq,
                io_dmem_req_bits_0_bits_uop_uses_stq,
                io_dmem_req_bits_0_bits_uop_is_sys_pc2epc,
                io_dmem_req_bits_0_bits_uop_is_unique,
                io_dmem_req_bits_0_bits_uop_flush_on_commit,
                io_dmem_req_bits_0_bits_uop_ldst_is_rs1,
  output [5:0]  io_dmem_req_bits_0_bits_uop_ldst,
                io_dmem_req_bits_0_bits_uop_lrs1,
                io_dmem_req_bits_0_bits_uop_lrs2,
                io_dmem_req_bits_0_bits_uop_lrs3,
  output        io_dmem_req_bits_0_bits_uop_ldst_val,
  output [1:0]  io_dmem_req_bits_0_bits_uop_dst_rtype,
                io_dmem_req_bits_0_bits_uop_lrs1_rtype,
                io_dmem_req_bits_0_bits_uop_lrs2_rtype,
  output        io_dmem_req_bits_0_bits_uop_frs3_en,
                io_dmem_req_bits_0_bits_uop_fp_val,
                io_dmem_req_bits_0_bits_uop_fp_single,
                io_dmem_req_bits_0_bits_uop_xcpt_pf_if,
                io_dmem_req_bits_0_bits_uop_xcpt_ae_if,
                io_dmem_req_bits_0_bits_uop_xcpt_ma_if,
                io_dmem_req_bits_0_bits_uop_bp_debug_if,
                io_dmem_req_bits_0_bits_uop_bp_xcpt_if,
  output [1:0]  io_dmem_req_bits_0_bits_uop_debug_fsrc,
                io_dmem_req_bits_0_bits_uop_debug_tsrc,
  output [39:0] io_dmem_req_bits_0_bits_addr,
  output [63:0] io_dmem_req_bits_0_bits_data,
  output        io_dmem_req_bits_0_bits_is_hella,
                io_dmem_req_bits_1_valid,
  output [6:0]  io_dmem_req_bits_1_bits_uop_uopc,
  output [31:0] io_dmem_req_bits_1_bits_uop_inst,
                io_dmem_req_bits_1_bits_uop_debug_inst,
  output        io_dmem_req_bits_1_bits_uop_is_rvc,
  output [39:0] io_dmem_req_bits_1_bits_uop_debug_pc,
  output [2:0]  io_dmem_req_bits_1_bits_uop_iq_type,
  output [9:0]  io_dmem_req_bits_1_bits_uop_fu_code,
  output [3:0]  io_dmem_req_bits_1_bits_uop_ctrl_br_type,
  output [1:0]  io_dmem_req_bits_1_bits_uop_ctrl_op1_sel,
  output [2:0]  io_dmem_req_bits_1_bits_uop_ctrl_op2_sel,
                io_dmem_req_bits_1_bits_uop_ctrl_imm_sel,
  output [3:0]  io_dmem_req_bits_1_bits_uop_ctrl_op_fcn,
  output        io_dmem_req_bits_1_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_dmem_req_bits_1_bits_uop_ctrl_csr_cmd,
  output        io_dmem_req_bits_1_bits_uop_ctrl_is_load,
                io_dmem_req_bits_1_bits_uop_ctrl_is_sta,
                io_dmem_req_bits_1_bits_uop_ctrl_is_std,
  output [1:0]  io_dmem_req_bits_1_bits_uop_iw_state,
  output        io_dmem_req_bits_1_bits_uop_iw_p1_poisoned,
                io_dmem_req_bits_1_bits_uop_iw_p2_poisoned,
                io_dmem_req_bits_1_bits_uop_is_br,
                io_dmem_req_bits_1_bits_uop_is_jalr,
                io_dmem_req_bits_1_bits_uop_is_jal,
                io_dmem_req_bits_1_bits_uop_is_sfb,
  output [19:0] io_dmem_req_bits_1_bits_uop_br_mask,
  output [4:0]  io_dmem_req_bits_1_bits_uop_br_tag,
  output [5:0]  io_dmem_req_bits_1_bits_uop_ftq_idx,
  output        io_dmem_req_bits_1_bits_uop_edge_inst,
  output [5:0]  io_dmem_req_bits_1_bits_uop_pc_lob,
  output        io_dmem_req_bits_1_bits_uop_taken,
  output [19:0] io_dmem_req_bits_1_bits_uop_imm_packed,
  output [11:0] io_dmem_req_bits_1_bits_uop_csr_addr,
  output [6:0]  io_dmem_req_bits_1_bits_uop_rob_idx,
  output [4:0]  io_dmem_req_bits_1_bits_uop_ldq_idx,
                io_dmem_req_bits_1_bits_uop_stq_idx,
  output [1:0]  io_dmem_req_bits_1_bits_uop_rxq_idx,
  output [6:0]  io_dmem_req_bits_1_bits_uop_pdst,
                io_dmem_req_bits_1_bits_uop_prs1,
                io_dmem_req_bits_1_bits_uop_prs2,
                io_dmem_req_bits_1_bits_uop_prs3,
  output [5:0]  io_dmem_req_bits_1_bits_uop_ppred,
  output        io_dmem_req_bits_1_bits_uop_prs1_busy,
                io_dmem_req_bits_1_bits_uop_prs2_busy,
                io_dmem_req_bits_1_bits_uop_prs3_busy,
                io_dmem_req_bits_1_bits_uop_ppred_busy,
  output [6:0]  io_dmem_req_bits_1_bits_uop_stale_pdst,
  output        io_dmem_req_bits_1_bits_uop_exception,
  output [63:0] io_dmem_req_bits_1_bits_uop_exc_cause,
  output        io_dmem_req_bits_1_bits_uop_bypassable,
  output [4:0]  io_dmem_req_bits_1_bits_uop_mem_cmd,
  output [1:0]  io_dmem_req_bits_1_bits_uop_mem_size,
  output        io_dmem_req_bits_1_bits_uop_mem_signed,
                io_dmem_req_bits_1_bits_uop_is_fence,
                io_dmem_req_bits_1_bits_uop_is_fencei,
                io_dmem_req_bits_1_bits_uop_is_amo,
                io_dmem_req_bits_1_bits_uop_uses_ldq,
                io_dmem_req_bits_1_bits_uop_uses_stq,
                io_dmem_req_bits_1_bits_uop_is_sys_pc2epc,
                io_dmem_req_bits_1_bits_uop_is_unique,
                io_dmem_req_bits_1_bits_uop_flush_on_commit,
                io_dmem_req_bits_1_bits_uop_ldst_is_rs1,
  output [5:0]  io_dmem_req_bits_1_bits_uop_ldst,
                io_dmem_req_bits_1_bits_uop_lrs1,
                io_dmem_req_bits_1_bits_uop_lrs2,
                io_dmem_req_bits_1_bits_uop_lrs3,
  output        io_dmem_req_bits_1_bits_uop_ldst_val,
  output [1:0]  io_dmem_req_bits_1_bits_uop_dst_rtype,
                io_dmem_req_bits_1_bits_uop_lrs1_rtype,
                io_dmem_req_bits_1_bits_uop_lrs2_rtype,
  output        io_dmem_req_bits_1_bits_uop_frs3_en,
                io_dmem_req_bits_1_bits_uop_fp_val,
                io_dmem_req_bits_1_bits_uop_fp_single,
                io_dmem_req_bits_1_bits_uop_xcpt_pf_if,
                io_dmem_req_bits_1_bits_uop_xcpt_ae_if,
                io_dmem_req_bits_1_bits_uop_xcpt_ma_if,
                io_dmem_req_bits_1_bits_uop_bp_debug_if,
                io_dmem_req_bits_1_bits_uop_bp_xcpt_if,
  output [1:0]  io_dmem_req_bits_1_bits_uop_debug_fsrc,
                io_dmem_req_bits_1_bits_uop_debug_tsrc,
  output [39:0] io_dmem_req_bits_1_bits_addr,
  output [63:0] io_dmem_req_bits_1_bits_data,
  output        io_dmem_req_bits_1_bits_is_hella,
                io_dmem_s1_kill_0,
                io_dmem_s1_kill_1,
  input         io_dmem_resp_0_valid,
  input  [4:0]  io_dmem_resp_0_bits_uop_ldq_idx,
                io_dmem_resp_0_bits_uop_stq_idx,
  input         io_dmem_resp_0_bits_uop_is_amo,
                io_dmem_resp_0_bits_uop_uses_ldq,
                io_dmem_resp_0_bits_uop_uses_stq,
  input  [63:0] io_dmem_resp_0_bits_data,
  input         io_dmem_resp_0_bits_is_hella,
                io_dmem_resp_1_valid,
  input  [4:0]  io_dmem_resp_1_bits_uop_ldq_idx,
                io_dmem_resp_1_bits_uop_stq_idx,
  input         io_dmem_resp_1_bits_uop_is_amo,
                io_dmem_resp_1_bits_uop_uses_ldq,
                io_dmem_resp_1_bits_uop_uses_stq,
  input  [63:0] io_dmem_resp_1_bits_data,
  input         io_dmem_resp_1_bits_is_hella,
                io_dmem_nack_0_valid,
  input  [4:0]  io_dmem_nack_0_bits_uop_ldq_idx,
                io_dmem_nack_0_bits_uop_stq_idx,
  input         io_dmem_nack_0_bits_uop_uses_ldq,
                io_dmem_nack_0_bits_uop_uses_stq,
                io_dmem_nack_0_bits_is_hella,
                io_dmem_nack_1_valid,
  input  [4:0]  io_dmem_nack_1_bits_uop_ldq_idx,
                io_dmem_nack_1_bits_uop_stq_idx,
  input         io_dmem_nack_1_bits_uop_uses_ldq,
                io_dmem_nack_1_bits_uop_uses_stq,
                io_dmem_nack_1_bits_is_hella,
  output [19:0] io_dmem_brupdate_b1_resolve_mask,
                io_dmem_brupdate_b1_mispredict_mask,
  output        io_dmem_exception,
                io_dmem_release_ready,
  input         io_dmem_release_valid,
  input  [32:0] io_dmem_release_bits_address,
  output        io_dmem_force_order,
  input         io_dmem_ordered,
  output        io_hellacache_req_ready,
  input         io_hellacache_req_valid,
  input  [39:0] io_hellacache_req_bits_addr,
  input         io_hellacache_s1_kill,
  output        io_hellacache_s2_nack,
                io_hellacache_resp_valid,
  output [63:0] io_hellacache_resp_bits_data,
  output        io_hellacache_s2_xcpt_ae_ld
);

  wire        _GEN;
  wire        _GEN_0;
  wire        store_needs_order;
  wire        nacking_loads_31;
  wire        nacking_loads_30;
  wire        nacking_loads_29;
  wire        nacking_loads_28;
  wire        nacking_loads_27;
  wire        nacking_loads_26;
  wire        nacking_loads_25;
  wire        nacking_loads_24;
  wire        nacking_loads_23;
  wire        nacking_loads_22;
  wire        nacking_loads_21;
  wire        nacking_loads_20;
  wire        nacking_loads_19;
  wire        nacking_loads_18;
  wire        nacking_loads_17;
  wire        nacking_loads_16;
  wire        nacking_loads_15;
  wire        nacking_loads_14;
  wire        nacking_loads_13;
  wire        nacking_loads_12;
  wire        nacking_loads_11;
  wire        nacking_loads_10;
  wire        nacking_loads_9;
  wire        nacking_loads_8;
  wire        nacking_loads_7;
  wire        nacking_loads_6;
  wire        nacking_loads_5;
  wire        nacking_loads_4;
  wire        nacking_loads_3;
  wire        nacking_loads_2;
  wire        nacking_loads_1;
  wire        nacking_loads_0;
  wire        dmem_req_1_valid;
  wire        dmem_req_0_valid;
  wire        _GEN_1;
  wire        _GEN_2;
  wire        mem_xcpt_valid;
  wire        _will_fire_store_commit_1_T_2;
  wire        _will_fire_store_commit_0_T_2;
  wire [4:0]  _forwarding_age_logic_1_io_forwarding_idx;
  wire [4:0]  _forwarding_age_logic_0_io_forwarding_idx;
  wire        _dtlb_io_miss_rdy;
  wire        _dtlb_io_resp_0_miss;
  wire [32:0] _dtlb_io_resp_0_paddr;
  wire        _dtlb_io_resp_0_pf_ld;
  wire        _dtlb_io_resp_0_pf_st;
  wire        _dtlb_io_resp_0_ae_ld;
  wire        _dtlb_io_resp_0_ae_st;
  wire        _dtlb_io_resp_0_cacheable;
  wire        _dtlb_io_resp_1_miss;
  wire [32:0] _dtlb_io_resp_1_paddr;
  wire        _dtlb_io_resp_1_pf_ld;
  wire        _dtlb_io_resp_1_pf_st;
  wire        _dtlb_io_resp_1_ae_ld;
  wire        _dtlb_io_resp_1_ae_st;
  wire        _dtlb_io_resp_1_ma_ld;
  wire        _dtlb_io_resp_1_ma_st;
  wire        _dtlb_io_resp_1_cacheable;
  wire        will_fire_release_0_will_fire = 1'h0;
  wire        will_fire_hella_incoming_0_will_fire = 1'h0;
  wire        will_fire_hella_wakeup_0_will_fire = 1'h0;
  wire        will_fire_load_retry_0_will_fire = 1'h0;
  wire        will_fire_sta_retry_0_will_fire = 1'h0;
  wire        will_fire_load_wakeup_0_will_fire = 1'h0;
  wire        will_fire_store_commit_1_will_fire = 1'h0;
  reg         ldq_0_valid;
  reg  [6:0]  ldq_0_bits_uop_uopc;
  reg  [31:0] ldq_0_bits_uop_inst;
  reg  [31:0] ldq_0_bits_uop_debug_inst;
  reg         ldq_0_bits_uop_is_rvc;
  reg  [39:0] ldq_0_bits_uop_debug_pc;
  reg  [2:0]  ldq_0_bits_uop_iq_type;
  reg  [9:0]  ldq_0_bits_uop_fu_code;
  reg  [3:0]  ldq_0_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_0_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_0_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_0_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_0_bits_uop_ctrl_op_fcn;
  reg         ldq_0_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_0_bits_uop_ctrl_csr_cmd;
  reg         ldq_0_bits_uop_ctrl_is_load;
  reg         ldq_0_bits_uop_ctrl_is_sta;
  reg         ldq_0_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_0_bits_uop_iw_state;
  reg         ldq_0_bits_uop_iw_p1_poisoned;
  reg         ldq_0_bits_uop_iw_p2_poisoned;
  reg         ldq_0_bits_uop_is_br;
  reg         ldq_0_bits_uop_is_jalr;
  reg         ldq_0_bits_uop_is_jal;
  reg         ldq_0_bits_uop_is_sfb;
  reg  [19:0] ldq_0_bits_uop_br_mask;
  reg  [4:0]  ldq_0_bits_uop_br_tag;
  reg  [5:0]  ldq_0_bits_uop_ftq_idx;
  reg         ldq_0_bits_uop_edge_inst;
  reg  [5:0]  ldq_0_bits_uop_pc_lob;
  reg         ldq_0_bits_uop_taken;
  reg  [19:0] ldq_0_bits_uop_imm_packed;
  reg  [11:0] ldq_0_bits_uop_csr_addr;
  reg  [6:0]  ldq_0_bits_uop_rob_idx;
  reg  [4:0]  ldq_0_bits_uop_ldq_idx;
  reg  [4:0]  ldq_0_bits_uop_stq_idx;
  reg  [1:0]  ldq_0_bits_uop_rxq_idx;
  reg  [6:0]  ldq_0_bits_uop_pdst;
  reg  [6:0]  ldq_0_bits_uop_prs1;
  reg  [6:0]  ldq_0_bits_uop_prs2;
  reg  [6:0]  ldq_0_bits_uop_prs3;
  reg         ldq_0_bits_uop_prs1_busy;
  reg         ldq_0_bits_uop_prs2_busy;
  reg         ldq_0_bits_uop_prs3_busy;
  reg  [6:0]  ldq_0_bits_uop_stale_pdst;
  reg         ldq_0_bits_uop_exception;
  reg  [63:0] ldq_0_bits_uop_exc_cause;
  reg         ldq_0_bits_uop_bypassable;
  reg  [4:0]  ldq_0_bits_uop_mem_cmd;
  reg  [1:0]  ldq_0_bits_uop_mem_size;
  reg         ldq_0_bits_uop_mem_signed;
  reg         ldq_0_bits_uop_is_fence;
  reg         ldq_0_bits_uop_is_fencei;
  reg         ldq_0_bits_uop_is_amo;
  reg         ldq_0_bits_uop_uses_ldq;
  reg         ldq_0_bits_uop_uses_stq;
  reg         ldq_0_bits_uop_is_sys_pc2epc;
  reg         ldq_0_bits_uop_is_unique;
  reg         ldq_0_bits_uop_flush_on_commit;
  reg         ldq_0_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_0_bits_uop_ldst;
  reg  [5:0]  ldq_0_bits_uop_lrs1;
  reg  [5:0]  ldq_0_bits_uop_lrs2;
  reg  [5:0]  ldq_0_bits_uop_lrs3;
  reg         ldq_0_bits_uop_ldst_val;
  reg  [1:0]  ldq_0_bits_uop_dst_rtype;
  reg  [1:0]  ldq_0_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_0_bits_uop_lrs2_rtype;
  reg         ldq_0_bits_uop_frs3_en;
  reg         ldq_0_bits_uop_fp_val;
  reg         ldq_0_bits_uop_fp_single;
  reg         ldq_0_bits_uop_xcpt_pf_if;
  reg         ldq_0_bits_uop_xcpt_ae_if;
  reg         ldq_0_bits_uop_xcpt_ma_if;
  reg         ldq_0_bits_uop_bp_debug_if;
  reg         ldq_0_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_0_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_0_bits_uop_debug_tsrc;
  reg         ldq_0_bits_addr_valid;
  reg  [39:0] ldq_0_bits_addr_bits;
  reg         ldq_0_bits_addr_is_virtual;
  reg         ldq_0_bits_addr_is_uncacheable;
  reg         ldq_0_bits_executed;
  reg         ldq_0_bits_succeeded;
  reg         ldq_0_bits_order_fail;
  reg         ldq_0_bits_observed;
  reg  [31:0] ldq_0_bits_st_dep_mask;
  reg  [4:0]  ldq_0_bits_youngest_stq_idx;
  reg         ldq_0_bits_forward_std_val;
  reg  [4:0]  ldq_0_bits_forward_stq_idx;
  reg         ldq_1_valid;
  reg  [6:0]  ldq_1_bits_uop_uopc;
  reg  [31:0] ldq_1_bits_uop_inst;
  reg  [31:0] ldq_1_bits_uop_debug_inst;
  reg         ldq_1_bits_uop_is_rvc;
  reg  [39:0] ldq_1_bits_uop_debug_pc;
  reg  [2:0]  ldq_1_bits_uop_iq_type;
  reg  [9:0]  ldq_1_bits_uop_fu_code;
  reg  [3:0]  ldq_1_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_1_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_1_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_1_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_1_bits_uop_ctrl_op_fcn;
  reg         ldq_1_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_1_bits_uop_ctrl_csr_cmd;
  reg         ldq_1_bits_uop_ctrl_is_load;
  reg         ldq_1_bits_uop_ctrl_is_sta;
  reg         ldq_1_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_1_bits_uop_iw_state;
  reg         ldq_1_bits_uop_iw_p1_poisoned;
  reg         ldq_1_bits_uop_iw_p2_poisoned;
  reg         ldq_1_bits_uop_is_br;
  reg         ldq_1_bits_uop_is_jalr;
  reg         ldq_1_bits_uop_is_jal;
  reg         ldq_1_bits_uop_is_sfb;
  reg  [19:0] ldq_1_bits_uop_br_mask;
  reg  [4:0]  ldq_1_bits_uop_br_tag;
  reg  [5:0]  ldq_1_bits_uop_ftq_idx;
  reg         ldq_1_bits_uop_edge_inst;
  reg  [5:0]  ldq_1_bits_uop_pc_lob;
  reg         ldq_1_bits_uop_taken;
  reg  [19:0] ldq_1_bits_uop_imm_packed;
  reg  [11:0] ldq_1_bits_uop_csr_addr;
  reg  [6:0]  ldq_1_bits_uop_rob_idx;
  reg  [4:0]  ldq_1_bits_uop_ldq_idx;
  reg  [4:0]  ldq_1_bits_uop_stq_idx;
  reg  [1:0]  ldq_1_bits_uop_rxq_idx;
  reg  [6:0]  ldq_1_bits_uop_pdst;
  reg  [6:0]  ldq_1_bits_uop_prs1;
  reg  [6:0]  ldq_1_bits_uop_prs2;
  reg  [6:0]  ldq_1_bits_uop_prs3;
  reg         ldq_1_bits_uop_prs1_busy;
  reg         ldq_1_bits_uop_prs2_busy;
  reg         ldq_1_bits_uop_prs3_busy;
  reg  [6:0]  ldq_1_bits_uop_stale_pdst;
  reg         ldq_1_bits_uop_exception;
  reg  [63:0] ldq_1_bits_uop_exc_cause;
  reg         ldq_1_bits_uop_bypassable;
  reg  [4:0]  ldq_1_bits_uop_mem_cmd;
  reg  [1:0]  ldq_1_bits_uop_mem_size;
  reg         ldq_1_bits_uop_mem_signed;
  reg         ldq_1_bits_uop_is_fence;
  reg         ldq_1_bits_uop_is_fencei;
  reg         ldq_1_bits_uop_is_amo;
  reg         ldq_1_bits_uop_uses_ldq;
  reg         ldq_1_bits_uop_uses_stq;
  reg         ldq_1_bits_uop_is_sys_pc2epc;
  reg         ldq_1_bits_uop_is_unique;
  reg         ldq_1_bits_uop_flush_on_commit;
  reg         ldq_1_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_1_bits_uop_ldst;
  reg  [5:0]  ldq_1_bits_uop_lrs1;
  reg  [5:0]  ldq_1_bits_uop_lrs2;
  reg  [5:0]  ldq_1_bits_uop_lrs3;
  reg         ldq_1_bits_uop_ldst_val;
  reg  [1:0]  ldq_1_bits_uop_dst_rtype;
  reg  [1:0]  ldq_1_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_1_bits_uop_lrs2_rtype;
  reg         ldq_1_bits_uop_frs3_en;
  reg         ldq_1_bits_uop_fp_val;
  reg         ldq_1_bits_uop_fp_single;
  reg         ldq_1_bits_uop_xcpt_pf_if;
  reg         ldq_1_bits_uop_xcpt_ae_if;
  reg         ldq_1_bits_uop_xcpt_ma_if;
  reg         ldq_1_bits_uop_bp_debug_if;
  reg         ldq_1_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_1_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_1_bits_uop_debug_tsrc;
  reg         ldq_1_bits_addr_valid;
  reg  [39:0] ldq_1_bits_addr_bits;
  reg         ldq_1_bits_addr_is_virtual;
  reg         ldq_1_bits_addr_is_uncacheable;
  reg         ldq_1_bits_executed;
  reg         ldq_1_bits_succeeded;
  reg         ldq_1_bits_order_fail;
  reg         ldq_1_bits_observed;
  reg  [31:0] ldq_1_bits_st_dep_mask;
  reg  [4:0]  ldq_1_bits_youngest_stq_idx;
  reg         ldq_1_bits_forward_std_val;
  reg  [4:0]  ldq_1_bits_forward_stq_idx;
  reg         ldq_2_valid;
  reg  [6:0]  ldq_2_bits_uop_uopc;
  reg  [31:0] ldq_2_bits_uop_inst;
  reg  [31:0] ldq_2_bits_uop_debug_inst;
  reg         ldq_2_bits_uop_is_rvc;
  reg  [39:0] ldq_2_bits_uop_debug_pc;
  reg  [2:0]  ldq_2_bits_uop_iq_type;
  reg  [9:0]  ldq_2_bits_uop_fu_code;
  reg  [3:0]  ldq_2_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_2_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_2_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_2_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_2_bits_uop_ctrl_op_fcn;
  reg         ldq_2_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_2_bits_uop_ctrl_csr_cmd;
  reg         ldq_2_bits_uop_ctrl_is_load;
  reg         ldq_2_bits_uop_ctrl_is_sta;
  reg         ldq_2_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_2_bits_uop_iw_state;
  reg         ldq_2_bits_uop_iw_p1_poisoned;
  reg         ldq_2_bits_uop_iw_p2_poisoned;
  reg         ldq_2_bits_uop_is_br;
  reg         ldq_2_bits_uop_is_jalr;
  reg         ldq_2_bits_uop_is_jal;
  reg         ldq_2_bits_uop_is_sfb;
  reg  [19:0] ldq_2_bits_uop_br_mask;
  reg  [4:0]  ldq_2_bits_uop_br_tag;
  reg  [5:0]  ldq_2_bits_uop_ftq_idx;
  reg         ldq_2_bits_uop_edge_inst;
  reg  [5:0]  ldq_2_bits_uop_pc_lob;
  reg         ldq_2_bits_uop_taken;
  reg  [19:0] ldq_2_bits_uop_imm_packed;
  reg  [11:0] ldq_2_bits_uop_csr_addr;
  reg  [6:0]  ldq_2_bits_uop_rob_idx;
  reg  [4:0]  ldq_2_bits_uop_ldq_idx;
  reg  [4:0]  ldq_2_bits_uop_stq_idx;
  reg  [1:0]  ldq_2_bits_uop_rxq_idx;
  reg  [6:0]  ldq_2_bits_uop_pdst;
  reg  [6:0]  ldq_2_bits_uop_prs1;
  reg  [6:0]  ldq_2_bits_uop_prs2;
  reg  [6:0]  ldq_2_bits_uop_prs3;
  reg         ldq_2_bits_uop_prs1_busy;
  reg         ldq_2_bits_uop_prs2_busy;
  reg         ldq_2_bits_uop_prs3_busy;
  reg  [6:0]  ldq_2_bits_uop_stale_pdst;
  reg         ldq_2_bits_uop_exception;
  reg  [63:0] ldq_2_bits_uop_exc_cause;
  reg         ldq_2_bits_uop_bypassable;
  reg  [4:0]  ldq_2_bits_uop_mem_cmd;
  reg  [1:0]  ldq_2_bits_uop_mem_size;
  reg         ldq_2_bits_uop_mem_signed;
  reg         ldq_2_bits_uop_is_fence;
  reg         ldq_2_bits_uop_is_fencei;
  reg         ldq_2_bits_uop_is_amo;
  reg         ldq_2_bits_uop_uses_ldq;
  reg         ldq_2_bits_uop_uses_stq;
  reg         ldq_2_bits_uop_is_sys_pc2epc;
  reg         ldq_2_bits_uop_is_unique;
  reg         ldq_2_bits_uop_flush_on_commit;
  reg         ldq_2_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_2_bits_uop_ldst;
  reg  [5:0]  ldq_2_bits_uop_lrs1;
  reg  [5:0]  ldq_2_bits_uop_lrs2;
  reg  [5:0]  ldq_2_bits_uop_lrs3;
  reg         ldq_2_bits_uop_ldst_val;
  reg  [1:0]  ldq_2_bits_uop_dst_rtype;
  reg  [1:0]  ldq_2_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_2_bits_uop_lrs2_rtype;
  reg         ldq_2_bits_uop_frs3_en;
  reg         ldq_2_bits_uop_fp_val;
  reg         ldq_2_bits_uop_fp_single;
  reg         ldq_2_bits_uop_xcpt_pf_if;
  reg         ldq_2_bits_uop_xcpt_ae_if;
  reg         ldq_2_bits_uop_xcpt_ma_if;
  reg         ldq_2_bits_uop_bp_debug_if;
  reg         ldq_2_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_2_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_2_bits_uop_debug_tsrc;
  reg         ldq_2_bits_addr_valid;
  reg  [39:0] ldq_2_bits_addr_bits;
  reg         ldq_2_bits_addr_is_virtual;
  reg         ldq_2_bits_addr_is_uncacheable;
  reg         ldq_2_bits_executed;
  reg         ldq_2_bits_succeeded;
  reg         ldq_2_bits_order_fail;
  reg         ldq_2_bits_observed;
  reg  [31:0] ldq_2_bits_st_dep_mask;
  reg  [4:0]  ldq_2_bits_youngest_stq_idx;
  reg         ldq_2_bits_forward_std_val;
  reg  [4:0]  ldq_2_bits_forward_stq_idx;
  reg         ldq_3_valid;
  reg  [6:0]  ldq_3_bits_uop_uopc;
  reg  [31:0] ldq_3_bits_uop_inst;
  reg  [31:0] ldq_3_bits_uop_debug_inst;
  reg         ldq_3_bits_uop_is_rvc;
  reg  [39:0] ldq_3_bits_uop_debug_pc;
  reg  [2:0]  ldq_3_bits_uop_iq_type;
  reg  [9:0]  ldq_3_bits_uop_fu_code;
  reg  [3:0]  ldq_3_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_3_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_3_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_3_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_3_bits_uop_ctrl_op_fcn;
  reg         ldq_3_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_3_bits_uop_ctrl_csr_cmd;
  reg         ldq_3_bits_uop_ctrl_is_load;
  reg         ldq_3_bits_uop_ctrl_is_sta;
  reg         ldq_3_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_3_bits_uop_iw_state;
  reg         ldq_3_bits_uop_iw_p1_poisoned;
  reg         ldq_3_bits_uop_iw_p2_poisoned;
  reg         ldq_3_bits_uop_is_br;
  reg         ldq_3_bits_uop_is_jalr;
  reg         ldq_3_bits_uop_is_jal;
  reg         ldq_3_bits_uop_is_sfb;
  reg  [19:0] ldq_3_bits_uop_br_mask;
  reg  [4:0]  ldq_3_bits_uop_br_tag;
  reg  [5:0]  ldq_3_bits_uop_ftq_idx;
  reg         ldq_3_bits_uop_edge_inst;
  reg  [5:0]  ldq_3_bits_uop_pc_lob;
  reg         ldq_3_bits_uop_taken;
  reg  [19:0] ldq_3_bits_uop_imm_packed;
  reg  [11:0] ldq_3_bits_uop_csr_addr;
  reg  [6:0]  ldq_3_bits_uop_rob_idx;
  reg  [4:0]  ldq_3_bits_uop_ldq_idx;
  reg  [4:0]  ldq_3_bits_uop_stq_idx;
  reg  [1:0]  ldq_3_bits_uop_rxq_idx;
  reg  [6:0]  ldq_3_bits_uop_pdst;
  reg  [6:0]  ldq_3_bits_uop_prs1;
  reg  [6:0]  ldq_3_bits_uop_prs2;
  reg  [6:0]  ldq_3_bits_uop_prs3;
  reg         ldq_3_bits_uop_prs1_busy;
  reg         ldq_3_bits_uop_prs2_busy;
  reg         ldq_3_bits_uop_prs3_busy;
  reg  [6:0]  ldq_3_bits_uop_stale_pdst;
  reg         ldq_3_bits_uop_exception;
  reg  [63:0] ldq_3_bits_uop_exc_cause;
  reg         ldq_3_bits_uop_bypassable;
  reg  [4:0]  ldq_3_bits_uop_mem_cmd;
  reg  [1:0]  ldq_3_bits_uop_mem_size;
  reg         ldq_3_bits_uop_mem_signed;
  reg         ldq_3_bits_uop_is_fence;
  reg         ldq_3_bits_uop_is_fencei;
  reg         ldq_3_bits_uop_is_amo;
  reg         ldq_3_bits_uop_uses_ldq;
  reg         ldq_3_bits_uop_uses_stq;
  reg         ldq_3_bits_uop_is_sys_pc2epc;
  reg         ldq_3_bits_uop_is_unique;
  reg         ldq_3_bits_uop_flush_on_commit;
  reg         ldq_3_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_3_bits_uop_ldst;
  reg  [5:0]  ldq_3_bits_uop_lrs1;
  reg  [5:0]  ldq_3_bits_uop_lrs2;
  reg  [5:0]  ldq_3_bits_uop_lrs3;
  reg         ldq_3_bits_uop_ldst_val;
  reg  [1:0]  ldq_3_bits_uop_dst_rtype;
  reg  [1:0]  ldq_3_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_3_bits_uop_lrs2_rtype;
  reg         ldq_3_bits_uop_frs3_en;
  reg         ldq_3_bits_uop_fp_val;
  reg         ldq_3_bits_uop_fp_single;
  reg         ldq_3_bits_uop_xcpt_pf_if;
  reg         ldq_3_bits_uop_xcpt_ae_if;
  reg         ldq_3_bits_uop_xcpt_ma_if;
  reg         ldq_3_bits_uop_bp_debug_if;
  reg         ldq_3_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_3_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_3_bits_uop_debug_tsrc;
  reg         ldq_3_bits_addr_valid;
  reg  [39:0] ldq_3_bits_addr_bits;
  reg         ldq_3_bits_addr_is_virtual;
  reg         ldq_3_bits_addr_is_uncacheable;
  reg         ldq_3_bits_executed;
  reg         ldq_3_bits_succeeded;
  reg         ldq_3_bits_order_fail;
  reg         ldq_3_bits_observed;
  reg  [31:0] ldq_3_bits_st_dep_mask;
  reg  [4:0]  ldq_3_bits_youngest_stq_idx;
  reg         ldq_3_bits_forward_std_val;
  reg  [4:0]  ldq_3_bits_forward_stq_idx;
  reg         ldq_4_valid;
  reg  [6:0]  ldq_4_bits_uop_uopc;
  reg  [31:0] ldq_4_bits_uop_inst;
  reg  [31:0] ldq_4_bits_uop_debug_inst;
  reg         ldq_4_bits_uop_is_rvc;
  reg  [39:0] ldq_4_bits_uop_debug_pc;
  reg  [2:0]  ldq_4_bits_uop_iq_type;
  reg  [9:0]  ldq_4_bits_uop_fu_code;
  reg  [3:0]  ldq_4_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_4_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_4_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_4_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_4_bits_uop_ctrl_op_fcn;
  reg         ldq_4_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_4_bits_uop_ctrl_csr_cmd;
  reg         ldq_4_bits_uop_ctrl_is_load;
  reg         ldq_4_bits_uop_ctrl_is_sta;
  reg         ldq_4_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_4_bits_uop_iw_state;
  reg         ldq_4_bits_uop_iw_p1_poisoned;
  reg         ldq_4_bits_uop_iw_p2_poisoned;
  reg         ldq_4_bits_uop_is_br;
  reg         ldq_4_bits_uop_is_jalr;
  reg         ldq_4_bits_uop_is_jal;
  reg         ldq_4_bits_uop_is_sfb;
  reg  [19:0] ldq_4_bits_uop_br_mask;
  reg  [4:0]  ldq_4_bits_uop_br_tag;
  reg  [5:0]  ldq_4_bits_uop_ftq_idx;
  reg         ldq_4_bits_uop_edge_inst;
  reg  [5:0]  ldq_4_bits_uop_pc_lob;
  reg         ldq_4_bits_uop_taken;
  reg  [19:0] ldq_4_bits_uop_imm_packed;
  reg  [11:0] ldq_4_bits_uop_csr_addr;
  reg  [6:0]  ldq_4_bits_uop_rob_idx;
  reg  [4:0]  ldq_4_bits_uop_ldq_idx;
  reg  [4:0]  ldq_4_bits_uop_stq_idx;
  reg  [1:0]  ldq_4_bits_uop_rxq_idx;
  reg  [6:0]  ldq_4_bits_uop_pdst;
  reg  [6:0]  ldq_4_bits_uop_prs1;
  reg  [6:0]  ldq_4_bits_uop_prs2;
  reg  [6:0]  ldq_4_bits_uop_prs3;
  reg         ldq_4_bits_uop_prs1_busy;
  reg         ldq_4_bits_uop_prs2_busy;
  reg         ldq_4_bits_uop_prs3_busy;
  reg  [6:0]  ldq_4_bits_uop_stale_pdst;
  reg         ldq_4_bits_uop_exception;
  reg  [63:0] ldq_4_bits_uop_exc_cause;
  reg         ldq_4_bits_uop_bypassable;
  reg  [4:0]  ldq_4_bits_uop_mem_cmd;
  reg  [1:0]  ldq_4_bits_uop_mem_size;
  reg         ldq_4_bits_uop_mem_signed;
  reg         ldq_4_bits_uop_is_fence;
  reg         ldq_4_bits_uop_is_fencei;
  reg         ldq_4_bits_uop_is_amo;
  reg         ldq_4_bits_uop_uses_ldq;
  reg         ldq_4_bits_uop_uses_stq;
  reg         ldq_4_bits_uop_is_sys_pc2epc;
  reg         ldq_4_bits_uop_is_unique;
  reg         ldq_4_bits_uop_flush_on_commit;
  reg         ldq_4_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_4_bits_uop_ldst;
  reg  [5:0]  ldq_4_bits_uop_lrs1;
  reg  [5:0]  ldq_4_bits_uop_lrs2;
  reg  [5:0]  ldq_4_bits_uop_lrs3;
  reg         ldq_4_bits_uop_ldst_val;
  reg  [1:0]  ldq_4_bits_uop_dst_rtype;
  reg  [1:0]  ldq_4_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_4_bits_uop_lrs2_rtype;
  reg         ldq_4_bits_uop_frs3_en;
  reg         ldq_4_bits_uop_fp_val;
  reg         ldq_4_bits_uop_fp_single;
  reg         ldq_4_bits_uop_xcpt_pf_if;
  reg         ldq_4_bits_uop_xcpt_ae_if;
  reg         ldq_4_bits_uop_xcpt_ma_if;
  reg         ldq_4_bits_uop_bp_debug_if;
  reg         ldq_4_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_4_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_4_bits_uop_debug_tsrc;
  reg         ldq_4_bits_addr_valid;
  reg  [39:0] ldq_4_bits_addr_bits;
  reg         ldq_4_bits_addr_is_virtual;
  reg         ldq_4_bits_addr_is_uncacheable;
  reg         ldq_4_bits_executed;
  reg         ldq_4_bits_succeeded;
  reg         ldq_4_bits_order_fail;
  reg         ldq_4_bits_observed;
  reg  [31:0] ldq_4_bits_st_dep_mask;
  reg  [4:0]  ldq_4_bits_youngest_stq_idx;
  reg         ldq_4_bits_forward_std_val;
  reg  [4:0]  ldq_4_bits_forward_stq_idx;
  reg         ldq_5_valid;
  reg  [6:0]  ldq_5_bits_uop_uopc;
  reg  [31:0] ldq_5_bits_uop_inst;
  reg  [31:0] ldq_5_bits_uop_debug_inst;
  reg         ldq_5_bits_uop_is_rvc;
  reg  [39:0] ldq_5_bits_uop_debug_pc;
  reg  [2:0]  ldq_5_bits_uop_iq_type;
  reg  [9:0]  ldq_5_bits_uop_fu_code;
  reg  [3:0]  ldq_5_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_5_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_5_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_5_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_5_bits_uop_ctrl_op_fcn;
  reg         ldq_5_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_5_bits_uop_ctrl_csr_cmd;
  reg         ldq_5_bits_uop_ctrl_is_load;
  reg         ldq_5_bits_uop_ctrl_is_sta;
  reg         ldq_5_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_5_bits_uop_iw_state;
  reg         ldq_5_bits_uop_iw_p1_poisoned;
  reg         ldq_5_bits_uop_iw_p2_poisoned;
  reg         ldq_5_bits_uop_is_br;
  reg         ldq_5_bits_uop_is_jalr;
  reg         ldq_5_bits_uop_is_jal;
  reg         ldq_5_bits_uop_is_sfb;
  reg  [19:0] ldq_5_bits_uop_br_mask;
  reg  [4:0]  ldq_5_bits_uop_br_tag;
  reg  [5:0]  ldq_5_bits_uop_ftq_idx;
  reg         ldq_5_bits_uop_edge_inst;
  reg  [5:0]  ldq_5_bits_uop_pc_lob;
  reg         ldq_5_bits_uop_taken;
  reg  [19:0] ldq_5_bits_uop_imm_packed;
  reg  [11:0] ldq_5_bits_uop_csr_addr;
  reg  [6:0]  ldq_5_bits_uop_rob_idx;
  reg  [4:0]  ldq_5_bits_uop_ldq_idx;
  reg  [4:0]  ldq_5_bits_uop_stq_idx;
  reg  [1:0]  ldq_5_bits_uop_rxq_idx;
  reg  [6:0]  ldq_5_bits_uop_pdst;
  reg  [6:0]  ldq_5_bits_uop_prs1;
  reg  [6:0]  ldq_5_bits_uop_prs2;
  reg  [6:0]  ldq_5_bits_uop_prs3;
  reg         ldq_5_bits_uop_prs1_busy;
  reg         ldq_5_bits_uop_prs2_busy;
  reg         ldq_5_bits_uop_prs3_busy;
  reg  [6:0]  ldq_5_bits_uop_stale_pdst;
  reg         ldq_5_bits_uop_exception;
  reg  [63:0] ldq_5_bits_uop_exc_cause;
  reg         ldq_5_bits_uop_bypassable;
  reg  [4:0]  ldq_5_bits_uop_mem_cmd;
  reg  [1:0]  ldq_5_bits_uop_mem_size;
  reg         ldq_5_bits_uop_mem_signed;
  reg         ldq_5_bits_uop_is_fence;
  reg         ldq_5_bits_uop_is_fencei;
  reg         ldq_5_bits_uop_is_amo;
  reg         ldq_5_bits_uop_uses_ldq;
  reg         ldq_5_bits_uop_uses_stq;
  reg         ldq_5_bits_uop_is_sys_pc2epc;
  reg         ldq_5_bits_uop_is_unique;
  reg         ldq_5_bits_uop_flush_on_commit;
  reg         ldq_5_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_5_bits_uop_ldst;
  reg  [5:0]  ldq_5_bits_uop_lrs1;
  reg  [5:0]  ldq_5_bits_uop_lrs2;
  reg  [5:0]  ldq_5_bits_uop_lrs3;
  reg         ldq_5_bits_uop_ldst_val;
  reg  [1:0]  ldq_5_bits_uop_dst_rtype;
  reg  [1:0]  ldq_5_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_5_bits_uop_lrs2_rtype;
  reg         ldq_5_bits_uop_frs3_en;
  reg         ldq_5_bits_uop_fp_val;
  reg         ldq_5_bits_uop_fp_single;
  reg         ldq_5_bits_uop_xcpt_pf_if;
  reg         ldq_5_bits_uop_xcpt_ae_if;
  reg         ldq_5_bits_uop_xcpt_ma_if;
  reg         ldq_5_bits_uop_bp_debug_if;
  reg         ldq_5_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_5_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_5_bits_uop_debug_tsrc;
  reg         ldq_5_bits_addr_valid;
  reg  [39:0] ldq_5_bits_addr_bits;
  reg         ldq_5_bits_addr_is_virtual;
  reg         ldq_5_bits_addr_is_uncacheable;
  reg         ldq_5_bits_executed;
  reg         ldq_5_bits_succeeded;
  reg         ldq_5_bits_order_fail;
  reg         ldq_5_bits_observed;
  reg  [31:0] ldq_5_bits_st_dep_mask;
  reg  [4:0]  ldq_5_bits_youngest_stq_idx;
  reg         ldq_5_bits_forward_std_val;
  reg  [4:0]  ldq_5_bits_forward_stq_idx;
  reg         ldq_6_valid;
  reg  [6:0]  ldq_6_bits_uop_uopc;
  reg  [31:0] ldq_6_bits_uop_inst;
  reg  [31:0] ldq_6_bits_uop_debug_inst;
  reg         ldq_6_bits_uop_is_rvc;
  reg  [39:0] ldq_6_bits_uop_debug_pc;
  reg  [2:0]  ldq_6_bits_uop_iq_type;
  reg  [9:0]  ldq_6_bits_uop_fu_code;
  reg  [3:0]  ldq_6_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_6_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_6_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_6_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_6_bits_uop_ctrl_op_fcn;
  reg         ldq_6_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_6_bits_uop_ctrl_csr_cmd;
  reg         ldq_6_bits_uop_ctrl_is_load;
  reg         ldq_6_bits_uop_ctrl_is_sta;
  reg         ldq_6_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_6_bits_uop_iw_state;
  reg         ldq_6_bits_uop_iw_p1_poisoned;
  reg         ldq_6_bits_uop_iw_p2_poisoned;
  reg         ldq_6_bits_uop_is_br;
  reg         ldq_6_bits_uop_is_jalr;
  reg         ldq_6_bits_uop_is_jal;
  reg         ldq_6_bits_uop_is_sfb;
  reg  [19:0] ldq_6_bits_uop_br_mask;
  reg  [4:0]  ldq_6_bits_uop_br_tag;
  reg  [5:0]  ldq_6_bits_uop_ftq_idx;
  reg         ldq_6_bits_uop_edge_inst;
  reg  [5:0]  ldq_6_bits_uop_pc_lob;
  reg         ldq_6_bits_uop_taken;
  reg  [19:0] ldq_6_bits_uop_imm_packed;
  reg  [11:0] ldq_6_bits_uop_csr_addr;
  reg  [6:0]  ldq_6_bits_uop_rob_idx;
  reg  [4:0]  ldq_6_bits_uop_ldq_idx;
  reg  [4:0]  ldq_6_bits_uop_stq_idx;
  reg  [1:0]  ldq_6_bits_uop_rxq_idx;
  reg  [6:0]  ldq_6_bits_uop_pdst;
  reg  [6:0]  ldq_6_bits_uop_prs1;
  reg  [6:0]  ldq_6_bits_uop_prs2;
  reg  [6:0]  ldq_6_bits_uop_prs3;
  reg         ldq_6_bits_uop_prs1_busy;
  reg         ldq_6_bits_uop_prs2_busy;
  reg         ldq_6_bits_uop_prs3_busy;
  reg  [6:0]  ldq_6_bits_uop_stale_pdst;
  reg         ldq_6_bits_uop_exception;
  reg  [63:0] ldq_6_bits_uop_exc_cause;
  reg         ldq_6_bits_uop_bypassable;
  reg  [4:0]  ldq_6_bits_uop_mem_cmd;
  reg  [1:0]  ldq_6_bits_uop_mem_size;
  reg         ldq_6_bits_uop_mem_signed;
  reg         ldq_6_bits_uop_is_fence;
  reg         ldq_6_bits_uop_is_fencei;
  reg         ldq_6_bits_uop_is_amo;
  reg         ldq_6_bits_uop_uses_ldq;
  reg         ldq_6_bits_uop_uses_stq;
  reg         ldq_6_bits_uop_is_sys_pc2epc;
  reg         ldq_6_bits_uop_is_unique;
  reg         ldq_6_bits_uop_flush_on_commit;
  reg         ldq_6_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_6_bits_uop_ldst;
  reg  [5:0]  ldq_6_bits_uop_lrs1;
  reg  [5:0]  ldq_6_bits_uop_lrs2;
  reg  [5:0]  ldq_6_bits_uop_lrs3;
  reg         ldq_6_bits_uop_ldst_val;
  reg  [1:0]  ldq_6_bits_uop_dst_rtype;
  reg  [1:0]  ldq_6_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_6_bits_uop_lrs2_rtype;
  reg         ldq_6_bits_uop_frs3_en;
  reg         ldq_6_bits_uop_fp_val;
  reg         ldq_6_bits_uop_fp_single;
  reg         ldq_6_bits_uop_xcpt_pf_if;
  reg         ldq_6_bits_uop_xcpt_ae_if;
  reg         ldq_6_bits_uop_xcpt_ma_if;
  reg         ldq_6_bits_uop_bp_debug_if;
  reg         ldq_6_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_6_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_6_bits_uop_debug_tsrc;
  reg         ldq_6_bits_addr_valid;
  reg  [39:0] ldq_6_bits_addr_bits;
  reg         ldq_6_bits_addr_is_virtual;
  reg         ldq_6_bits_addr_is_uncacheable;
  reg         ldq_6_bits_executed;
  reg         ldq_6_bits_succeeded;
  reg         ldq_6_bits_order_fail;
  reg         ldq_6_bits_observed;
  reg  [31:0] ldq_6_bits_st_dep_mask;
  reg  [4:0]  ldq_6_bits_youngest_stq_idx;
  reg         ldq_6_bits_forward_std_val;
  reg  [4:0]  ldq_6_bits_forward_stq_idx;
  reg         ldq_7_valid;
  reg  [6:0]  ldq_7_bits_uop_uopc;
  reg  [31:0] ldq_7_bits_uop_inst;
  reg  [31:0] ldq_7_bits_uop_debug_inst;
  reg         ldq_7_bits_uop_is_rvc;
  reg  [39:0] ldq_7_bits_uop_debug_pc;
  reg  [2:0]  ldq_7_bits_uop_iq_type;
  reg  [9:0]  ldq_7_bits_uop_fu_code;
  reg  [3:0]  ldq_7_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_7_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_7_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_7_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_7_bits_uop_ctrl_op_fcn;
  reg         ldq_7_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_7_bits_uop_ctrl_csr_cmd;
  reg         ldq_7_bits_uop_ctrl_is_load;
  reg         ldq_7_bits_uop_ctrl_is_sta;
  reg         ldq_7_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_7_bits_uop_iw_state;
  reg         ldq_7_bits_uop_iw_p1_poisoned;
  reg         ldq_7_bits_uop_iw_p2_poisoned;
  reg         ldq_7_bits_uop_is_br;
  reg         ldq_7_bits_uop_is_jalr;
  reg         ldq_7_bits_uop_is_jal;
  reg         ldq_7_bits_uop_is_sfb;
  reg  [19:0] ldq_7_bits_uop_br_mask;
  reg  [4:0]  ldq_7_bits_uop_br_tag;
  reg  [5:0]  ldq_7_bits_uop_ftq_idx;
  reg         ldq_7_bits_uop_edge_inst;
  reg  [5:0]  ldq_7_bits_uop_pc_lob;
  reg         ldq_7_bits_uop_taken;
  reg  [19:0] ldq_7_bits_uop_imm_packed;
  reg  [11:0] ldq_7_bits_uop_csr_addr;
  reg  [6:0]  ldq_7_bits_uop_rob_idx;
  reg  [4:0]  ldq_7_bits_uop_ldq_idx;
  reg  [4:0]  ldq_7_bits_uop_stq_idx;
  reg  [1:0]  ldq_7_bits_uop_rxq_idx;
  reg  [6:0]  ldq_7_bits_uop_pdst;
  reg  [6:0]  ldq_7_bits_uop_prs1;
  reg  [6:0]  ldq_7_bits_uop_prs2;
  reg  [6:0]  ldq_7_bits_uop_prs3;
  reg         ldq_7_bits_uop_prs1_busy;
  reg         ldq_7_bits_uop_prs2_busy;
  reg         ldq_7_bits_uop_prs3_busy;
  reg  [6:0]  ldq_7_bits_uop_stale_pdst;
  reg         ldq_7_bits_uop_exception;
  reg  [63:0] ldq_7_bits_uop_exc_cause;
  reg         ldq_7_bits_uop_bypassable;
  reg  [4:0]  ldq_7_bits_uop_mem_cmd;
  reg  [1:0]  ldq_7_bits_uop_mem_size;
  reg         ldq_7_bits_uop_mem_signed;
  reg         ldq_7_bits_uop_is_fence;
  reg         ldq_7_bits_uop_is_fencei;
  reg         ldq_7_bits_uop_is_amo;
  reg         ldq_7_bits_uop_uses_ldq;
  reg         ldq_7_bits_uop_uses_stq;
  reg         ldq_7_bits_uop_is_sys_pc2epc;
  reg         ldq_7_bits_uop_is_unique;
  reg         ldq_7_bits_uop_flush_on_commit;
  reg         ldq_7_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_7_bits_uop_ldst;
  reg  [5:0]  ldq_7_bits_uop_lrs1;
  reg  [5:0]  ldq_7_bits_uop_lrs2;
  reg  [5:0]  ldq_7_bits_uop_lrs3;
  reg         ldq_7_bits_uop_ldst_val;
  reg  [1:0]  ldq_7_bits_uop_dst_rtype;
  reg  [1:0]  ldq_7_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_7_bits_uop_lrs2_rtype;
  reg         ldq_7_bits_uop_frs3_en;
  reg         ldq_7_bits_uop_fp_val;
  reg         ldq_7_bits_uop_fp_single;
  reg         ldq_7_bits_uop_xcpt_pf_if;
  reg         ldq_7_bits_uop_xcpt_ae_if;
  reg         ldq_7_bits_uop_xcpt_ma_if;
  reg         ldq_7_bits_uop_bp_debug_if;
  reg         ldq_7_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_7_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_7_bits_uop_debug_tsrc;
  reg         ldq_7_bits_addr_valid;
  reg  [39:0] ldq_7_bits_addr_bits;
  reg         ldq_7_bits_addr_is_virtual;
  reg         ldq_7_bits_addr_is_uncacheable;
  reg         ldq_7_bits_executed;
  reg         ldq_7_bits_succeeded;
  reg         ldq_7_bits_order_fail;
  reg         ldq_7_bits_observed;
  reg  [31:0] ldq_7_bits_st_dep_mask;
  reg  [4:0]  ldq_7_bits_youngest_stq_idx;
  reg         ldq_7_bits_forward_std_val;
  reg  [4:0]  ldq_7_bits_forward_stq_idx;
  reg         ldq_8_valid;
  reg  [6:0]  ldq_8_bits_uop_uopc;
  reg  [31:0] ldq_8_bits_uop_inst;
  reg  [31:0] ldq_8_bits_uop_debug_inst;
  reg         ldq_8_bits_uop_is_rvc;
  reg  [39:0] ldq_8_bits_uop_debug_pc;
  reg  [2:0]  ldq_8_bits_uop_iq_type;
  reg  [9:0]  ldq_8_bits_uop_fu_code;
  reg  [3:0]  ldq_8_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_8_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_8_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_8_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_8_bits_uop_ctrl_op_fcn;
  reg         ldq_8_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_8_bits_uop_ctrl_csr_cmd;
  reg         ldq_8_bits_uop_ctrl_is_load;
  reg         ldq_8_bits_uop_ctrl_is_sta;
  reg         ldq_8_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_8_bits_uop_iw_state;
  reg         ldq_8_bits_uop_iw_p1_poisoned;
  reg         ldq_8_bits_uop_iw_p2_poisoned;
  reg         ldq_8_bits_uop_is_br;
  reg         ldq_8_bits_uop_is_jalr;
  reg         ldq_8_bits_uop_is_jal;
  reg         ldq_8_bits_uop_is_sfb;
  reg  [19:0] ldq_8_bits_uop_br_mask;
  reg  [4:0]  ldq_8_bits_uop_br_tag;
  reg  [5:0]  ldq_8_bits_uop_ftq_idx;
  reg         ldq_8_bits_uop_edge_inst;
  reg  [5:0]  ldq_8_bits_uop_pc_lob;
  reg         ldq_8_bits_uop_taken;
  reg  [19:0] ldq_8_bits_uop_imm_packed;
  reg  [11:0] ldq_8_bits_uop_csr_addr;
  reg  [6:0]  ldq_8_bits_uop_rob_idx;
  reg  [4:0]  ldq_8_bits_uop_ldq_idx;
  reg  [4:0]  ldq_8_bits_uop_stq_idx;
  reg  [1:0]  ldq_8_bits_uop_rxq_idx;
  reg  [6:0]  ldq_8_bits_uop_pdst;
  reg  [6:0]  ldq_8_bits_uop_prs1;
  reg  [6:0]  ldq_8_bits_uop_prs2;
  reg  [6:0]  ldq_8_bits_uop_prs3;
  reg         ldq_8_bits_uop_prs1_busy;
  reg         ldq_8_bits_uop_prs2_busy;
  reg         ldq_8_bits_uop_prs3_busy;
  reg  [6:0]  ldq_8_bits_uop_stale_pdst;
  reg         ldq_8_bits_uop_exception;
  reg  [63:0] ldq_8_bits_uop_exc_cause;
  reg         ldq_8_bits_uop_bypassable;
  reg  [4:0]  ldq_8_bits_uop_mem_cmd;
  reg  [1:0]  ldq_8_bits_uop_mem_size;
  reg         ldq_8_bits_uop_mem_signed;
  reg         ldq_8_bits_uop_is_fence;
  reg         ldq_8_bits_uop_is_fencei;
  reg         ldq_8_bits_uop_is_amo;
  reg         ldq_8_bits_uop_uses_ldq;
  reg         ldq_8_bits_uop_uses_stq;
  reg         ldq_8_bits_uop_is_sys_pc2epc;
  reg         ldq_8_bits_uop_is_unique;
  reg         ldq_8_bits_uop_flush_on_commit;
  reg         ldq_8_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_8_bits_uop_ldst;
  reg  [5:0]  ldq_8_bits_uop_lrs1;
  reg  [5:0]  ldq_8_bits_uop_lrs2;
  reg  [5:0]  ldq_8_bits_uop_lrs3;
  reg         ldq_8_bits_uop_ldst_val;
  reg  [1:0]  ldq_8_bits_uop_dst_rtype;
  reg  [1:0]  ldq_8_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_8_bits_uop_lrs2_rtype;
  reg         ldq_8_bits_uop_frs3_en;
  reg         ldq_8_bits_uop_fp_val;
  reg         ldq_8_bits_uop_fp_single;
  reg         ldq_8_bits_uop_xcpt_pf_if;
  reg         ldq_8_bits_uop_xcpt_ae_if;
  reg         ldq_8_bits_uop_xcpt_ma_if;
  reg         ldq_8_bits_uop_bp_debug_if;
  reg         ldq_8_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_8_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_8_bits_uop_debug_tsrc;
  reg         ldq_8_bits_addr_valid;
  reg  [39:0] ldq_8_bits_addr_bits;
  reg         ldq_8_bits_addr_is_virtual;
  reg         ldq_8_bits_addr_is_uncacheable;
  reg         ldq_8_bits_executed;
  reg         ldq_8_bits_succeeded;
  reg         ldq_8_bits_order_fail;
  reg         ldq_8_bits_observed;
  reg  [31:0] ldq_8_bits_st_dep_mask;
  reg  [4:0]  ldq_8_bits_youngest_stq_idx;
  reg         ldq_8_bits_forward_std_val;
  reg  [4:0]  ldq_8_bits_forward_stq_idx;
  reg         ldq_9_valid;
  reg  [6:0]  ldq_9_bits_uop_uopc;
  reg  [31:0] ldq_9_bits_uop_inst;
  reg  [31:0] ldq_9_bits_uop_debug_inst;
  reg         ldq_9_bits_uop_is_rvc;
  reg  [39:0] ldq_9_bits_uop_debug_pc;
  reg  [2:0]  ldq_9_bits_uop_iq_type;
  reg  [9:0]  ldq_9_bits_uop_fu_code;
  reg  [3:0]  ldq_9_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_9_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_9_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_9_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_9_bits_uop_ctrl_op_fcn;
  reg         ldq_9_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_9_bits_uop_ctrl_csr_cmd;
  reg         ldq_9_bits_uop_ctrl_is_load;
  reg         ldq_9_bits_uop_ctrl_is_sta;
  reg         ldq_9_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_9_bits_uop_iw_state;
  reg         ldq_9_bits_uop_iw_p1_poisoned;
  reg         ldq_9_bits_uop_iw_p2_poisoned;
  reg         ldq_9_bits_uop_is_br;
  reg         ldq_9_bits_uop_is_jalr;
  reg         ldq_9_bits_uop_is_jal;
  reg         ldq_9_bits_uop_is_sfb;
  reg  [19:0] ldq_9_bits_uop_br_mask;
  reg  [4:0]  ldq_9_bits_uop_br_tag;
  reg  [5:0]  ldq_9_bits_uop_ftq_idx;
  reg         ldq_9_bits_uop_edge_inst;
  reg  [5:0]  ldq_9_bits_uop_pc_lob;
  reg         ldq_9_bits_uop_taken;
  reg  [19:0] ldq_9_bits_uop_imm_packed;
  reg  [11:0] ldq_9_bits_uop_csr_addr;
  reg  [6:0]  ldq_9_bits_uop_rob_idx;
  reg  [4:0]  ldq_9_bits_uop_ldq_idx;
  reg  [4:0]  ldq_9_bits_uop_stq_idx;
  reg  [1:0]  ldq_9_bits_uop_rxq_idx;
  reg  [6:0]  ldq_9_bits_uop_pdst;
  reg  [6:0]  ldq_9_bits_uop_prs1;
  reg  [6:0]  ldq_9_bits_uop_prs2;
  reg  [6:0]  ldq_9_bits_uop_prs3;
  reg         ldq_9_bits_uop_prs1_busy;
  reg         ldq_9_bits_uop_prs2_busy;
  reg         ldq_9_bits_uop_prs3_busy;
  reg  [6:0]  ldq_9_bits_uop_stale_pdst;
  reg         ldq_9_bits_uop_exception;
  reg  [63:0] ldq_9_bits_uop_exc_cause;
  reg         ldq_9_bits_uop_bypassable;
  reg  [4:0]  ldq_9_bits_uop_mem_cmd;
  reg  [1:0]  ldq_9_bits_uop_mem_size;
  reg         ldq_9_bits_uop_mem_signed;
  reg         ldq_9_bits_uop_is_fence;
  reg         ldq_9_bits_uop_is_fencei;
  reg         ldq_9_bits_uop_is_amo;
  reg         ldq_9_bits_uop_uses_ldq;
  reg         ldq_9_bits_uop_uses_stq;
  reg         ldq_9_bits_uop_is_sys_pc2epc;
  reg         ldq_9_bits_uop_is_unique;
  reg         ldq_9_bits_uop_flush_on_commit;
  reg         ldq_9_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_9_bits_uop_ldst;
  reg  [5:0]  ldq_9_bits_uop_lrs1;
  reg  [5:0]  ldq_9_bits_uop_lrs2;
  reg  [5:0]  ldq_9_bits_uop_lrs3;
  reg         ldq_9_bits_uop_ldst_val;
  reg  [1:0]  ldq_9_bits_uop_dst_rtype;
  reg  [1:0]  ldq_9_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_9_bits_uop_lrs2_rtype;
  reg         ldq_9_bits_uop_frs3_en;
  reg         ldq_9_bits_uop_fp_val;
  reg         ldq_9_bits_uop_fp_single;
  reg         ldq_9_bits_uop_xcpt_pf_if;
  reg         ldq_9_bits_uop_xcpt_ae_if;
  reg         ldq_9_bits_uop_xcpt_ma_if;
  reg         ldq_9_bits_uop_bp_debug_if;
  reg         ldq_9_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_9_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_9_bits_uop_debug_tsrc;
  reg         ldq_9_bits_addr_valid;
  reg  [39:0] ldq_9_bits_addr_bits;
  reg         ldq_9_bits_addr_is_virtual;
  reg         ldq_9_bits_addr_is_uncacheable;
  reg         ldq_9_bits_executed;
  reg         ldq_9_bits_succeeded;
  reg         ldq_9_bits_order_fail;
  reg         ldq_9_bits_observed;
  reg  [31:0] ldq_9_bits_st_dep_mask;
  reg  [4:0]  ldq_9_bits_youngest_stq_idx;
  reg         ldq_9_bits_forward_std_val;
  reg  [4:0]  ldq_9_bits_forward_stq_idx;
  reg         ldq_10_valid;
  reg  [6:0]  ldq_10_bits_uop_uopc;
  reg  [31:0] ldq_10_bits_uop_inst;
  reg  [31:0] ldq_10_bits_uop_debug_inst;
  reg         ldq_10_bits_uop_is_rvc;
  reg  [39:0] ldq_10_bits_uop_debug_pc;
  reg  [2:0]  ldq_10_bits_uop_iq_type;
  reg  [9:0]  ldq_10_bits_uop_fu_code;
  reg  [3:0]  ldq_10_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_10_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_10_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_10_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_10_bits_uop_ctrl_op_fcn;
  reg         ldq_10_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_10_bits_uop_ctrl_csr_cmd;
  reg         ldq_10_bits_uop_ctrl_is_load;
  reg         ldq_10_bits_uop_ctrl_is_sta;
  reg         ldq_10_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_10_bits_uop_iw_state;
  reg         ldq_10_bits_uop_iw_p1_poisoned;
  reg         ldq_10_bits_uop_iw_p2_poisoned;
  reg         ldq_10_bits_uop_is_br;
  reg         ldq_10_bits_uop_is_jalr;
  reg         ldq_10_bits_uop_is_jal;
  reg         ldq_10_bits_uop_is_sfb;
  reg  [19:0] ldq_10_bits_uop_br_mask;
  reg  [4:0]  ldq_10_bits_uop_br_tag;
  reg  [5:0]  ldq_10_bits_uop_ftq_idx;
  reg         ldq_10_bits_uop_edge_inst;
  reg  [5:0]  ldq_10_bits_uop_pc_lob;
  reg         ldq_10_bits_uop_taken;
  reg  [19:0] ldq_10_bits_uop_imm_packed;
  reg  [11:0] ldq_10_bits_uop_csr_addr;
  reg  [6:0]  ldq_10_bits_uop_rob_idx;
  reg  [4:0]  ldq_10_bits_uop_ldq_idx;
  reg  [4:0]  ldq_10_bits_uop_stq_idx;
  reg  [1:0]  ldq_10_bits_uop_rxq_idx;
  reg  [6:0]  ldq_10_bits_uop_pdst;
  reg  [6:0]  ldq_10_bits_uop_prs1;
  reg  [6:0]  ldq_10_bits_uop_prs2;
  reg  [6:0]  ldq_10_bits_uop_prs3;
  reg         ldq_10_bits_uop_prs1_busy;
  reg         ldq_10_bits_uop_prs2_busy;
  reg         ldq_10_bits_uop_prs3_busy;
  reg  [6:0]  ldq_10_bits_uop_stale_pdst;
  reg         ldq_10_bits_uop_exception;
  reg  [63:0] ldq_10_bits_uop_exc_cause;
  reg         ldq_10_bits_uop_bypassable;
  reg  [4:0]  ldq_10_bits_uop_mem_cmd;
  reg  [1:0]  ldq_10_bits_uop_mem_size;
  reg         ldq_10_bits_uop_mem_signed;
  reg         ldq_10_bits_uop_is_fence;
  reg         ldq_10_bits_uop_is_fencei;
  reg         ldq_10_bits_uop_is_amo;
  reg         ldq_10_bits_uop_uses_ldq;
  reg         ldq_10_bits_uop_uses_stq;
  reg         ldq_10_bits_uop_is_sys_pc2epc;
  reg         ldq_10_bits_uop_is_unique;
  reg         ldq_10_bits_uop_flush_on_commit;
  reg         ldq_10_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_10_bits_uop_ldst;
  reg  [5:0]  ldq_10_bits_uop_lrs1;
  reg  [5:0]  ldq_10_bits_uop_lrs2;
  reg  [5:0]  ldq_10_bits_uop_lrs3;
  reg         ldq_10_bits_uop_ldst_val;
  reg  [1:0]  ldq_10_bits_uop_dst_rtype;
  reg  [1:0]  ldq_10_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_10_bits_uop_lrs2_rtype;
  reg         ldq_10_bits_uop_frs3_en;
  reg         ldq_10_bits_uop_fp_val;
  reg         ldq_10_bits_uop_fp_single;
  reg         ldq_10_bits_uop_xcpt_pf_if;
  reg         ldq_10_bits_uop_xcpt_ae_if;
  reg         ldq_10_bits_uop_xcpt_ma_if;
  reg         ldq_10_bits_uop_bp_debug_if;
  reg         ldq_10_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_10_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_10_bits_uop_debug_tsrc;
  reg         ldq_10_bits_addr_valid;
  reg  [39:0] ldq_10_bits_addr_bits;
  reg         ldq_10_bits_addr_is_virtual;
  reg         ldq_10_bits_addr_is_uncacheable;
  reg         ldq_10_bits_executed;
  reg         ldq_10_bits_succeeded;
  reg         ldq_10_bits_order_fail;
  reg         ldq_10_bits_observed;
  reg  [31:0] ldq_10_bits_st_dep_mask;
  reg  [4:0]  ldq_10_bits_youngest_stq_idx;
  reg         ldq_10_bits_forward_std_val;
  reg  [4:0]  ldq_10_bits_forward_stq_idx;
  reg         ldq_11_valid;
  reg  [6:0]  ldq_11_bits_uop_uopc;
  reg  [31:0] ldq_11_bits_uop_inst;
  reg  [31:0] ldq_11_bits_uop_debug_inst;
  reg         ldq_11_bits_uop_is_rvc;
  reg  [39:0] ldq_11_bits_uop_debug_pc;
  reg  [2:0]  ldq_11_bits_uop_iq_type;
  reg  [9:0]  ldq_11_bits_uop_fu_code;
  reg  [3:0]  ldq_11_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_11_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_11_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_11_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_11_bits_uop_ctrl_op_fcn;
  reg         ldq_11_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_11_bits_uop_ctrl_csr_cmd;
  reg         ldq_11_bits_uop_ctrl_is_load;
  reg         ldq_11_bits_uop_ctrl_is_sta;
  reg         ldq_11_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_11_bits_uop_iw_state;
  reg         ldq_11_bits_uop_iw_p1_poisoned;
  reg         ldq_11_bits_uop_iw_p2_poisoned;
  reg         ldq_11_bits_uop_is_br;
  reg         ldq_11_bits_uop_is_jalr;
  reg         ldq_11_bits_uop_is_jal;
  reg         ldq_11_bits_uop_is_sfb;
  reg  [19:0] ldq_11_bits_uop_br_mask;
  reg  [4:0]  ldq_11_bits_uop_br_tag;
  reg  [5:0]  ldq_11_bits_uop_ftq_idx;
  reg         ldq_11_bits_uop_edge_inst;
  reg  [5:0]  ldq_11_bits_uop_pc_lob;
  reg         ldq_11_bits_uop_taken;
  reg  [19:0] ldq_11_bits_uop_imm_packed;
  reg  [11:0] ldq_11_bits_uop_csr_addr;
  reg  [6:0]  ldq_11_bits_uop_rob_idx;
  reg  [4:0]  ldq_11_bits_uop_ldq_idx;
  reg  [4:0]  ldq_11_bits_uop_stq_idx;
  reg  [1:0]  ldq_11_bits_uop_rxq_idx;
  reg  [6:0]  ldq_11_bits_uop_pdst;
  reg  [6:0]  ldq_11_bits_uop_prs1;
  reg  [6:0]  ldq_11_bits_uop_prs2;
  reg  [6:0]  ldq_11_bits_uop_prs3;
  reg         ldq_11_bits_uop_prs1_busy;
  reg         ldq_11_bits_uop_prs2_busy;
  reg         ldq_11_bits_uop_prs3_busy;
  reg  [6:0]  ldq_11_bits_uop_stale_pdst;
  reg         ldq_11_bits_uop_exception;
  reg  [63:0] ldq_11_bits_uop_exc_cause;
  reg         ldq_11_bits_uop_bypassable;
  reg  [4:0]  ldq_11_bits_uop_mem_cmd;
  reg  [1:0]  ldq_11_bits_uop_mem_size;
  reg         ldq_11_bits_uop_mem_signed;
  reg         ldq_11_bits_uop_is_fence;
  reg         ldq_11_bits_uop_is_fencei;
  reg         ldq_11_bits_uop_is_amo;
  reg         ldq_11_bits_uop_uses_ldq;
  reg         ldq_11_bits_uop_uses_stq;
  reg         ldq_11_bits_uop_is_sys_pc2epc;
  reg         ldq_11_bits_uop_is_unique;
  reg         ldq_11_bits_uop_flush_on_commit;
  reg         ldq_11_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_11_bits_uop_ldst;
  reg  [5:0]  ldq_11_bits_uop_lrs1;
  reg  [5:0]  ldq_11_bits_uop_lrs2;
  reg  [5:0]  ldq_11_bits_uop_lrs3;
  reg         ldq_11_bits_uop_ldst_val;
  reg  [1:0]  ldq_11_bits_uop_dst_rtype;
  reg  [1:0]  ldq_11_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_11_bits_uop_lrs2_rtype;
  reg         ldq_11_bits_uop_frs3_en;
  reg         ldq_11_bits_uop_fp_val;
  reg         ldq_11_bits_uop_fp_single;
  reg         ldq_11_bits_uop_xcpt_pf_if;
  reg         ldq_11_bits_uop_xcpt_ae_if;
  reg         ldq_11_bits_uop_xcpt_ma_if;
  reg         ldq_11_bits_uop_bp_debug_if;
  reg         ldq_11_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_11_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_11_bits_uop_debug_tsrc;
  reg         ldq_11_bits_addr_valid;
  reg  [39:0] ldq_11_bits_addr_bits;
  reg         ldq_11_bits_addr_is_virtual;
  reg         ldq_11_bits_addr_is_uncacheable;
  reg         ldq_11_bits_executed;
  reg         ldq_11_bits_succeeded;
  reg         ldq_11_bits_order_fail;
  reg         ldq_11_bits_observed;
  reg  [31:0] ldq_11_bits_st_dep_mask;
  reg  [4:0]  ldq_11_bits_youngest_stq_idx;
  reg         ldq_11_bits_forward_std_val;
  reg  [4:0]  ldq_11_bits_forward_stq_idx;
  reg         ldq_12_valid;
  reg  [6:0]  ldq_12_bits_uop_uopc;
  reg  [31:0] ldq_12_bits_uop_inst;
  reg  [31:0] ldq_12_bits_uop_debug_inst;
  reg         ldq_12_bits_uop_is_rvc;
  reg  [39:0] ldq_12_bits_uop_debug_pc;
  reg  [2:0]  ldq_12_bits_uop_iq_type;
  reg  [9:0]  ldq_12_bits_uop_fu_code;
  reg  [3:0]  ldq_12_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_12_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_12_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_12_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_12_bits_uop_ctrl_op_fcn;
  reg         ldq_12_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_12_bits_uop_ctrl_csr_cmd;
  reg         ldq_12_bits_uop_ctrl_is_load;
  reg         ldq_12_bits_uop_ctrl_is_sta;
  reg         ldq_12_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_12_bits_uop_iw_state;
  reg         ldq_12_bits_uop_iw_p1_poisoned;
  reg         ldq_12_bits_uop_iw_p2_poisoned;
  reg         ldq_12_bits_uop_is_br;
  reg         ldq_12_bits_uop_is_jalr;
  reg         ldq_12_bits_uop_is_jal;
  reg         ldq_12_bits_uop_is_sfb;
  reg  [19:0] ldq_12_bits_uop_br_mask;
  reg  [4:0]  ldq_12_bits_uop_br_tag;
  reg  [5:0]  ldq_12_bits_uop_ftq_idx;
  reg         ldq_12_bits_uop_edge_inst;
  reg  [5:0]  ldq_12_bits_uop_pc_lob;
  reg         ldq_12_bits_uop_taken;
  reg  [19:0] ldq_12_bits_uop_imm_packed;
  reg  [11:0] ldq_12_bits_uop_csr_addr;
  reg  [6:0]  ldq_12_bits_uop_rob_idx;
  reg  [4:0]  ldq_12_bits_uop_ldq_idx;
  reg  [4:0]  ldq_12_bits_uop_stq_idx;
  reg  [1:0]  ldq_12_bits_uop_rxq_idx;
  reg  [6:0]  ldq_12_bits_uop_pdst;
  reg  [6:0]  ldq_12_bits_uop_prs1;
  reg  [6:0]  ldq_12_bits_uop_prs2;
  reg  [6:0]  ldq_12_bits_uop_prs3;
  reg         ldq_12_bits_uop_prs1_busy;
  reg         ldq_12_bits_uop_prs2_busy;
  reg         ldq_12_bits_uop_prs3_busy;
  reg  [6:0]  ldq_12_bits_uop_stale_pdst;
  reg         ldq_12_bits_uop_exception;
  reg  [63:0] ldq_12_bits_uop_exc_cause;
  reg         ldq_12_bits_uop_bypassable;
  reg  [4:0]  ldq_12_bits_uop_mem_cmd;
  reg  [1:0]  ldq_12_bits_uop_mem_size;
  reg         ldq_12_bits_uop_mem_signed;
  reg         ldq_12_bits_uop_is_fence;
  reg         ldq_12_bits_uop_is_fencei;
  reg         ldq_12_bits_uop_is_amo;
  reg         ldq_12_bits_uop_uses_ldq;
  reg         ldq_12_bits_uop_uses_stq;
  reg         ldq_12_bits_uop_is_sys_pc2epc;
  reg         ldq_12_bits_uop_is_unique;
  reg         ldq_12_bits_uop_flush_on_commit;
  reg         ldq_12_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_12_bits_uop_ldst;
  reg  [5:0]  ldq_12_bits_uop_lrs1;
  reg  [5:0]  ldq_12_bits_uop_lrs2;
  reg  [5:0]  ldq_12_bits_uop_lrs3;
  reg         ldq_12_bits_uop_ldst_val;
  reg  [1:0]  ldq_12_bits_uop_dst_rtype;
  reg  [1:0]  ldq_12_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_12_bits_uop_lrs2_rtype;
  reg         ldq_12_bits_uop_frs3_en;
  reg         ldq_12_bits_uop_fp_val;
  reg         ldq_12_bits_uop_fp_single;
  reg         ldq_12_bits_uop_xcpt_pf_if;
  reg         ldq_12_bits_uop_xcpt_ae_if;
  reg         ldq_12_bits_uop_xcpt_ma_if;
  reg         ldq_12_bits_uop_bp_debug_if;
  reg         ldq_12_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_12_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_12_bits_uop_debug_tsrc;
  reg         ldq_12_bits_addr_valid;
  reg  [39:0] ldq_12_bits_addr_bits;
  reg         ldq_12_bits_addr_is_virtual;
  reg         ldq_12_bits_addr_is_uncacheable;
  reg         ldq_12_bits_executed;
  reg         ldq_12_bits_succeeded;
  reg         ldq_12_bits_order_fail;
  reg         ldq_12_bits_observed;
  reg  [31:0] ldq_12_bits_st_dep_mask;
  reg  [4:0]  ldq_12_bits_youngest_stq_idx;
  reg         ldq_12_bits_forward_std_val;
  reg  [4:0]  ldq_12_bits_forward_stq_idx;
  reg         ldq_13_valid;
  reg  [6:0]  ldq_13_bits_uop_uopc;
  reg  [31:0] ldq_13_bits_uop_inst;
  reg  [31:0] ldq_13_bits_uop_debug_inst;
  reg         ldq_13_bits_uop_is_rvc;
  reg  [39:0] ldq_13_bits_uop_debug_pc;
  reg  [2:0]  ldq_13_bits_uop_iq_type;
  reg  [9:0]  ldq_13_bits_uop_fu_code;
  reg  [3:0]  ldq_13_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_13_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_13_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_13_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_13_bits_uop_ctrl_op_fcn;
  reg         ldq_13_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_13_bits_uop_ctrl_csr_cmd;
  reg         ldq_13_bits_uop_ctrl_is_load;
  reg         ldq_13_bits_uop_ctrl_is_sta;
  reg         ldq_13_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_13_bits_uop_iw_state;
  reg         ldq_13_bits_uop_iw_p1_poisoned;
  reg         ldq_13_bits_uop_iw_p2_poisoned;
  reg         ldq_13_bits_uop_is_br;
  reg         ldq_13_bits_uop_is_jalr;
  reg         ldq_13_bits_uop_is_jal;
  reg         ldq_13_bits_uop_is_sfb;
  reg  [19:0] ldq_13_bits_uop_br_mask;
  reg  [4:0]  ldq_13_bits_uop_br_tag;
  reg  [5:0]  ldq_13_bits_uop_ftq_idx;
  reg         ldq_13_bits_uop_edge_inst;
  reg  [5:0]  ldq_13_bits_uop_pc_lob;
  reg         ldq_13_bits_uop_taken;
  reg  [19:0] ldq_13_bits_uop_imm_packed;
  reg  [11:0] ldq_13_bits_uop_csr_addr;
  reg  [6:0]  ldq_13_bits_uop_rob_idx;
  reg  [4:0]  ldq_13_bits_uop_ldq_idx;
  reg  [4:0]  ldq_13_bits_uop_stq_idx;
  reg  [1:0]  ldq_13_bits_uop_rxq_idx;
  reg  [6:0]  ldq_13_bits_uop_pdst;
  reg  [6:0]  ldq_13_bits_uop_prs1;
  reg  [6:0]  ldq_13_bits_uop_prs2;
  reg  [6:0]  ldq_13_bits_uop_prs3;
  reg         ldq_13_bits_uop_prs1_busy;
  reg         ldq_13_bits_uop_prs2_busy;
  reg         ldq_13_bits_uop_prs3_busy;
  reg  [6:0]  ldq_13_bits_uop_stale_pdst;
  reg         ldq_13_bits_uop_exception;
  reg  [63:0] ldq_13_bits_uop_exc_cause;
  reg         ldq_13_bits_uop_bypassable;
  reg  [4:0]  ldq_13_bits_uop_mem_cmd;
  reg  [1:0]  ldq_13_bits_uop_mem_size;
  reg         ldq_13_bits_uop_mem_signed;
  reg         ldq_13_bits_uop_is_fence;
  reg         ldq_13_bits_uop_is_fencei;
  reg         ldq_13_bits_uop_is_amo;
  reg         ldq_13_bits_uop_uses_ldq;
  reg         ldq_13_bits_uop_uses_stq;
  reg         ldq_13_bits_uop_is_sys_pc2epc;
  reg         ldq_13_bits_uop_is_unique;
  reg         ldq_13_bits_uop_flush_on_commit;
  reg         ldq_13_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_13_bits_uop_ldst;
  reg  [5:0]  ldq_13_bits_uop_lrs1;
  reg  [5:0]  ldq_13_bits_uop_lrs2;
  reg  [5:0]  ldq_13_bits_uop_lrs3;
  reg         ldq_13_bits_uop_ldst_val;
  reg  [1:0]  ldq_13_bits_uop_dst_rtype;
  reg  [1:0]  ldq_13_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_13_bits_uop_lrs2_rtype;
  reg         ldq_13_bits_uop_frs3_en;
  reg         ldq_13_bits_uop_fp_val;
  reg         ldq_13_bits_uop_fp_single;
  reg         ldq_13_bits_uop_xcpt_pf_if;
  reg         ldq_13_bits_uop_xcpt_ae_if;
  reg         ldq_13_bits_uop_xcpt_ma_if;
  reg         ldq_13_bits_uop_bp_debug_if;
  reg         ldq_13_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_13_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_13_bits_uop_debug_tsrc;
  reg         ldq_13_bits_addr_valid;
  reg  [39:0] ldq_13_bits_addr_bits;
  reg         ldq_13_bits_addr_is_virtual;
  reg         ldq_13_bits_addr_is_uncacheable;
  reg         ldq_13_bits_executed;
  reg         ldq_13_bits_succeeded;
  reg         ldq_13_bits_order_fail;
  reg         ldq_13_bits_observed;
  reg  [31:0] ldq_13_bits_st_dep_mask;
  reg  [4:0]  ldq_13_bits_youngest_stq_idx;
  reg         ldq_13_bits_forward_std_val;
  reg  [4:0]  ldq_13_bits_forward_stq_idx;
  reg         ldq_14_valid;
  reg  [6:0]  ldq_14_bits_uop_uopc;
  reg  [31:0] ldq_14_bits_uop_inst;
  reg  [31:0] ldq_14_bits_uop_debug_inst;
  reg         ldq_14_bits_uop_is_rvc;
  reg  [39:0] ldq_14_bits_uop_debug_pc;
  reg  [2:0]  ldq_14_bits_uop_iq_type;
  reg  [9:0]  ldq_14_bits_uop_fu_code;
  reg  [3:0]  ldq_14_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_14_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_14_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_14_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_14_bits_uop_ctrl_op_fcn;
  reg         ldq_14_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_14_bits_uop_ctrl_csr_cmd;
  reg         ldq_14_bits_uop_ctrl_is_load;
  reg         ldq_14_bits_uop_ctrl_is_sta;
  reg         ldq_14_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_14_bits_uop_iw_state;
  reg         ldq_14_bits_uop_iw_p1_poisoned;
  reg         ldq_14_bits_uop_iw_p2_poisoned;
  reg         ldq_14_bits_uop_is_br;
  reg         ldq_14_bits_uop_is_jalr;
  reg         ldq_14_bits_uop_is_jal;
  reg         ldq_14_bits_uop_is_sfb;
  reg  [19:0] ldq_14_bits_uop_br_mask;
  reg  [4:0]  ldq_14_bits_uop_br_tag;
  reg  [5:0]  ldq_14_bits_uop_ftq_idx;
  reg         ldq_14_bits_uop_edge_inst;
  reg  [5:0]  ldq_14_bits_uop_pc_lob;
  reg         ldq_14_bits_uop_taken;
  reg  [19:0] ldq_14_bits_uop_imm_packed;
  reg  [11:0] ldq_14_bits_uop_csr_addr;
  reg  [6:0]  ldq_14_bits_uop_rob_idx;
  reg  [4:0]  ldq_14_bits_uop_ldq_idx;
  reg  [4:0]  ldq_14_bits_uop_stq_idx;
  reg  [1:0]  ldq_14_bits_uop_rxq_idx;
  reg  [6:0]  ldq_14_bits_uop_pdst;
  reg  [6:0]  ldq_14_bits_uop_prs1;
  reg  [6:0]  ldq_14_bits_uop_prs2;
  reg  [6:0]  ldq_14_bits_uop_prs3;
  reg         ldq_14_bits_uop_prs1_busy;
  reg         ldq_14_bits_uop_prs2_busy;
  reg         ldq_14_bits_uop_prs3_busy;
  reg  [6:0]  ldq_14_bits_uop_stale_pdst;
  reg         ldq_14_bits_uop_exception;
  reg  [63:0] ldq_14_bits_uop_exc_cause;
  reg         ldq_14_bits_uop_bypassable;
  reg  [4:0]  ldq_14_bits_uop_mem_cmd;
  reg  [1:0]  ldq_14_bits_uop_mem_size;
  reg         ldq_14_bits_uop_mem_signed;
  reg         ldq_14_bits_uop_is_fence;
  reg         ldq_14_bits_uop_is_fencei;
  reg         ldq_14_bits_uop_is_amo;
  reg         ldq_14_bits_uop_uses_ldq;
  reg         ldq_14_bits_uop_uses_stq;
  reg         ldq_14_bits_uop_is_sys_pc2epc;
  reg         ldq_14_bits_uop_is_unique;
  reg         ldq_14_bits_uop_flush_on_commit;
  reg         ldq_14_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_14_bits_uop_ldst;
  reg  [5:0]  ldq_14_bits_uop_lrs1;
  reg  [5:0]  ldq_14_bits_uop_lrs2;
  reg  [5:0]  ldq_14_bits_uop_lrs3;
  reg         ldq_14_bits_uop_ldst_val;
  reg  [1:0]  ldq_14_bits_uop_dst_rtype;
  reg  [1:0]  ldq_14_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_14_bits_uop_lrs2_rtype;
  reg         ldq_14_bits_uop_frs3_en;
  reg         ldq_14_bits_uop_fp_val;
  reg         ldq_14_bits_uop_fp_single;
  reg         ldq_14_bits_uop_xcpt_pf_if;
  reg         ldq_14_bits_uop_xcpt_ae_if;
  reg         ldq_14_bits_uop_xcpt_ma_if;
  reg         ldq_14_bits_uop_bp_debug_if;
  reg         ldq_14_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_14_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_14_bits_uop_debug_tsrc;
  reg         ldq_14_bits_addr_valid;
  reg  [39:0] ldq_14_bits_addr_bits;
  reg         ldq_14_bits_addr_is_virtual;
  reg         ldq_14_bits_addr_is_uncacheable;
  reg         ldq_14_bits_executed;
  reg         ldq_14_bits_succeeded;
  reg         ldq_14_bits_order_fail;
  reg         ldq_14_bits_observed;
  reg  [31:0] ldq_14_bits_st_dep_mask;
  reg  [4:0]  ldq_14_bits_youngest_stq_idx;
  reg         ldq_14_bits_forward_std_val;
  reg  [4:0]  ldq_14_bits_forward_stq_idx;
  reg         ldq_15_valid;
  reg  [6:0]  ldq_15_bits_uop_uopc;
  reg  [31:0] ldq_15_bits_uop_inst;
  reg  [31:0] ldq_15_bits_uop_debug_inst;
  reg         ldq_15_bits_uop_is_rvc;
  reg  [39:0] ldq_15_bits_uop_debug_pc;
  reg  [2:0]  ldq_15_bits_uop_iq_type;
  reg  [9:0]  ldq_15_bits_uop_fu_code;
  reg  [3:0]  ldq_15_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_15_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_15_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_15_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_15_bits_uop_ctrl_op_fcn;
  reg         ldq_15_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_15_bits_uop_ctrl_csr_cmd;
  reg         ldq_15_bits_uop_ctrl_is_load;
  reg         ldq_15_bits_uop_ctrl_is_sta;
  reg         ldq_15_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_15_bits_uop_iw_state;
  reg         ldq_15_bits_uop_iw_p1_poisoned;
  reg         ldq_15_bits_uop_iw_p2_poisoned;
  reg         ldq_15_bits_uop_is_br;
  reg         ldq_15_bits_uop_is_jalr;
  reg         ldq_15_bits_uop_is_jal;
  reg         ldq_15_bits_uop_is_sfb;
  reg  [19:0] ldq_15_bits_uop_br_mask;
  reg  [4:0]  ldq_15_bits_uop_br_tag;
  reg  [5:0]  ldq_15_bits_uop_ftq_idx;
  reg         ldq_15_bits_uop_edge_inst;
  reg  [5:0]  ldq_15_bits_uop_pc_lob;
  reg         ldq_15_bits_uop_taken;
  reg  [19:0] ldq_15_bits_uop_imm_packed;
  reg  [11:0] ldq_15_bits_uop_csr_addr;
  reg  [6:0]  ldq_15_bits_uop_rob_idx;
  reg  [4:0]  ldq_15_bits_uop_ldq_idx;
  reg  [4:0]  ldq_15_bits_uop_stq_idx;
  reg  [1:0]  ldq_15_bits_uop_rxq_idx;
  reg  [6:0]  ldq_15_bits_uop_pdst;
  reg  [6:0]  ldq_15_bits_uop_prs1;
  reg  [6:0]  ldq_15_bits_uop_prs2;
  reg  [6:0]  ldq_15_bits_uop_prs3;
  reg         ldq_15_bits_uop_prs1_busy;
  reg         ldq_15_bits_uop_prs2_busy;
  reg         ldq_15_bits_uop_prs3_busy;
  reg  [6:0]  ldq_15_bits_uop_stale_pdst;
  reg         ldq_15_bits_uop_exception;
  reg  [63:0] ldq_15_bits_uop_exc_cause;
  reg         ldq_15_bits_uop_bypassable;
  reg  [4:0]  ldq_15_bits_uop_mem_cmd;
  reg  [1:0]  ldq_15_bits_uop_mem_size;
  reg         ldq_15_bits_uop_mem_signed;
  reg         ldq_15_bits_uop_is_fence;
  reg         ldq_15_bits_uop_is_fencei;
  reg         ldq_15_bits_uop_is_amo;
  reg         ldq_15_bits_uop_uses_ldq;
  reg         ldq_15_bits_uop_uses_stq;
  reg         ldq_15_bits_uop_is_sys_pc2epc;
  reg         ldq_15_bits_uop_is_unique;
  reg         ldq_15_bits_uop_flush_on_commit;
  reg         ldq_15_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_15_bits_uop_ldst;
  reg  [5:0]  ldq_15_bits_uop_lrs1;
  reg  [5:0]  ldq_15_bits_uop_lrs2;
  reg  [5:0]  ldq_15_bits_uop_lrs3;
  reg         ldq_15_bits_uop_ldst_val;
  reg  [1:0]  ldq_15_bits_uop_dst_rtype;
  reg  [1:0]  ldq_15_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_15_bits_uop_lrs2_rtype;
  reg         ldq_15_bits_uop_frs3_en;
  reg         ldq_15_bits_uop_fp_val;
  reg         ldq_15_bits_uop_fp_single;
  reg         ldq_15_bits_uop_xcpt_pf_if;
  reg         ldq_15_bits_uop_xcpt_ae_if;
  reg         ldq_15_bits_uop_xcpt_ma_if;
  reg         ldq_15_bits_uop_bp_debug_if;
  reg         ldq_15_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_15_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_15_bits_uop_debug_tsrc;
  reg         ldq_15_bits_addr_valid;
  reg  [39:0] ldq_15_bits_addr_bits;
  reg         ldq_15_bits_addr_is_virtual;
  reg         ldq_15_bits_addr_is_uncacheable;
  reg         ldq_15_bits_executed;
  reg         ldq_15_bits_succeeded;
  reg         ldq_15_bits_order_fail;
  reg         ldq_15_bits_observed;
  reg  [31:0] ldq_15_bits_st_dep_mask;
  reg  [4:0]  ldq_15_bits_youngest_stq_idx;
  reg         ldq_15_bits_forward_std_val;
  reg  [4:0]  ldq_15_bits_forward_stq_idx;
  reg         ldq_16_valid;
  reg  [6:0]  ldq_16_bits_uop_uopc;
  reg  [31:0] ldq_16_bits_uop_inst;
  reg  [31:0] ldq_16_bits_uop_debug_inst;
  reg         ldq_16_bits_uop_is_rvc;
  reg  [39:0] ldq_16_bits_uop_debug_pc;
  reg  [2:0]  ldq_16_bits_uop_iq_type;
  reg  [9:0]  ldq_16_bits_uop_fu_code;
  reg  [3:0]  ldq_16_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_16_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_16_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_16_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_16_bits_uop_ctrl_op_fcn;
  reg         ldq_16_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_16_bits_uop_ctrl_csr_cmd;
  reg         ldq_16_bits_uop_ctrl_is_load;
  reg         ldq_16_bits_uop_ctrl_is_sta;
  reg         ldq_16_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_16_bits_uop_iw_state;
  reg         ldq_16_bits_uop_iw_p1_poisoned;
  reg         ldq_16_bits_uop_iw_p2_poisoned;
  reg         ldq_16_bits_uop_is_br;
  reg         ldq_16_bits_uop_is_jalr;
  reg         ldq_16_bits_uop_is_jal;
  reg         ldq_16_bits_uop_is_sfb;
  reg  [19:0] ldq_16_bits_uop_br_mask;
  reg  [4:0]  ldq_16_bits_uop_br_tag;
  reg  [5:0]  ldq_16_bits_uop_ftq_idx;
  reg         ldq_16_bits_uop_edge_inst;
  reg  [5:0]  ldq_16_bits_uop_pc_lob;
  reg         ldq_16_bits_uop_taken;
  reg  [19:0] ldq_16_bits_uop_imm_packed;
  reg  [11:0] ldq_16_bits_uop_csr_addr;
  reg  [6:0]  ldq_16_bits_uop_rob_idx;
  reg  [4:0]  ldq_16_bits_uop_ldq_idx;
  reg  [4:0]  ldq_16_bits_uop_stq_idx;
  reg  [1:0]  ldq_16_bits_uop_rxq_idx;
  reg  [6:0]  ldq_16_bits_uop_pdst;
  reg  [6:0]  ldq_16_bits_uop_prs1;
  reg  [6:0]  ldq_16_bits_uop_prs2;
  reg  [6:0]  ldq_16_bits_uop_prs3;
  reg         ldq_16_bits_uop_prs1_busy;
  reg         ldq_16_bits_uop_prs2_busy;
  reg         ldq_16_bits_uop_prs3_busy;
  reg  [6:0]  ldq_16_bits_uop_stale_pdst;
  reg         ldq_16_bits_uop_exception;
  reg  [63:0] ldq_16_bits_uop_exc_cause;
  reg         ldq_16_bits_uop_bypassable;
  reg  [4:0]  ldq_16_bits_uop_mem_cmd;
  reg  [1:0]  ldq_16_bits_uop_mem_size;
  reg         ldq_16_bits_uop_mem_signed;
  reg         ldq_16_bits_uop_is_fence;
  reg         ldq_16_bits_uop_is_fencei;
  reg         ldq_16_bits_uop_is_amo;
  reg         ldq_16_bits_uop_uses_ldq;
  reg         ldq_16_bits_uop_uses_stq;
  reg         ldq_16_bits_uop_is_sys_pc2epc;
  reg         ldq_16_bits_uop_is_unique;
  reg         ldq_16_bits_uop_flush_on_commit;
  reg         ldq_16_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_16_bits_uop_ldst;
  reg  [5:0]  ldq_16_bits_uop_lrs1;
  reg  [5:0]  ldq_16_bits_uop_lrs2;
  reg  [5:0]  ldq_16_bits_uop_lrs3;
  reg         ldq_16_bits_uop_ldst_val;
  reg  [1:0]  ldq_16_bits_uop_dst_rtype;
  reg  [1:0]  ldq_16_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_16_bits_uop_lrs2_rtype;
  reg         ldq_16_bits_uop_frs3_en;
  reg         ldq_16_bits_uop_fp_val;
  reg         ldq_16_bits_uop_fp_single;
  reg         ldq_16_bits_uop_xcpt_pf_if;
  reg         ldq_16_bits_uop_xcpt_ae_if;
  reg         ldq_16_bits_uop_xcpt_ma_if;
  reg         ldq_16_bits_uop_bp_debug_if;
  reg         ldq_16_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_16_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_16_bits_uop_debug_tsrc;
  reg         ldq_16_bits_addr_valid;
  reg  [39:0] ldq_16_bits_addr_bits;
  reg         ldq_16_bits_addr_is_virtual;
  reg         ldq_16_bits_addr_is_uncacheable;
  reg         ldq_16_bits_executed;
  reg         ldq_16_bits_succeeded;
  reg         ldq_16_bits_order_fail;
  reg         ldq_16_bits_observed;
  reg  [31:0] ldq_16_bits_st_dep_mask;
  reg  [4:0]  ldq_16_bits_youngest_stq_idx;
  reg         ldq_16_bits_forward_std_val;
  reg  [4:0]  ldq_16_bits_forward_stq_idx;
  reg         ldq_17_valid;
  reg  [6:0]  ldq_17_bits_uop_uopc;
  reg  [31:0] ldq_17_bits_uop_inst;
  reg  [31:0] ldq_17_bits_uop_debug_inst;
  reg         ldq_17_bits_uop_is_rvc;
  reg  [39:0] ldq_17_bits_uop_debug_pc;
  reg  [2:0]  ldq_17_bits_uop_iq_type;
  reg  [9:0]  ldq_17_bits_uop_fu_code;
  reg  [3:0]  ldq_17_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_17_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_17_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_17_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_17_bits_uop_ctrl_op_fcn;
  reg         ldq_17_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_17_bits_uop_ctrl_csr_cmd;
  reg         ldq_17_bits_uop_ctrl_is_load;
  reg         ldq_17_bits_uop_ctrl_is_sta;
  reg         ldq_17_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_17_bits_uop_iw_state;
  reg         ldq_17_bits_uop_iw_p1_poisoned;
  reg         ldq_17_bits_uop_iw_p2_poisoned;
  reg         ldq_17_bits_uop_is_br;
  reg         ldq_17_bits_uop_is_jalr;
  reg         ldq_17_bits_uop_is_jal;
  reg         ldq_17_bits_uop_is_sfb;
  reg  [19:0] ldq_17_bits_uop_br_mask;
  reg  [4:0]  ldq_17_bits_uop_br_tag;
  reg  [5:0]  ldq_17_bits_uop_ftq_idx;
  reg         ldq_17_bits_uop_edge_inst;
  reg  [5:0]  ldq_17_bits_uop_pc_lob;
  reg         ldq_17_bits_uop_taken;
  reg  [19:0] ldq_17_bits_uop_imm_packed;
  reg  [11:0] ldq_17_bits_uop_csr_addr;
  reg  [6:0]  ldq_17_bits_uop_rob_idx;
  reg  [4:0]  ldq_17_bits_uop_ldq_idx;
  reg  [4:0]  ldq_17_bits_uop_stq_idx;
  reg  [1:0]  ldq_17_bits_uop_rxq_idx;
  reg  [6:0]  ldq_17_bits_uop_pdst;
  reg  [6:0]  ldq_17_bits_uop_prs1;
  reg  [6:0]  ldq_17_bits_uop_prs2;
  reg  [6:0]  ldq_17_bits_uop_prs3;
  reg         ldq_17_bits_uop_prs1_busy;
  reg         ldq_17_bits_uop_prs2_busy;
  reg         ldq_17_bits_uop_prs3_busy;
  reg  [6:0]  ldq_17_bits_uop_stale_pdst;
  reg         ldq_17_bits_uop_exception;
  reg  [63:0] ldq_17_bits_uop_exc_cause;
  reg         ldq_17_bits_uop_bypassable;
  reg  [4:0]  ldq_17_bits_uop_mem_cmd;
  reg  [1:0]  ldq_17_bits_uop_mem_size;
  reg         ldq_17_bits_uop_mem_signed;
  reg         ldq_17_bits_uop_is_fence;
  reg         ldq_17_bits_uop_is_fencei;
  reg         ldq_17_bits_uop_is_amo;
  reg         ldq_17_bits_uop_uses_ldq;
  reg         ldq_17_bits_uop_uses_stq;
  reg         ldq_17_bits_uop_is_sys_pc2epc;
  reg         ldq_17_bits_uop_is_unique;
  reg         ldq_17_bits_uop_flush_on_commit;
  reg         ldq_17_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_17_bits_uop_ldst;
  reg  [5:0]  ldq_17_bits_uop_lrs1;
  reg  [5:0]  ldq_17_bits_uop_lrs2;
  reg  [5:0]  ldq_17_bits_uop_lrs3;
  reg         ldq_17_bits_uop_ldst_val;
  reg  [1:0]  ldq_17_bits_uop_dst_rtype;
  reg  [1:0]  ldq_17_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_17_bits_uop_lrs2_rtype;
  reg         ldq_17_bits_uop_frs3_en;
  reg         ldq_17_bits_uop_fp_val;
  reg         ldq_17_bits_uop_fp_single;
  reg         ldq_17_bits_uop_xcpt_pf_if;
  reg         ldq_17_bits_uop_xcpt_ae_if;
  reg         ldq_17_bits_uop_xcpt_ma_if;
  reg         ldq_17_bits_uop_bp_debug_if;
  reg         ldq_17_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_17_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_17_bits_uop_debug_tsrc;
  reg         ldq_17_bits_addr_valid;
  reg  [39:0] ldq_17_bits_addr_bits;
  reg         ldq_17_bits_addr_is_virtual;
  reg         ldq_17_bits_addr_is_uncacheable;
  reg         ldq_17_bits_executed;
  reg         ldq_17_bits_succeeded;
  reg         ldq_17_bits_order_fail;
  reg         ldq_17_bits_observed;
  reg  [31:0] ldq_17_bits_st_dep_mask;
  reg  [4:0]  ldq_17_bits_youngest_stq_idx;
  reg         ldq_17_bits_forward_std_val;
  reg  [4:0]  ldq_17_bits_forward_stq_idx;
  reg         ldq_18_valid;
  reg  [6:0]  ldq_18_bits_uop_uopc;
  reg  [31:0] ldq_18_bits_uop_inst;
  reg  [31:0] ldq_18_bits_uop_debug_inst;
  reg         ldq_18_bits_uop_is_rvc;
  reg  [39:0] ldq_18_bits_uop_debug_pc;
  reg  [2:0]  ldq_18_bits_uop_iq_type;
  reg  [9:0]  ldq_18_bits_uop_fu_code;
  reg  [3:0]  ldq_18_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_18_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_18_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_18_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_18_bits_uop_ctrl_op_fcn;
  reg         ldq_18_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_18_bits_uop_ctrl_csr_cmd;
  reg         ldq_18_bits_uop_ctrl_is_load;
  reg         ldq_18_bits_uop_ctrl_is_sta;
  reg         ldq_18_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_18_bits_uop_iw_state;
  reg         ldq_18_bits_uop_iw_p1_poisoned;
  reg         ldq_18_bits_uop_iw_p2_poisoned;
  reg         ldq_18_bits_uop_is_br;
  reg         ldq_18_bits_uop_is_jalr;
  reg         ldq_18_bits_uop_is_jal;
  reg         ldq_18_bits_uop_is_sfb;
  reg  [19:0] ldq_18_bits_uop_br_mask;
  reg  [4:0]  ldq_18_bits_uop_br_tag;
  reg  [5:0]  ldq_18_bits_uop_ftq_idx;
  reg         ldq_18_bits_uop_edge_inst;
  reg  [5:0]  ldq_18_bits_uop_pc_lob;
  reg         ldq_18_bits_uop_taken;
  reg  [19:0] ldq_18_bits_uop_imm_packed;
  reg  [11:0] ldq_18_bits_uop_csr_addr;
  reg  [6:0]  ldq_18_bits_uop_rob_idx;
  reg  [4:0]  ldq_18_bits_uop_ldq_idx;
  reg  [4:0]  ldq_18_bits_uop_stq_idx;
  reg  [1:0]  ldq_18_bits_uop_rxq_idx;
  reg  [6:0]  ldq_18_bits_uop_pdst;
  reg  [6:0]  ldq_18_bits_uop_prs1;
  reg  [6:0]  ldq_18_bits_uop_prs2;
  reg  [6:0]  ldq_18_bits_uop_prs3;
  reg         ldq_18_bits_uop_prs1_busy;
  reg         ldq_18_bits_uop_prs2_busy;
  reg         ldq_18_bits_uop_prs3_busy;
  reg  [6:0]  ldq_18_bits_uop_stale_pdst;
  reg         ldq_18_bits_uop_exception;
  reg  [63:0] ldq_18_bits_uop_exc_cause;
  reg         ldq_18_bits_uop_bypassable;
  reg  [4:0]  ldq_18_bits_uop_mem_cmd;
  reg  [1:0]  ldq_18_bits_uop_mem_size;
  reg         ldq_18_bits_uop_mem_signed;
  reg         ldq_18_bits_uop_is_fence;
  reg         ldq_18_bits_uop_is_fencei;
  reg         ldq_18_bits_uop_is_amo;
  reg         ldq_18_bits_uop_uses_ldq;
  reg         ldq_18_bits_uop_uses_stq;
  reg         ldq_18_bits_uop_is_sys_pc2epc;
  reg         ldq_18_bits_uop_is_unique;
  reg         ldq_18_bits_uop_flush_on_commit;
  reg         ldq_18_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_18_bits_uop_ldst;
  reg  [5:0]  ldq_18_bits_uop_lrs1;
  reg  [5:0]  ldq_18_bits_uop_lrs2;
  reg  [5:0]  ldq_18_bits_uop_lrs3;
  reg         ldq_18_bits_uop_ldst_val;
  reg  [1:0]  ldq_18_bits_uop_dst_rtype;
  reg  [1:0]  ldq_18_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_18_bits_uop_lrs2_rtype;
  reg         ldq_18_bits_uop_frs3_en;
  reg         ldq_18_bits_uop_fp_val;
  reg         ldq_18_bits_uop_fp_single;
  reg         ldq_18_bits_uop_xcpt_pf_if;
  reg         ldq_18_bits_uop_xcpt_ae_if;
  reg         ldq_18_bits_uop_xcpt_ma_if;
  reg         ldq_18_bits_uop_bp_debug_if;
  reg         ldq_18_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_18_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_18_bits_uop_debug_tsrc;
  reg         ldq_18_bits_addr_valid;
  reg  [39:0] ldq_18_bits_addr_bits;
  reg         ldq_18_bits_addr_is_virtual;
  reg         ldq_18_bits_addr_is_uncacheable;
  reg         ldq_18_bits_executed;
  reg         ldq_18_bits_succeeded;
  reg         ldq_18_bits_order_fail;
  reg         ldq_18_bits_observed;
  reg  [31:0] ldq_18_bits_st_dep_mask;
  reg  [4:0]  ldq_18_bits_youngest_stq_idx;
  reg         ldq_18_bits_forward_std_val;
  reg  [4:0]  ldq_18_bits_forward_stq_idx;
  reg         ldq_19_valid;
  reg  [6:0]  ldq_19_bits_uop_uopc;
  reg  [31:0] ldq_19_bits_uop_inst;
  reg  [31:0] ldq_19_bits_uop_debug_inst;
  reg         ldq_19_bits_uop_is_rvc;
  reg  [39:0] ldq_19_bits_uop_debug_pc;
  reg  [2:0]  ldq_19_bits_uop_iq_type;
  reg  [9:0]  ldq_19_bits_uop_fu_code;
  reg  [3:0]  ldq_19_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_19_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_19_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_19_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_19_bits_uop_ctrl_op_fcn;
  reg         ldq_19_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_19_bits_uop_ctrl_csr_cmd;
  reg         ldq_19_bits_uop_ctrl_is_load;
  reg         ldq_19_bits_uop_ctrl_is_sta;
  reg         ldq_19_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_19_bits_uop_iw_state;
  reg         ldq_19_bits_uop_iw_p1_poisoned;
  reg         ldq_19_bits_uop_iw_p2_poisoned;
  reg         ldq_19_bits_uop_is_br;
  reg         ldq_19_bits_uop_is_jalr;
  reg         ldq_19_bits_uop_is_jal;
  reg         ldq_19_bits_uop_is_sfb;
  reg  [19:0] ldq_19_bits_uop_br_mask;
  reg  [4:0]  ldq_19_bits_uop_br_tag;
  reg  [5:0]  ldq_19_bits_uop_ftq_idx;
  reg         ldq_19_bits_uop_edge_inst;
  reg  [5:0]  ldq_19_bits_uop_pc_lob;
  reg         ldq_19_bits_uop_taken;
  reg  [19:0] ldq_19_bits_uop_imm_packed;
  reg  [11:0] ldq_19_bits_uop_csr_addr;
  reg  [6:0]  ldq_19_bits_uop_rob_idx;
  reg  [4:0]  ldq_19_bits_uop_ldq_idx;
  reg  [4:0]  ldq_19_bits_uop_stq_idx;
  reg  [1:0]  ldq_19_bits_uop_rxq_idx;
  reg  [6:0]  ldq_19_bits_uop_pdst;
  reg  [6:0]  ldq_19_bits_uop_prs1;
  reg  [6:0]  ldq_19_bits_uop_prs2;
  reg  [6:0]  ldq_19_bits_uop_prs3;
  reg         ldq_19_bits_uop_prs1_busy;
  reg         ldq_19_bits_uop_prs2_busy;
  reg         ldq_19_bits_uop_prs3_busy;
  reg  [6:0]  ldq_19_bits_uop_stale_pdst;
  reg         ldq_19_bits_uop_exception;
  reg  [63:0] ldq_19_bits_uop_exc_cause;
  reg         ldq_19_bits_uop_bypassable;
  reg  [4:0]  ldq_19_bits_uop_mem_cmd;
  reg  [1:0]  ldq_19_bits_uop_mem_size;
  reg         ldq_19_bits_uop_mem_signed;
  reg         ldq_19_bits_uop_is_fence;
  reg         ldq_19_bits_uop_is_fencei;
  reg         ldq_19_bits_uop_is_amo;
  reg         ldq_19_bits_uop_uses_ldq;
  reg         ldq_19_bits_uop_uses_stq;
  reg         ldq_19_bits_uop_is_sys_pc2epc;
  reg         ldq_19_bits_uop_is_unique;
  reg         ldq_19_bits_uop_flush_on_commit;
  reg         ldq_19_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_19_bits_uop_ldst;
  reg  [5:0]  ldq_19_bits_uop_lrs1;
  reg  [5:0]  ldq_19_bits_uop_lrs2;
  reg  [5:0]  ldq_19_bits_uop_lrs3;
  reg         ldq_19_bits_uop_ldst_val;
  reg  [1:0]  ldq_19_bits_uop_dst_rtype;
  reg  [1:0]  ldq_19_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_19_bits_uop_lrs2_rtype;
  reg         ldq_19_bits_uop_frs3_en;
  reg         ldq_19_bits_uop_fp_val;
  reg         ldq_19_bits_uop_fp_single;
  reg         ldq_19_bits_uop_xcpt_pf_if;
  reg         ldq_19_bits_uop_xcpt_ae_if;
  reg         ldq_19_bits_uop_xcpt_ma_if;
  reg         ldq_19_bits_uop_bp_debug_if;
  reg         ldq_19_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_19_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_19_bits_uop_debug_tsrc;
  reg         ldq_19_bits_addr_valid;
  reg  [39:0] ldq_19_bits_addr_bits;
  reg         ldq_19_bits_addr_is_virtual;
  reg         ldq_19_bits_addr_is_uncacheable;
  reg         ldq_19_bits_executed;
  reg         ldq_19_bits_succeeded;
  reg         ldq_19_bits_order_fail;
  reg         ldq_19_bits_observed;
  reg  [31:0] ldq_19_bits_st_dep_mask;
  reg  [4:0]  ldq_19_bits_youngest_stq_idx;
  reg         ldq_19_bits_forward_std_val;
  reg  [4:0]  ldq_19_bits_forward_stq_idx;
  reg         ldq_20_valid;
  reg  [6:0]  ldq_20_bits_uop_uopc;
  reg  [31:0] ldq_20_bits_uop_inst;
  reg  [31:0] ldq_20_bits_uop_debug_inst;
  reg         ldq_20_bits_uop_is_rvc;
  reg  [39:0] ldq_20_bits_uop_debug_pc;
  reg  [2:0]  ldq_20_bits_uop_iq_type;
  reg  [9:0]  ldq_20_bits_uop_fu_code;
  reg  [3:0]  ldq_20_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_20_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_20_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_20_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_20_bits_uop_ctrl_op_fcn;
  reg         ldq_20_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_20_bits_uop_ctrl_csr_cmd;
  reg         ldq_20_bits_uop_ctrl_is_load;
  reg         ldq_20_bits_uop_ctrl_is_sta;
  reg         ldq_20_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_20_bits_uop_iw_state;
  reg         ldq_20_bits_uop_iw_p1_poisoned;
  reg         ldq_20_bits_uop_iw_p2_poisoned;
  reg         ldq_20_bits_uop_is_br;
  reg         ldq_20_bits_uop_is_jalr;
  reg         ldq_20_bits_uop_is_jal;
  reg         ldq_20_bits_uop_is_sfb;
  reg  [19:0] ldq_20_bits_uop_br_mask;
  reg  [4:0]  ldq_20_bits_uop_br_tag;
  reg  [5:0]  ldq_20_bits_uop_ftq_idx;
  reg         ldq_20_bits_uop_edge_inst;
  reg  [5:0]  ldq_20_bits_uop_pc_lob;
  reg         ldq_20_bits_uop_taken;
  reg  [19:0] ldq_20_bits_uop_imm_packed;
  reg  [11:0] ldq_20_bits_uop_csr_addr;
  reg  [6:0]  ldq_20_bits_uop_rob_idx;
  reg  [4:0]  ldq_20_bits_uop_ldq_idx;
  reg  [4:0]  ldq_20_bits_uop_stq_idx;
  reg  [1:0]  ldq_20_bits_uop_rxq_idx;
  reg  [6:0]  ldq_20_bits_uop_pdst;
  reg  [6:0]  ldq_20_bits_uop_prs1;
  reg  [6:0]  ldq_20_bits_uop_prs2;
  reg  [6:0]  ldq_20_bits_uop_prs3;
  reg         ldq_20_bits_uop_prs1_busy;
  reg         ldq_20_bits_uop_prs2_busy;
  reg         ldq_20_bits_uop_prs3_busy;
  reg  [6:0]  ldq_20_bits_uop_stale_pdst;
  reg         ldq_20_bits_uop_exception;
  reg  [63:0] ldq_20_bits_uop_exc_cause;
  reg         ldq_20_bits_uop_bypassable;
  reg  [4:0]  ldq_20_bits_uop_mem_cmd;
  reg  [1:0]  ldq_20_bits_uop_mem_size;
  reg         ldq_20_bits_uop_mem_signed;
  reg         ldq_20_bits_uop_is_fence;
  reg         ldq_20_bits_uop_is_fencei;
  reg         ldq_20_bits_uop_is_amo;
  reg         ldq_20_bits_uop_uses_ldq;
  reg         ldq_20_bits_uop_uses_stq;
  reg         ldq_20_bits_uop_is_sys_pc2epc;
  reg         ldq_20_bits_uop_is_unique;
  reg         ldq_20_bits_uop_flush_on_commit;
  reg         ldq_20_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_20_bits_uop_ldst;
  reg  [5:0]  ldq_20_bits_uop_lrs1;
  reg  [5:0]  ldq_20_bits_uop_lrs2;
  reg  [5:0]  ldq_20_bits_uop_lrs3;
  reg         ldq_20_bits_uop_ldst_val;
  reg  [1:0]  ldq_20_bits_uop_dst_rtype;
  reg  [1:0]  ldq_20_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_20_bits_uop_lrs2_rtype;
  reg         ldq_20_bits_uop_frs3_en;
  reg         ldq_20_bits_uop_fp_val;
  reg         ldq_20_bits_uop_fp_single;
  reg         ldq_20_bits_uop_xcpt_pf_if;
  reg         ldq_20_bits_uop_xcpt_ae_if;
  reg         ldq_20_bits_uop_xcpt_ma_if;
  reg         ldq_20_bits_uop_bp_debug_if;
  reg         ldq_20_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_20_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_20_bits_uop_debug_tsrc;
  reg         ldq_20_bits_addr_valid;
  reg  [39:0] ldq_20_bits_addr_bits;
  reg         ldq_20_bits_addr_is_virtual;
  reg         ldq_20_bits_addr_is_uncacheable;
  reg         ldq_20_bits_executed;
  reg         ldq_20_bits_succeeded;
  reg         ldq_20_bits_order_fail;
  reg         ldq_20_bits_observed;
  reg  [31:0] ldq_20_bits_st_dep_mask;
  reg  [4:0]  ldq_20_bits_youngest_stq_idx;
  reg         ldq_20_bits_forward_std_val;
  reg  [4:0]  ldq_20_bits_forward_stq_idx;
  reg         ldq_21_valid;
  reg  [6:0]  ldq_21_bits_uop_uopc;
  reg  [31:0] ldq_21_bits_uop_inst;
  reg  [31:0] ldq_21_bits_uop_debug_inst;
  reg         ldq_21_bits_uop_is_rvc;
  reg  [39:0] ldq_21_bits_uop_debug_pc;
  reg  [2:0]  ldq_21_bits_uop_iq_type;
  reg  [9:0]  ldq_21_bits_uop_fu_code;
  reg  [3:0]  ldq_21_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_21_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_21_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_21_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_21_bits_uop_ctrl_op_fcn;
  reg         ldq_21_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_21_bits_uop_ctrl_csr_cmd;
  reg         ldq_21_bits_uop_ctrl_is_load;
  reg         ldq_21_bits_uop_ctrl_is_sta;
  reg         ldq_21_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_21_bits_uop_iw_state;
  reg         ldq_21_bits_uop_iw_p1_poisoned;
  reg         ldq_21_bits_uop_iw_p2_poisoned;
  reg         ldq_21_bits_uop_is_br;
  reg         ldq_21_bits_uop_is_jalr;
  reg         ldq_21_bits_uop_is_jal;
  reg         ldq_21_bits_uop_is_sfb;
  reg  [19:0] ldq_21_bits_uop_br_mask;
  reg  [4:0]  ldq_21_bits_uop_br_tag;
  reg  [5:0]  ldq_21_bits_uop_ftq_idx;
  reg         ldq_21_bits_uop_edge_inst;
  reg  [5:0]  ldq_21_bits_uop_pc_lob;
  reg         ldq_21_bits_uop_taken;
  reg  [19:0] ldq_21_bits_uop_imm_packed;
  reg  [11:0] ldq_21_bits_uop_csr_addr;
  reg  [6:0]  ldq_21_bits_uop_rob_idx;
  reg  [4:0]  ldq_21_bits_uop_ldq_idx;
  reg  [4:0]  ldq_21_bits_uop_stq_idx;
  reg  [1:0]  ldq_21_bits_uop_rxq_idx;
  reg  [6:0]  ldq_21_bits_uop_pdst;
  reg  [6:0]  ldq_21_bits_uop_prs1;
  reg  [6:0]  ldq_21_bits_uop_prs2;
  reg  [6:0]  ldq_21_bits_uop_prs3;
  reg         ldq_21_bits_uop_prs1_busy;
  reg         ldq_21_bits_uop_prs2_busy;
  reg         ldq_21_bits_uop_prs3_busy;
  reg  [6:0]  ldq_21_bits_uop_stale_pdst;
  reg         ldq_21_bits_uop_exception;
  reg  [63:0] ldq_21_bits_uop_exc_cause;
  reg         ldq_21_bits_uop_bypassable;
  reg  [4:0]  ldq_21_bits_uop_mem_cmd;
  reg  [1:0]  ldq_21_bits_uop_mem_size;
  reg         ldq_21_bits_uop_mem_signed;
  reg         ldq_21_bits_uop_is_fence;
  reg         ldq_21_bits_uop_is_fencei;
  reg         ldq_21_bits_uop_is_amo;
  reg         ldq_21_bits_uop_uses_ldq;
  reg         ldq_21_bits_uop_uses_stq;
  reg         ldq_21_bits_uop_is_sys_pc2epc;
  reg         ldq_21_bits_uop_is_unique;
  reg         ldq_21_bits_uop_flush_on_commit;
  reg         ldq_21_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_21_bits_uop_ldst;
  reg  [5:0]  ldq_21_bits_uop_lrs1;
  reg  [5:0]  ldq_21_bits_uop_lrs2;
  reg  [5:0]  ldq_21_bits_uop_lrs3;
  reg         ldq_21_bits_uop_ldst_val;
  reg  [1:0]  ldq_21_bits_uop_dst_rtype;
  reg  [1:0]  ldq_21_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_21_bits_uop_lrs2_rtype;
  reg         ldq_21_bits_uop_frs3_en;
  reg         ldq_21_bits_uop_fp_val;
  reg         ldq_21_bits_uop_fp_single;
  reg         ldq_21_bits_uop_xcpt_pf_if;
  reg         ldq_21_bits_uop_xcpt_ae_if;
  reg         ldq_21_bits_uop_xcpt_ma_if;
  reg         ldq_21_bits_uop_bp_debug_if;
  reg         ldq_21_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_21_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_21_bits_uop_debug_tsrc;
  reg         ldq_21_bits_addr_valid;
  reg  [39:0] ldq_21_bits_addr_bits;
  reg         ldq_21_bits_addr_is_virtual;
  reg         ldq_21_bits_addr_is_uncacheable;
  reg         ldq_21_bits_executed;
  reg         ldq_21_bits_succeeded;
  reg         ldq_21_bits_order_fail;
  reg         ldq_21_bits_observed;
  reg  [31:0] ldq_21_bits_st_dep_mask;
  reg  [4:0]  ldq_21_bits_youngest_stq_idx;
  reg         ldq_21_bits_forward_std_val;
  reg  [4:0]  ldq_21_bits_forward_stq_idx;
  reg         ldq_22_valid;
  reg  [6:0]  ldq_22_bits_uop_uopc;
  reg  [31:0] ldq_22_bits_uop_inst;
  reg  [31:0] ldq_22_bits_uop_debug_inst;
  reg         ldq_22_bits_uop_is_rvc;
  reg  [39:0] ldq_22_bits_uop_debug_pc;
  reg  [2:0]  ldq_22_bits_uop_iq_type;
  reg  [9:0]  ldq_22_bits_uop_fu_code;
  reg  [3:0]  ldq_22_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_22_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_22_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_22_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_22_bits_uop_ctrl_op_fcn;
  reg         ldq_22_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_22_bits_uop_ctrl_csr_cmd;
  reg         ldq_22_bits_uop_ctrl_is_load;
  reg         ldq_22_bits_uop_ctrl_is_sta;
  reg         ldq_22_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_22_bits_uop_iw_state;
  reg         ldq_22_bits_uop_iw_p1_poisoned;
  reg         ldq_22_bits_uop_iw_p2_poisoned;
  reg         ldq_22_bits_uop_is_br;
  reg         ldq_22_bits_uop_is_jalr;
  reg         ldq_22_bits_uop_is_jal;
  reg         ldq_22_bits_uop_is_sfb;
  reg  [19:0] ldq_22_bits_uop_br_mask;
  reg  [4:0]  ldq_22_bits_uop_br_tag;
  reg  [5:0]  ldq_22_bits_uop_ftq_idx;
  reg         ldq_22_bits_uop_edge_inst;
  reg  [5:0]  ldq_22_bits_uop_pc_lob;
  reg         ldq_22_bits_uop_taken;
  reg  [19:0] ldq_22_bits_uop_imm_packed;
  reg  [11:0] ldq_22_bits_uop_csr_addr;
  reg  [6:0]  ldq_22_bits_uop_rob_idx;
  reg  [4:0]  ldq_22_bits_uop_ldq_idx;
  reg  [4:0]  ldq_22_bits_uop_stq_idx;
  reg  [1:0]  ldq_22_bits_uop_rxq_idx;
  reg  [6:0]  ldq_22_bits_uop_pdst;
  reg  [6:0]  ldq_22_bits_uop_prs1;
  reg  [6:0]  ldq_22_bits_uop_prs2;
  reg  [6:0]  ldq_22_bits_uop_prs3;
  reg         ldq_22_bits_uop_prs1_busy;
  reg         ldq_22_bits_uop_prs2_busy;
  reg         ldq_22_bits_uop_prs3_busy;
  reg  [6:0]  ldq_22_bits_uop_stale_pdst;
  reg         ldq_22_bits_uop_exception;
  reg  [63:0] ldq_22_bits_uop_exc_cause;
  reg         ldq_22_bits_uop_bypassable;
  reg  [4:0]  ldq_22_bits_uop_mem_cmd;
  reg  [1:0]  ldq_22_bits_uop_mem_size;
  reg         ldq_22_bits_uop_mem_signed;
  reg         ldq_22_bits_uop_is_fence;
  reg         ldq_22_bits_uop_is_fencei;
  reg         ldq_22_bits_uop_is_amo;
  reg         ldq_22_bits_uop_uses_ldq;
  reg         ldq_22_bits_uop_uses_stq;
  reg         ldq_22_bits_uop_is_sys_pc2epc;
  reg         ldq_22_bits_uop_is_unique;
  reg         ldq_22_bits_uop_flush_on_commit;
  reg         ldq_22_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_22_bits_uop_ldst;
  reg  [5:0]  ldq_22_bits_uop_lrs1;
  reg  [5:0]  ldq_22_bits_uop_lrs2;
  reg  [5:0]  ldq_22_bits_uop_lrs3;
  reg         ldq_22_bits_uop_ldst_val;
  reg  [1:0]  ldq_22_bits_uop_dst_rtype;
  reg  [1:0]  ldq_22_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_22_bits_uop_lrs2_rtype;
  reg         ldq_22_bits_uop_frs3_en;
  reg         ldq_22_bits_uop_fp_val;
  reg         ldq_22_bits_uop_fp_single;
  reg         ldq_22_bits_uop_xcpt_pf_if;
  reg         ldq_22_bits_uop_xcpt_ae_if;
  reg         ldq_22_bits_uop_xcpt_ma_if;
  reg         ldq_22_bits_uop_bp_debug_if;
  reg         ldq_22_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_22_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_22_bits_uop_debug_tsrc;
  reg         ldq_22_bits_addr_valid;
  reg  [39:0] ldq_22_bits_addr_bits;
  reg         ldq_22_bits_addr_is_virtual;
  reg         ldq_22_bits_addr_is_uncacheable;
  reg         ldq_22_bits_executed;
  reg         ldq_22_bits_succeeded;
  reg         ldq_22_bits_order_fail;
  reg         ldq_22_bits_observed;
  reg  [31:0] ldq_22_bits_st_dep_mask;
  reg  [4:0]  ldq_22_bits_youngest_stq_idx;
  reg         ldq_22_bits_forward_std_val;
  reg  [4:0]  ldq_22_bits_forward_stq_idx;
  reg         ldq_23_valid;
  reg  [6:0]  ldq_23_bits_uop_uopc;
  reg  [31:0] ldq_23_bits_uop_inst;
  reg  [31:0] ldq_23_bits_uop_debug_inst;
  reg         ldq_23_bits_uop_is_rvc;
  reg  [39:0] ldq_23_bits_uop_debug_pc;
  reg  [2:0]  ldq_23_bits_uop_iq_type;
  reg  [9:0]  ldq_23_bits_uop_fu_code;
  reg  [3:0]  ldq_23_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_23_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_23_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_23_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_23_bits_uop_ctrl_op_fcn;
  reg         ldq_23_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_23_bits_uop_ctrl_csr_cmd;
  reg         ldq_23_bits_uop_ctrl_is_load;
  reg         ldq_23_bits_uop_ctrl_is_sta;
  reg         ldq_23_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_23_bits_uop_iw_state;
  reg         ldq_23_bits_uop_iw_p1_poisoned;
  reg         ldq_23_bits_uop_iw_p2_poisoned;
  reg         ldq_23_bits_uop_is_br;
  reg         ldq_23_bits_uop_is_jalr;
  reg         ldq_23_bits_uop_is_jal;
  reg         ldq_23_bits_uop_is_sfb;
  reg  [19:0] ldq_23_bits_uop_br_mask;
  reg  [4:0]  ldq_23_bits_uop_br_tag;
  reg  [5:0]  ldq_23_bits_uop_ftq_idx;
  reg         ldq_23_bits_uop_edge_inst;
  reg  [5:0]  ldq_23_bits_uop_pc_lob;
  reg         ldq_23_bits_uop_taken;
  reg  [19:0] ldq_23_bits_uop_imm_packed;
  reg  [11:0] ldq_23_bits_uop_csr_addr;
  reg  [6:0]  ldq_23_bits_uop_rob_idx;
  reg  [4:0]  ldq_23_bits_uop_ldq_idx;
  reg  [4:0]  ldq_23_bits_uop_stq_idx;
  reg  [1:0]  ldq_23_bits_uop_rxq_idx;
  reg  [6:0]  ldq_23_bits_uop_pdst;
  reg  [6:0]  ldq_23_bits_uop_prs1;
  reg  [6:0]  ldq_23_bits_uop_prs2;
  reg  [6:0]  ldq_23_bits_uop_prs3;
  reg         ldq_23_bits_uop_prs1_busy;
  reg         ldq_23_bits_uop_prs2_busy;
  reg         ldq_23_bits_uop_prs3_busy;
  reg  [6:0]  ldq_23_bits_uop_stale_pdst;
  reg         ldq_23_bits_uop_exception;
  reg  [63:0] ldq_23_bits_uop_exc_cause;
  reg         ldq_23_bits_uop_bypassable;
  reg  [4:0]  ldq_23_bits_uop_mem_cmd;
  reg  [1:0]  ldq_23_bits_uop_mem_size;
  reg         ldq_23_bits_uop_mem_signed;
  reg         ldq_23_bits_uop_is_fence;
  reg         ldq_23_bits_uop_is_fencei;
  reg         ldq_23_bits_uop_is_amo;
  reg         ldq_23_bits_uop_uses_ldq;
  reg         ldq_23_bits_uop_uses_stq;
  reg         ldq_23_bits_uop_is_sys_pc2epc;
  reg         ldq_23_bits_uop_is_unique;
  reg         ldq_23_bits_uop_flush_on_commit;
  reg         ldq_23_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_23_bits_uop_ldst;
  reg  [5:0]  ldq_23_bits_uop_lrs1;
  reg  [5:0]  ldq_23_bits_uop_lrs2;
  reg  [5:0]  ldq_23_bits_uop_lrs3;
  reg         ldq_23_bits_uop_ldst_val;
  reg  [1:0]  ldq_23_bits_uop_dst_rtype;
  reg  [1:0]  ldq_23_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_23_bits_uop_lrs2_rtype;
  reg         ldq_23_bits_uop_frs3_en;
  reg         ldq_23_bits_uop_fp_val;
  reg         ldq_23_bits_uop_fp_single;
  reg         ldq_23_bits_uop_xcpt_pf_if;
  reg         ldq_23_bits_uop_xcpt_ae_if;
  reg         ldq_23_bits_uop_xcpt_ma_if;
  reg         ldq_23_bits_uop_bp_debug_if;
  reg         ldq_23_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_23_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_23_bits_uop_debug_tsrc;
  reg         ldq_23_bits_addr_valid;
  reg  [39:0] ldq_23_bits_addr_bits;
  reg         ldq_23_bits_addr_is_virtual;
  reg         ldq_23_bits_addr_is_uncacheable;
  reg         ldq_23_bits_executed;
  reg         ldq_23_bits_succeeded;
  reg         ldq_23_bits_order_fail;
  reg         ldq_23_bits_observed;
  reg  [31:0] ldq_23_bits_st_dep_mask;
  reg  [4:0]  ldq_23_bits_youngest_stq_idx;
  reg         ldq_23_bits_forward_std_val;
  reg  [4:0]  ldq_23_bits_forward_stq_idx;
  reg         ldq_24_valid;
  reg  [6:0]  ldq_24_bits_uop_uopc;
  reg  [31:0] ldq_24_bits_uop_inst;
  reg  [31:0] ldq_24_bits_uop_debug_inst;
  reg         ldq_24_bits_uop_is_rvc;
  reg  [39:0] ldq_24_bits_uop_debug_pc;
  reg  [2:0]  ldq_24_bits_uop_iq_type;
  reg  [9:0]  ldq_24_bits_uop_fu_code;
  reg  [3:0]  ldq_24_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_24_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_24_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_24_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_24_bits_uop_ctrl_op_fcn;
  reg         ldq_24_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_24_bits_uop_ctrl_csr_cmd;
  reg         ldq_24_bits_uop_ctrl_is_load;
  reg         ldq_24_bits_uop_ctrl_is_sta;
  reg         ldq_24_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_24_bits_uop_iw_state;
  reg         ldq_24_bits_uop_iw_p1_poisoned;
  reg         ldq_24_bits_uop_iw_p2_poisoned;
  reg         ldq_24_bits_uop_is_br;
  reg         ldq_24_bits_uop_is_jalr;
  reg         ldq_24_bits_uop_is_jal;
  reg         ldq_24_bits_uop_is_sfb;
  reg  [19:0] ldq_24_bits_uop_br_mask;
  reg  [4:0]  ldq_24_bits_uop_br_tag;
  reg  [5:0]  ldq_24_bits_uop_ftq_idx;
  reg         ldq_24_bits_uop_edge_inst;
  reg  [5:0]  ldq_24_bits_uop_pc_lob;
  reg         ldq_24_bits_uop_taken;
  reg  [19:0] ldq_24_bits_uop_imm_packed;
  reg  [11:0] ldq_24_bits_uop_csr_addr;
  reg  [6:0]  ldq_24_bits_uop_rob_idx;
  reg  [4:0]  ldq_24_bits_uop_ldq_idx;
  reg  [4:0]  ldq_24_bits_uop_stq_idx;
  reg  [1:0]  ldq_24_bits_uop_rxq_idx;
  reg  [6:0]  ldq_24_bits_uop_pdst;
  reg  [6:0]  ldq_24_bits_uop_prs1;
  reg  [6:0]  ldq_24_bits_uop_prs2;
  reg  [6:0]  ldq_24_bits_uop_prs3;
  reg         ldq_24_bits_uop_prs1_busy;
  reg         ldq_24_bits_uop_prs2_busy;
  reg         ldq_24_bits_uop_prs3_busy;
  reg  [6:0]  ldq_24_bits_uop_stale_pdst;
  reg         ldq_24_bits_uop_exception;
  reg  [63:0] ldq_24_bits_uop_exc_cause;
  reg         ldq_24_bits_uop_bypassable;
  reg  [4:0]  ldq_24_bits_uop_mem_cmd;
  reg  [1:0]  ldq_24_bits_uop_mem_size;
  reg         ldq_24_bits_uop_mem_signed;
  reg         ldq_24_bits_uop_is_fence;
  reg         ldq_24_bits_uop_is_fencei;
  reg         ldq_24_bits_uop_is_amo;
  reg         ldq_24_bits_uop_uses_ldq;
  reg         ldq_24_bits_uop_uses_stq;
  reg         ldq_24_bits_uop_is_sys_pc2epc;
  reg         ldq_24_bits_uop_is_unique;
  reg         ldq_24_bits_uop_flush_on_commit;
  reg         ldq_24_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_24_bits_uop_ldst;
  reg  [5:0]  ldq_24_bits_uop_lrs1;
  reg  [5:0]  ldq_24_bits_uop_lrs2;
  reg  [5:0]  ldq_24_bits_uop_lrs3;
  reg         ldq_24_bits_uop_ldst_val;
  reg  [1:0]  ldq_24_bits_uop_dst_rtype;
  reg  [1:0]  ldq_24_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_24_bits_uop_lrs2_rtype;
  reg         ldq_24_bits_uop_frs3_en;
  reg         ldq_24_bits_uop_fp_val;
  reg         ldq_24_bits_uop_fp_single;
  reg         ldq_24_bits_uop_xcpt_pf_if;
  reg         ldq_24_bits_uop_xcpt_ae_if;
  reg         ldq_24_bits_uop_xcpt_ma_if;
  reg         ldq_24_bits_uop_bp_debug_if;
  reg         ldq_24_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_24_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_24_bits_uop_debug_tsrc;
  reg         ldq_24_bits_addr_valid;
  reg  [39:0] ldq_24_bits_addr_bits;
  reg         ldq_24_bits_addr_is_virtual;
  reg         ldq_24_bits_addr_is_uncacheable;
  reg         ldq_24_bits_executed;
  reg         ldq_24_bits_succeeded;
  reg         ldq_24_bits_order_fail;
  reg         ldq_24_bits_observed;
  reg  [31:0] ldq_24_bits_st_dep_mask;
  reg  [4:0]  ldq_24_bits_youngest_stq_idx;
  reg         ldq_24_bits_forward_std_val;
  reg  [4:0]  ldq_24_bits_forward_stq_idx;
  reg         ldq_25_valid;
  reg  [6:0]  ldq_25_bits_uop_uopc;
  reg  [31:0] ldq_25_bits_uop_inst;
  reg  [31:0] ldq_25_bits_uop_debug_inst;
  reg         ldq_25_bits_uop_is_rvc;
  reg  [39:0] ldq_25_bits_uop_debug_pc;
  reg  [2:0]  ldq_25_bits_uop_iq_type;
  reg  [9:0]  ldq_25_bits_uop_fu_code;
  reg  [3:0]  ldq_25_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_25_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_25_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_25_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_25_bits_uop_ctrl_op_fcn;
  reg         ldq_25_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_25_bits_uop_ctrl_csr_cmd;
  reg         ldq_25_bits_uop_ctrl_is_load;
  reg         ldq_25_bits_uop_ctrl_is_sta;
  reg         ldq_25_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_25_bits_uop_iw_state;
  reg         ldq_25_bits_uop_iw_p1_poisoned;
  reg         ldq_25_bits_uop_iw_p2_poisoned;
  reg         ldq_25_bits_uop_is_br;
  reg         ldq_25_bits_uop_is_jalr;
  reg         ldq_25_bits_uop_is_jal;
  reg         ldq_25_bits_uop_is_sfb;
  reg  [19:0] ldq_25_bits_uop_br_mask;
  reg  [4:0]  ldq_25_bits_uop_br_tag;
  reg  [5:0]  ldq_25_bits_uop_ftq_idx;
  reg         ldq_25_bits_uop_edge_inst;
  reg  [5:0]  ldq_25_bits_uop_pc_lob;
  reg         ldq_25_bits_uop_taken;
  reg  [19:0] ldq_25_bits_uop_imm_packed;
  reg  [11:0] ldq_25_bits_uop_csr_addr;
  reg  [6:0]  ldq_25_bits_uop_rob_idx;
  reg  [4:0]  ldq_25_bits_uop_ldq_idx;
  reg  [4:0]  ldq_25_bits_uop_stq_idx;
  reg  [1:0]  ldq_25_bits_uop_rxq_idx;
  reg  [6:0]  ldq_25_bits_uop_pdst;
  reg  [6:0]  ldq_25_bits_uop_prs1;
  reg  [6:0]  ldq_25_bits_uop_prs2;
  reg  [6:0]  ldq_25_bits_uop_prs3;
  reg         ldq_25_bits_uop_prs1_busy;
  reg         ldq_25_bits_uop_prs2_busy;
  reg         ldq_25_bits_uop_prs3_busy;
  reg  [6:0]  ldq_25_bits_uop_stale_pdst;
  reg         ldq_25_bits_uop_exception;
  reg  [63:0] ldq_25_bits_uop_exc_cause;
  reg         ldq_25_bits_uop_bypassable;
  reg  [4:0]  ldq_25_bits_uop_mem_cmd;
  reg  [1:0]  ldq_25_bits_uop_mem_size;
  reg         ldq_25_bits_uop_mem_signed;
  reg         ldq_25_bits_uop_is_fence;
  reg         ldq_25_bits_uop_is_fencei;
  reg         ldq_25_bits_uop_is_amo;
  reg         ldq_25_bits_uop_uses_ldq;
  reg         ldq_25_bits_uop_uses_stq;
  reg         ldq_25_bits_uop_is_sys_pc2epc;
  reg         ldq_25_bits_uop_is_unique;
  reg         ldq_25_bits_uop_flush_on_commit;
  reg         ldq_25_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_25_bits_uop_ldst;
  reg  [5:0]  ldq_25_bits_uop_lrs1;
  reg  [5:0]  ldq_25_bits_uop_lrs2;
  reg  [5:0]  ldq_25_bits_uop_lrs3;
  reg         ldq_25_bits_uop_ldst_val;
  reg  [1:0]  ldq_25_bits_uop_dst_rtype;
  reg  [1:0]  ldq_25_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_25_bits_uop_lrs2_rtype;
  reg         ldq_25_bits_uop_frs3_en;
  reg         ldq_25_bits_uop_fp_val;
  reg         ldq_25_bits_uop_fp_single;
  reg         ldq_25_bits_uop_xcpt_pf_if;
  reg         ldq_25_bits_uop_xcpt_ae_if;
  reg         ldq_25_bits_uop_xcpt_ma_if;
  reg         ldq_25_bits_uop_bp_debug_if;
  reg         ldq_25_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_25_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_25_bits_uop_debug_tsrc;
  reg         ldq_25_bits_addr_valid;
  reg  [39:0] ldq_25_bits_addr_bits;
  reg         ldq_25_bits_addr_is_virtual;
  reg         ldq_25_bits_addr_is_uncacheable;
  reg         ldq_25_bits_executed;
  reg         ldq_25_bits_succeeded;
  reg         ldq_25_bits_order_fail;
  reg         ldq_25_bits_observed;
  reg  [31:0] ldq_25_bits_st_dep_mask;
  reg  [4:0]  ldq_25_bits_youngest_stq_idx;
  reg         ldq_25_bits_forward_std_val;
  reg  [4:0]  ldq_25_bits_forward_stq_idx;
  reg         ldq_26_valid;
  reg  [6:0]  ldq_26_bits_uop_uopc;
  reg  [31:0] ldq_26_bits_uop_inst;
  reg  [31:0] ldq_26_bits_uop_debug_inst;
  reg         ldq_26_bits_uop_is_rvc;
  reg  [39:0] ldq_26_bits_uop_debug_pc;
  reg  [2:0]  ldq_26_bits_uop_iq_type;
  reg  [9:0]  ldq_26_bits_uop_fu_code;
  reg  [3:0]  ldq_26_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_26_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_26_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_26_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_26_bits_uop_ctrl_op_fcn;
  reg         ldq_26_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_26_bits_uop_ctrl_csr_cmd;
  reg         ldq_26_bits_uop_ctrl_is_load;
  reg         ldq_26_bits_uop_ctrl_is_sta;
  reg         ldq_26_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_26_bits_uop_iw_state;
  reg         ldq_26_bits_uop_iw_p1_poisoned;
  reg         ldq_26_bits_uop_iw_p2_poisoned;
  reg         ldq_26_bits_uop_is_br;
  reg         ldq_26_bits_uop_is_jalr;
  reg         ldq_26_bits_uop_is_jal;
  reg         ldq_26_bits_uop_is_sfb;
  reg  [19:0] ldq_26_bits_uop_br_mask;
  reg  [4:0]  ldq_26_bits_uop_br_tag;
  reg  [5:0]  ldq_26_bits_uop_ftq_idx;
  reg         ldq_26_bits_uop_edge_inst;
  reg  [5:0]  ldq_26_bits_uop_pc_lob;
  reg         ldq_26_bits_uop_taken;
  reg  [19:0] ldq_26_bits_uop_imm_packed;
  reg  [11:0] ldq_26_bits_uop_csr_addr;
  reg  [6:0]  ldq_26_bits_uop_rob_idx;
  reg  [4:0]  ldq_26_bits_uop_ldq_idx;
  reg  [4:0]  ldq_26_bits_uop_stq_idx;
  reg  [1:0]  ldq_26_bits_uop_rxq_idx;
  reg  [6:0]  ldq_26_bits_uop_pdst;
  reg  [6:0]  ldq_26_bits_uop_prs1;
  reg  [6:0]  ldq_26_bits_uop_prs2;
  reg  [6:0]  ldq_26_bits_uop_prs3;
  reg         ldq_26_bits_uop_prs1_busy;
  reg         ldq_26_bits_uop_prs2_busy;
  reg         ldq_26_bits_uop_prs3_busy;
  reg  [6:0]  ldq_26_bits_uop_stale_pdst;
  reg         ldq_26_bits_uop_exception;
  reg  [63:0] ldq_26_bits_uop_exc_cause;
  reg         ldq_26_bits_uop_bypassable;
  reg  [4:0]  ldq_26_bits_uop_mem_cmd;
  reg  [1:0]  ldq_26_bits_uop_mem_size;
  reg         ldq_26_bits_uop_mem_signed;
  reg         ldq_26_bits_uop_is_fence;
  reg         ldq_26_bits_uop_is_fencei;
  reg         ldq_26_bits_uop_is_amo;
  reg         ldq_26_bits_uop_uses_ldq;
  reg         ldq_26_bits_uop_uses_stq;
  reg         ldq_26_bits_uop_is_sys_pc2epc;
  reg         ldq_26_bits_uop_is_unique;
  reg         ldq_26_bits_uop_flush_on_commit;
  reg         ldq_26_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_26_bits_uop_ldst;
  reg  [5:0]  ldq_26_bits_uop_lrs1;
  reg  [5:0]  ldq_26_bits_uop_lrs2;
  reg  [5:0]  ldq_26_bits_uop_lrs3;
  reg         ldq_26_bits_uop_ldst_val;
  reg  [1:0]  ldq_26_bits_uop_dst_rtype;
  reg  [1:0]  ldq_26_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_26_bits_uop_lrs2_rtype;
  reg         ldq_26_bits_uop_frs3_en;
  reg         ldq_26_bits_uop_fp_val;
  reg         ldq_26_bits_uop_fp_single;
  reg         ldq_26_bits_uop_xcpt_pf_if;
  reg         ldq_26_bits_uop_xcpt_ae_if;
  reg         ldq_26_bits_uop_xcpt_ma_if;
  reg         ldq_26_bits_uop_bp_debug_if;
  reg         ldq_26_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_26_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_26_bits_uop_debug_tsrc;
  reg         ldq_26_bits_addr_valid;
  reg  [39:0] ldq_26_bits_addr_bits;
  reg         ldq_26_bits_addr_is_virtual;
  reg         ldq_26_bits_addr_is_uncacheable;
  reg         ldq_26_bits_executed;
  reg         ldq_26_bits_succeeded;
  reg         ldq_26_bits_order_fail;
  reg         ldq_26_bits_observed;
  reg  [31:0] ldq_26_bits_st_dep_mask;
  reg  [4:0]  ldq_26_bits_youngest_stq_idx;
  reg         ldq_26_bits_forward_std_val;
  reg  [4:0]  ldq_26_bits_forward_stq_idx;
  reg         ldq_27_valid;
  reg  [6:0]  ldq_27_bits_uop_uopc;
  reg  [31:0] ldq_27_bits_uop_inst;
  reg  [31:0] ldq_27_bits_uop_debug_inst;
  reg         ldq_27_bits_uop_is_rvc;
  reg  [39:0] ldq_27_bits_uop_debug_pc;
  reg  [2:0]  ldq_27_bits_uop_iq_type;
  reg  [9:0]  ldq_27_bits_uop_fu_code;
  reg  [3:0]  ldq_27_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_27_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_27_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_27_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_27_bits_uop_ctrl_op_fcn;
  reg         ldq_27_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_27_bits_uop_ctrl_csr_cmd;
  reg         ldq_27_bits_uop_ctrl_is_load;
  reg         ldq_27_bits_uop_ctrl_is_sta;
  reg         ldq_27_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_27_bits_uop_iw_state;
  reg         ldq_27_bits_uop_iw_p1_poisoned;
  reg         ldq_27_bits_uop_iw_p2_poisoned;
  reg         ldq_27_bits_uop_is_br;
  reg         ldq_27_bits_uop_is_jalr;
  reg         ldq_27_bits_uop_is_jal;
  reg         ldq_27_bits_uop_is_sfb;
  reg  [19:0] ldq_27_bits_uop_br_mask;
  reg  [4:0]  ldq_27_bits_uop_br_tag;
  reg  [5:0]  ldq_27_bits_uop_ftq_idx;
  reg         ldq_27_bits_uop_edge_inst;
  reg  [5:0]  ldq_27_bits_uop_pc_lob;
  reg         ldq_27_bits_uop_taken;
  reg  [19:0] ldq_27_bits_uop_imm_packed;
  reg  [11:0] ldq_27_bits_uop_csr_addr;
  reg  [6:0]  ldq_27_bits_uop_rob_idx;
  reg  [4:0]  ldq_27_bits_uop_ldq_idx;
  reg  [4:0]  ldq_27_bits_uop_stq_idx;
  reg  [1:0]  ldq_27_bits_uop_rxq_idx;
  reg  [6:0]  ldq_27_bits_uop_pdst;
  reg  [6:0]  ldq_27_bits_uop_prs1;
  reg  [6:0]  ldq_27_bits_uop_prs2;
  reg  [6:0]  ldq_27_bits_uop_prs3;
  reg         ldq_27_bits_uop_prs1_busy;
  reg         ldq_27_bits_uop_prs2_busy;
  reg         ldq_27_bits_uop_prs3_busy;
  reg  [6:0]  ldq_27_bits_uop_stale_pdst;
  reg         ldq_27_bits_uop_exception;
  reg  [63:0] ldq_27_bits_uop_exc_cause;
  reg         ldq_27_bits_uop_bypassable;
  reg  [4:0]  ldq_27_bits_uop_mem_cmd;
  reg  [1:0]  ldq_27_bits_uop_mem_size;
  reg         ldq_27_bits_uop_mem_signed;
  reg         ldq_27_bits_uop_is_fence;
  reg         ldq_27_bits_uop_is_fencei;
  reg         ldq_27_bits_uop_is_amo;
  reg         ldq_27_bits_uop_uses_ldq;
  reg         ldq_27_bits_uop_uses_stq;
  reg         ldq_27_bits_uop_is_sys_pc2epc;
  reg         ldq_27_bits_uop_is_unique;
  reg         ldq_27_bits_uop_flush_on_commit;
  reg         ldq_27_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_27_bits_uop_ldst;
  reg  [5:0]  ldq_27_bits_uop_lrs1;
  reg  [5:0]  ldq_27_bits_uop_lrs2;
  reg  [5:0]  ldq_27_bits_uop_lrs3;
  reg         ldq_27_bits_uop_ldst_val;
  reg  [1:0]  ldq_27_bits_uop_dst_rtype;
  reg  [1:0]  ldq_27_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_27_bits_uop_lrs2_rtype;
  reg         ldq_27_bits_uop_frs3_en;
  reg         ldq_27_bits_uop_fp_val;
  reg         ldq_27_bits_uop_fp_single;
  reg         ldq_27_bits_uop_xcpt_pf_if;
  reg         ldq_27_bits_uop_xcpt_ae_if;
  reg         ldq_27_bits_uop_xcpt_ma_if;
  reg         ldq_27_bits_uop_bp_debug_if;
  reg         ldq_27_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_27_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_27_bits_uop_debug_tsrc;
  reg         ldq_27_bits_addr_valid;
  reg  [39:0] ldq_27_bits_addr_bits;
  reg         ldq_27_bits_addr_is_virtual;
  reg         ldq_27_bits_addr_is_uncacheable;
  reg         ldq_27_bits_executed;
  reg         ldq_27_bits_succeeded;
  reg         ldq_27_bits_order_fail;
  reg         ldq_27_bits_observed;
  reg  [31:0] ldq_27_bits_st_dep_mask;
  reg  [4:0]  ldq_27_bits_youngest_stq_idx;
  reg         ldq_27_bits_forward_std_val;
  reg  [4:0]  ldq_27_bits_forward_stq_idx;
  reg         ldq_28_valid;
  reg  [6:0]  ldq_28_bits_uop_uopc;
  reg  [31:0] ldq_28_bits_uop_inst;
  reg  [31:0] ldq_28_bits_uop_debug_inst;
  reg         ldq_28_bits_uop_is_rvc;
  reg  [39:0] ldq_28_bits_uop_debug_pc;
  reg  [2:0]  ldq_28_bits_uop_iq_type;
  reg  [9:0]  ldq_28_bits_uop_fu_code;
  reg  [3:0]  ldq_28_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_28_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_28_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_28_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_28_bits_uop_ctrl_op_fcn;
  reg         ldq_28_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_28_bits_uop_ctrl_csr_cmd;
  reg         ldq_28_bits_uop_ctrl_is_load;
  reg         ldq_28_bits_uop_ctrl_is_sta;
  reg         ldq_28_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_28_bits_uop_iw_state;
  reg         ldq_28_bits_uop_iw_p1_poisoned;
  reg         ldq_28_bits_uop_iw_p2_poisoned;
  reg         ldq_28_bits_uop_is_br;
  reg         ldq_28_bits_uop_is_jalr;
  reg         ldq_28_bits_uop_is_jal;
  reg         ldq_28_bits_uop_is_sfb;
  reg  [19:0] ldq_28_bits_uop_br_mask;
  reg  [4:0]  ldq_28_bits_uop_br_tag;
  reg  [5:0]  ldq_28_bits_uop_ftq_idx;
  reg         ldq_28_bits_uop_edge_inst;
  reg  [5:0]  ldq_28_bits_uop_pc_lob;
  reg         ldq_28_bits_uop_taken;
  reg  [19:0] ldq_28_bits_uop_imm_packed;
  reg  [11:0] ldq_28_bits_uop_csr_addr;
  reg  [6:0]  ldq_28_bits_uop_rob_idx;
  reg  [4:0]  ldq_28_bits_uop_ldq_idx;
  reg  [4:0]  ldq_28_bits_uop_stq_idx;
  reg  [1:0]  ldq_28_bits_uop_rxq_idx;
  reg  [6:0]  ldq_28_bits_uop_pdst;
  reg  [6:0]  ldq_28_bits_uop_prs1;
  reg  [6:0]  ldq_28_bits_uop_prs2;
  reg  [6:0]  ldq_28_bits_uop_prs3;
  reg         ldq_28_bits_uop_prs1_busy;
  reg         ldq_28_bits_uop_prs2_busy;
  reg         ldq_28_bits_uop_prs3_busy;
  reg  [6:0]  ldq_28_bits_uop_stale_pdst;
  reg         ldq_28_bits_uop_exception;
  reg  [63:0] ldq_28_bits_uop_exc_cause;
  reg         ldq_28_bits_uop_bypassable;
  reg  [4:0]  ldq_28_bits_uop_mem_cmd;
  reg  [1:0]  ldq_28_bits_uop_mem_size;
  reg         ldq_28_bits_uop_mem_signed;
  reg         ldq_28_bits_uop_is_fence;
  reg         ldq_28_bits_uop_is_fencei;
  reg         ldq_28_bits_uop_is_amo;
  reg         ldq_28_bits_uop_uses_ldq;
  reg         ldq_28_bits_uop_uses_stq;
  reg         ldq_28_bits_uop_is_sys_pc2epc;
  reg         ldq_28_bits_uop_is_unique;
  reg         ldq_28_bits_uop_flush_on_commit;
  reg         ldq_28_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_28_bits_uop_ldst;
  reg  [5:0]  ldq_28_bits_uop_lrs1;
  reg  [5:0]  ldq_28_bits_uop_lrs2;
  reg  [5:0]  ldq_28_bits_uop_lrs3;
  reg         ldq_28_bits_uop_ldst_val;
  reg  [1:0]  ldq_28_bits_uop_dst_rtype;
  reg  [1:0]  ldq_28_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_28_bits_uop_lrs2_rtype;
  reg         ldq_28_bits_uop_frs3_en;
  reg         ldq_28_bits_uop_fp_val;
  reg         ldq_28_bits_uop_fp_single;
  reg         ldq_28_bits_uop_xcpt_pf_if;
  reg         ldq_28_bits_uop_xcpt_ae_if;
  reg         ldq_28_bits_uop_xcpt_ma_if;
  reg         ldq_28_bits_uop_bp_debug_if;
  reg         ldq_28_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_28_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_28_bits_uop_debug_tsrc;
  reg         ldq_28_bits_addr_valid;
  reg  [39:0] ldq_28_bits_addr_bits;
  reg         ldq_28_bits_addr_is_virtual;
  reg         ldq_28_bits_addr_is_uncacheable;
  reg         ldq_28_bits_executed;
  reg         ldq_28_bits_succeeded;
  reg         ldq_28_bits_order_fail;
  reg         ldq_28_bits_observed;
  reg  [31:0] ldq_28_bits_st_dep_mask;
  reg  [4:0]  ldq_28_bits_youngest_stq_idx;
  reg         ldq_28_bits_forward_std_val;
  reg  [4:0]  ldq_28_bits_forward_stq_idx;
  reg         ldq_29_valid;
  reg  [6:0]  ldq_29_bits_uop_uopc;
  reg  [31:0] ldq_29_bits_uop_inst;
  reg  [31:0] ldq_29_bits_uop_debug_inst;
  reg         ldq_29_bits_uop_is_rvc;
  reg  [39:0] ldq_29_bits_uop_debug_pc;
  reg  [2:0]  ldq_29_bits_uop_iq_type;
  reg  [9:0]  ldq_29_bits_uop_fu_code;
  reg  [3:0]  ldq_29_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_29_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_29_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_29_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_29_bits_uop_ctrl_op_fcn;
  reg         ldq_29_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_29_bits_uop_ctrl_csr_cmd;
  reg         ldq_29_bits_uop_ctrl_is_load;
  reg         ldq_29_bits_uop_ctrl_is_sta;
  reg         ldq_29_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_29_bits_uop_iw_state;
  reg         ldq_29_bits_uop_iw_p1_poisoned;
  reg         ldq_29_bits_uop_iw_p2_poisoned;
  reg         ldq_29_bits_uop_is_br;
  reg         ldq_29_bits_uop_is_jalr;
  reg         ldq_29_bits_uop_is_jal;
  reg         ldq_29_bits_uop_is_sfb;
  reg  [19:0] ldq_29_bits_uop_br_mask;
  reg  [4:0]  ldq_29_bits_uop_br_tag;
  reg  [5:0]  ldq_29_bits_uop_ftq_idx;
  reg         ldq_29_bits_uop_edge_inst;
  reg  [5:0]  ldq_29_bits_uop_pc_lob;
  reg         ldq_29_bits_uop_taken;
  reg  [19:0] ldq_29_bits_uop_imm_packed;
  reg  [11:0] ldq_29_bits_uop_csr_addr;
  reg  [6:0]  ldq_29_bits_uop_rob_idx;
  reg  [4:0]  ldq_29_bits_uop_ldq_idx;
  reg  [4:0]  ldq_29_bits_uop_stq_idx;
  reg  [1:0]  ldq_29_bits_uop_rxq_idx;
  reg  [6:0]  ldq_29_bits_uop_pdst;
  reg  [6:0]  ldq_29_bits_uop_prs1;
  reg  [6:0]  ldq_29_bits_uop_prs2;
  reg  [6:0]  ldq_29_bits_uop_prs3;
  reg         ldq_29_bits_uop_prs1_busy;
  reg         ldq_29_bits_uop_prs2_busy;
  reg         ldq_29_bits_uop_prs3_busy;
  reg  [6:0]  ldq_29_bits_uop_stale_pdst;
  reg         ldq_29_bits_uop_exception;
  reg  [63:0] ldq_29_bits_uop_exc_cause;
  reg         ldq_29_bits_uop_bypassable;
  reg  [4:0]  ldq_29_bits_uop_mem_cmd;
  reg  [1:0]  ldq_29_bits_uop_mem_size;
  reg         ldq_29_bits_uop_mem_signed;
  reg         ldq_29_bits_uop_is_fence;
  reg         ldq_29_bits_uop_is_fencei;
  reg         ldq_29_bits_uop_is_amo;
  reg         ldq_29_bits_uop_uses_ldq;
  reg         ldq_29_bits_uop_uses_stq;
  reg         ldq_29_bits_uop_is_sys_pc2epc;
  reg         ldq_29_bits_uop_is_unique;
  reg         ldq_29_bits_uop_flush_on_commit;
  reg         ldq_29_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_29_bits_uop_ldst;
  reg  [5:0]  ldq_29_bits_uop_lrs1;
  reg  [5:0]  ldq_29_bits_uop_lrs2;
  reg  [5:0]  ldq_29_bits_uop_lrs3;
  reg         ldq_29_bits_uop_ldst_val;
  reg  [1:0]  ldq_29_bits_uop_dst_rtype;
  reg  [1:0]  ldq_29_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_29_bits_uop_lrs2_rtype;
  reg         ldq_29_bits_uop_frs3_en;
  reg         ldq_29_bits_uop_fp_val;
  reg         ldq_29_bits_uop_fp_single;
  reg         ldq_29_bits_uop_xcpt_pf_if;
  reg         ldq_29_bits_uop_xcpt_ae_if;
  reg         ldq_29_bits_uop_xcpt_ma_if;
  reg         ldq_29_bits_uop_bp_debug_if;
  reg         ldq_29_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_29_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_29_bits_uop_debug_tsrc;
  reg         ldq_29_bits_addr_valid;
  reg  [39:0] ldq_29_bits_addr_bits;
  reg         ldq_29_bits_addr_is_virtual;
  reg         ldq_29_bits_addr_is_uncacheable;
  reg         ldq_29_bits_executed;
  reg         ldq_29_bits_succeeded;
  reg         ldq_29_bits_order_fail;
  reg         ldq_29_bits_observed;
  reg  [31:0] ldq_29_bits_st_dep_mask;
  reg  [4:0]  ldq_29_bits_youngest_stq_idx;
  reg         ldq_29_bits_forward_std_val;
  reg  [4:0]  ldq_29_bits_forward_stq_idx;
  reg         ldq_30_valid;
  reg  [6:0]  ldq_30_bits_uop_uopc;
  reg  [31:0] ldq_30_bits_uop_inst;
  reg  [31:0] ldq_30_bits_uop_debug_inst;
  reg         ldq_30_bits_uop_is_rvc;
  reg  [39:0] ldq_30_bits_uop_debug_pc;
  reg  [2:0]  ldq_30_bits_uop_iq_type;
  reg  [9:0]  ldq_30_bits_uop_fu_code;
  reg  [3:0]  ldq_30_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_30_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_30_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_30_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_30_bits_uop_ctrl_op_fcn;
  reg         ldq_30_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_30_bits_uop_ctrl_csr_cmd;
  reg         ldq_30_bits_uop_ctrl_is_load;
  reg         ldq_30_bits_uop_ctrl_is_sta;
  reg         ldq_30_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_30_bits_uop_iw_state;
  reg         ldq_30_bits_uop_iw_p1_poisoned;
  reg         ldq_30_bits_uop_iw_p2_poisoned;
  reg         ldq_30_bits_uop_is_br;
  reg         ldq_30_bits_uop_is_jalr;
  reg         ldq_30_bits_uop_is_jal;
  reg         ldq_30_bits_uop_is_sfb;
  reg  [19:0] ldq_30_bits_uop_br_mask;
  reg  [4:0]  ldq_30_bits_uop_br_tag;
  reg  [5:0]  ldq_30_bits_uop_ftq_idx;
  reg         ldq_30_bits_uop_edge_inst;
  reg  [5:0]  ldq_30_bits_uop_pc_lob;
  reg         ldq_30_bits_uop_taken;
  reg  [19:0] ldq_30_bits_uop_imm_packed;
  reg  [11:0] ldq_30_bits_uop_csr_addr;
  reg  [6:0]  ldq_30_bits_uop_rob_idx;
  reg  [4:0]  ldq_30_bits_uop_ldq_idx;
  reg  [4:0]  ldq_30_bits_uop_stq_idx;
  reg  [1:0]  ldq_30_bits_uop_rxq_idx;
  reg  [6:0]  ldq_30_bits_uop_pdst;
  reg  [6:0]  ldq_30_bits_uop_prs1;
  reg  [6:0]  ldq_30_bits_uop_prs2;
  reg  [6:0]  ldq_30_bits_uop_prs3;
  reg         ldq_30_bits_uop_prs1_busy;
  reg         ldq_30_bits_uop_prs2_busy;
  reg         ldq_30_bits_uop_prs3_busy;
  reg  [6:0]  ldq_30_bits_uop_stale_pdst;
  reg         ldq_30_bits_uop_exception;
  reg  [63:0] ldq_30_bits_uop_exc_cause;
  reg         ldq_30_bits_uop_bypassable;
  reg  [4:0]  ldq_30_bits_uop_mem_cmd;
  reg  [1:0]  ldq_30_bits_uop_mem_size;
  reg         ldq_30_bits_uop_mem_signed;
  reg         ldq_30_bits_uop_is_fence;
  reg         ldq_30_bits_uop_is_fencei;
  reg         ldq_30_bits_uop_is_amo;
  reg         ldq_30_bits_uop_uses_ldq;
  reg         ldq_30_bits_uop_uses_stq;
  reg         ldq_30_bits_uop_is_sys_pc2epc;
  reg         ldq_30_bits_uop_is_unique;
  reg         ldq_30_bits_uop_flush_on_commit;
  reg         ldq_30_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_30_bits_uop_ldst;
  reg  [5:0]  ldq_30_bits_uop_lrs1;
  reg  [5:0]  ldq_30_bits_uop_lrs2;
  reg  [5:0]  ldq_30_bits_uop_lrs3;
  reg         ldq_30_bits_uop_ldst_val;
  reg  [1:0]  ldq_30_bits_uop_dst_rtype;
  reg  [1:0]  ldq_30_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_30_bits_uop_lrs2_rtype;
  reg         ldq_30_bits_uop_frs3_en;
  reg         ldq_30_bits_uop_fp_val;
  reg         ldq_30_bits_uop_fp_single;
  reg         ldq_30_bits_uop_xcpt_pf_if;
  reg         ldq_30_bits_uop_xcpt_ae_if;
  reg         ldq_30_bits_uop_xcpt_ma_if;
  reg         ldq_30_bits_uop_bp_debug_if;
  reg         ldq_30_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_30_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_30_bits_uop_debug_tsrc;
  reg         ldq_30_bits_addr_valid;
  reg  [39:0] ldq_30_bits_addr_bits;
  reg         ldq_30_bits_addr_is_virtual;
  reg         ldq_30_bits_addr_is_uncacheable;
  reg         ldq_30_bits_executed;
  reg         ldq_30_bits_succeeded;
  reg         ldq_30_bits_order_fail;
  reg         ldq_30_bits_observed;
  reg  [31:0] ldq_30_bits_st_dep_mask;
  reg  [4:0]  ldq_30_bits_youngest_stq_idx;
  reg         ldq_30_bits_forward_std_val;
  reg  [4:0]  ldq_30_bits_forward_stq_idx;
  reg         ldq_31_valid;
  reg  [6:0]  ldq_31_bits_uop_uopc;
  reg  [31:0] ldq_31_bits_uop_inst;
  reg  [31:0] ldq_31_bits_uop_debug_inst;
  reg         ldq_31_bits_uop_is_rvc;
  reg  [39:0] ldq_31_bits_uop_debug_pc;
  reg  [2:0]  ldq_31_bits_uop_iq_type;
  reg  [9:0]  ldq_31_bits_uop_fu_code;
  reg  [3:0]  ldq_31_bits_uop_ctrl_br_type;
  reg  [1:0]  ldq_31_bits_uop_ctrl_op1_sel;
  reg  [2:0]  ldq_31_bits_uop_ctrl_op2_sel;
  reg  [2:0]  ldq_31_bits_uop_ctrl_imm_sel;
  reg  [3:0]  ldq_31_bits_uop_ctrl_op_fcn;
  reg         ldq_31_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  ldq_31_bits_uop_ctrl_csr_cmd;
  reg         ldq_31_bits_uop_ctrl_is_load;
  reg         ldq_31_bits_uop_ctrl_is_sta;
  reg         ldq_31_bits_uop_ctrl_is_std;
  reg  [1:0]  ldq_31_bits_uop_iw_state;
  reg         ldq_31_bits_uop_iw_p1_poisoned;
  reg         ldq_31_bits_uop_iw_p2_poisoned;
  reg         ldq_31_bits_uop_is_br;
  reg         ldq_31_bits_uop_is_jalr;
  reg         ldq_31_bits_uop_is_jal;
  reg         ldq_31_bits_uop_is_sfb;
  reg  [19:0] ldq_31_bits_uop_br_mask;
  reg  [4:0]  ldq_31_bits_uop_br_tag;
  reg  [5:0]  ldq_31_bits_uop_ftq_idx;
  reg         ldq_31_bits_uop_edge_inst;
  reg  [5:0]  ldq_31_bits_uop_pc_lob;
  reg         ldq_31_bits_uop_taken;
  reg  [19:0] ldq_31_bits_uop_imm_packed;
  reg  [11:0] ldq_31_bits_uop_csr_addr;
  reg  [6:0]  ldq_31_bits_uop_rob_idx;
  reg  [4:0]  ldq_31_bits_uop_ldq_idx;
  reg  [4:0]  ldq_31_bits_uop_stq_idx;
  reg  [1:0]  ldq_31_bits_uop_rxq_idx;
  reg  [6:0]  ldq_31_bits_uop_pdst;
  reg  [6:0]  ldq_31_bits_uop_prs1;
  reg  [6:0]  ldq_31_bits_uop_prs2;
  reg  [6:0]  ldq_31_bits_uop_prs3;
  reg         ldq_31_bits_uop_prs1_busy;
  reg         ldq_31_bits_uop_prs2_busy;
  reg         ldq_31_bits_uop_prs3_busy;
  reg  [6:0]  ldq_31_bits_uop_stale_pdst;
  reg         ldq_31_bits_uop_exception;
  reg  [63:0] ldq_31_bits_uop_exc_cause;
  reg         ldq_31_bits_uop_bypassable;
  reg  [4:0]  ldq_31_bits_uop_mem_cmd;
  reg  [1:0]  ldq_31_bits_uop_mem_size;
  reg         ldq_31_bits_uop_mem_signed;
  reg         ldq_31_bits_uop_is_fence;
  reg         ldq_31_bits_uop_is_fencei;
  reg         ldq_31_bits_uop_is_amo;
  reg         ldq_31_bits_uop_uses_ldq;
  reg         ldq_31_bits_uop_uses_stq;
  reg         ldq_31_bits_uop_is_sys_pc2epc;
  reg         ldq_31_bits_uop_is_unique;
  reg         ldq_31_bits_uop_flush_on_commit;
  reg         ldq_31_bits_uop_ldst_is_rs1;
  reg  [5:0]  ldq_31_bits_uop_ldst;
  reg  [5:0]  ldq_31_bits_uop_lrs1;
  reg  [5:0]  ldq_31_bits_uop_lrs2;
  reg  [5:0]  ldq_31_bits_uop_lrs3;
  reg         ldq_31_bits_uop_ldst_val;
  reg  [1:0]  ldq_31_bits_uop_dst_rtype;
  reg  [1:0]  ldq_31_bits_uop_lrs1_rtype;
  reg  [1:0]  ldq_31_bits_uop_lrs2_rtype;
  reg         ldq_31_bits_uop_frs3_en;
  reg         ldq_31_bits_uop_fp_val;
  reg         ldq_31_bits_uop_fp_single;
  reg         ldq_31_bits_uop_xcpt_pf_if;
  reg         ldq_31_bits_uop_xcpt_ae_if;
  reg         ldq_31_bits_uop_xcpt_ma_if;
  reg         ldq_31_bits_uop_bp_debug_if;
  reg         ldq_31_bits_uop_bp_xcpt_if;
  reg  [1:0]  ldq_31_bits_uop_debug_fsrc;
  reg  [1:0]  ldq_31_bits_uop_debug_tsrc;
  reg         ldq_31_bits_addr_valid;
  reg  [39:0] ldq_31_bits_addr_bits;
  reg         ldq_31_bits_addr_is_virtual;
  reg         ldq_31_bits_addr_is_uncacheable;
  reg         ldq_31_bits_executed;
  reg         ldq_31_bits_succeeded;
  reg         ldq_31_bits_order_fail;
  reg         ldq_31_bits_observed;
  reg  [31:0] ldq_31_bits_st_dep_mask;
  reg  [4:0]  ldq_31_bits_youngest_stq_idx;
  reg         ldq_31_bits_forward_std_val;
  reg  [4:0]  ldq_31_bits_forward_stq_idx;
  reg         stq_0_valid;
  reg  [6:0]  stq_0_bits_uop_uopc;
  reg  [31:0] stq_0_bits_uop_inst;
  reg  [31:0] stq_0_bits_uop_debug_inst;
  reg         stq_0_bits_uop_is_rvc;
  reg  [39:0] stq_0_bits_uop_debug_pc;
  reg  [2:0]  stq_0_bits_uop_iq_type;
  reg  [9:0]  stq_0_bits_uop_fu_code;
  reg  [3:0]  stq_0_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_0_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_0_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_0_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_0_bits_uop_ctrl_op_fcn;
  reg         stq_0_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_0_bits_uop_ctrl_csr_cmd;
  reg         stq_0_bits_uop_ctrl_is_load;
  reg         stq_0_bits_uop_ctrl_is_sta;
  reg         stq_0_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_0_bits_uop_iw_state;
  reg         stq_0_bits_uop_iw_p1_poisoned;
  reg         stq_0_bits_uop_iw_p2_poisoned;
  reg         stq_0_bits_uop_is_br;
  reg         stq_0_bits_uop_is_jalr;
  reg         stq_0_bits_uop_is_jal;
  reg         stq_0_bits_uop_is_sfb;
  reg  [19:0] stq_0_bits_uop_br_mask;
  reg  [4:0]  stq_0_bits_uop_br_tag;
  reg  [5:0]  stq_0_bits_uop_ftq_idx;
  reg         stq_0_bits_uop_edge_inst;
  reg  [5:0]  stq_0_bits_uop_pc_lob;
  reg         stq_0_bits_uop_taken;
  reg  [19:0] stq_0_bits_uop_imm_packed;
  reg  [11:0] stq_0_bits_uop_csr_addr;
  reg  [6:0]  stq_0_bits_uop_rob_idx;
  reg  [4:0]  stq_0_bits_uop_ldq_idx;
  reg  [4:0]  stq_0_bits_uop_stq_idx;
  reg  [1:0]  stq_0_bits_uop_rxq_idx;
  reg  [6:0]  stq_0_bits_uop_pdst;
  reg  [6:0]  stq_0_bits_uop_prs1;
  reg  [6:0]  stq_0_bits_uop_prs2;
  reg  [6:0]  stq_0_bits_uop_prs3;
  reg  [5:0]  stq_0_bits_uop_ppred;
  reg         stq_0_bits_uop_prs1_busy;
  reg         stq_0_bits_uop_prs2_busy;
  reg         stq_0_bits_uop_prs3_busy;
  reg         stq_0_bits_uop_ppred_busy;
  reg  [6:0]  stq_0_bits_uop_stale_pdst;
  reg         stq_0_bits_uop_exception;
  reg  [63:0] stq_0_bits_uop_exc_cause;
  reg         stq_0_bits_uop_bypassable;
  reg  [4:0]  stq_0_bits_uop_mem_cmd;
  reg  [1:0]  stq_0_bits_uop_mem_size;
  reg         stq_0_bits_uop_mem_signed;
  reg         stq_0_bits_uop_is_fence;
  reg         stq_0_bits_uop_is_fencei;
  reg         stq_0_bits_uop_is_amo;
  reg         stq_0_bits_uop_uses_ldq;
  reg         stq_0_bits_uop_uses_stq;
  reg         stq_0_bits_uop_is_sys_pc2epc;
  reg         stq_0_bits_uop_is_unique;
  reg         stq_0_bits_uop_flush_on_commit;
  reg         stq_0_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_0_bits_uop_ldst;
  reg  [5:0]  stq_0_bits_uop_lrs1;
  reg  [5:0]  stq_0_bits_uop_lrs2;
  reg  [5:0]  stq_0_bits_uop_lrs3;
  reg         stq_0_bits_uop_ldst_val;
  reg  [1:0]  stq_0_bits_uop_dst_rtype;
  reg  [1:0]  stq_0_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_0_bits_uop_lrs2_rtype;
  reg         stq_0_bits_uop_frs3_en;
  reg         stq_0_bits_uop_fp_val;
  reg         stq_0_bits_uop_fp_single;
  reg         stq_0_bits_uop_xcpt_pf_if;
  reg         stq_0_bits_uop_xcpt_ae_if;
  reg         stq_0_bits_uop_xcpt_ma_if;
  reg         stq_0_bits_uop_bp_debug_if;
  reg         stq_0_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_0_bits_uop_debug_fsrc;
  reg  [1:0]  stq_0_bits_uop_debug_tsrc;
  reg         stq_0_bits_addr_valid;
  reg  [39:0] stq_0_bits_addr_bits;
  reg         stq_0_bits_addr_is_virtual;
  reg         stq_0_bits_data_valid;
  reg  [63:0] stq_0_bits_data_bits;
  reg         stq_0_bits_committed;
  reg         stq_0_bits_succeeded;
  reg         stq_1_valid;
  reg  [6:0]  stq_1_bits_uop_uopc;
  reg  [31:0] stq_1_bits_uop_inst;
  reg  [31:0] stq_1_bits_uop_debug_inst;
  reg         stq_1_bits_uop_is_rvc;
  reg  [39:0] stq_1_bits_uop_debug_pc;
  reg  [2:0]  stq_1_bits_uop_iq_type;
  reg  [9:0]  stq_1_bits_uop_fu_code;
  reg  [3:0]  stq_1_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_1_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_1_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_1_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_1_bits_uop_ctrl_op_fcn;
  reg         stq_1_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_1_bits_uop_ctrl_csr_cmd;
  reg         stq_1_bits_uop_ctrl_is_load;
  reg         stq_1_bits_uop_ctrl_is_sta;
  reg         stq_1_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_1_bits_uop_iw_state;
  reg         stq_1_bits_uop_iw_p1_poisoned;
  reg         stq_1_bits_uop_iw_p2_poisoned;
  reg         stq_1_bits_uop_is_br;
  reg         stq_1_bits_uop_is_jalr;
  reg         stq_1_bits_uop_is_jal;
  reg         stq_1_bits_uop_is_sfb;
  reg  [19:0] stq_1_bits_uop_br_mask;
  reg  [4:0]  stq_1_bits_uop_br_tag;
  reg  [5:0]  stq_1_bits_uop_ftq_idx;
  reg         stq_1_bits_uop_edge_inst;
  reg  [5:0]  stq_1_bits_uop_pc_lob;
  reg         stq_1_bits_uop_taken;
  reg  [19:0] stq_1_bits_uop_imm_packed;
  reg  [11:0] stq_1_bits_uop_csr_addr;
  reg  [6:0]  stq_1_bits_uop_rob_idx;
  reg  [4:0]  stq_1_bits_uop_ldq_idx;
  reg  [4:0]  stq_1_bits_uop_stq_idx;
  reg  [1:0]  stq_1_bits_uop_rxq_idx;
  reg  [6:0]  stq_1_bits_uop_pdst;
  reg  [6:0]  stq_1_bits_uop_prs1;
  reg  [6:0]  stq_1_bits_uop_prs2;
  reg  [6:0]  stq_1_bits_uop_prs3;
  reg  [5:0]  stq_1_bits_uop_ppred;
  reg         stq_1_bits_uop_prs1_busy;
  reg         stq_1_bits_uop_prs2_busy;
  reg         stq_1_bits_uop_prs3_busy;
  reg         stq_1_bits_uop_ppred_busy;
  reg  [6:0]  stq_1_bits_uop_stale_pdst;
  reg         stq_1_bits_uop_exception;
  reg  [63:0] stq_1_bits_uop_exc_cause;
  reg         stq_1_bits_uop_bypassable;
  reg  [4:0]  stq_1_bits_uop_mem_cmd;
  reg  [1:0]  stq_1_bits_uop_mem_size;
  reg         stq_1_bits_uop_mem_signed;
  reg         stq_1_bits_uop_is_fence;
  reg         stq_1_bits_uop_is_fencei;
  reg         stq_1_bits_uop_is_amo;
  reg         stq_1_bits_uop_uses_ldq;
  reg         stq_1_bits_uop_uses_stq;
  reg         stq_1_bits_uop_is_sys_pc2epc;
  reg         stq_1_bits_uop_is_unique;
  reg         stq_1_bits_uop_flush_on_commit;
  reg         stq_1_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_1_bits_uop_ldst;
  reg  [5:0]  stq_1_bits_uop_lrs1;
  reg  [5:0]  stq_1_bits_uop_lrs2;
  reg  [5:0]  stq_1_bits_uop_lrs3;
  reg         stq_1_bits_uop_ldst_val;
  reg  [1:0]  stq_1_bits_uop_dst_rtype;
  reg  [1:0]  stq_1_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_1_bits_uop_lrs2_rtype;
  reg         stq_1_bits_uop_frs3_en;
  reg         stq_1_bits_uop_fp_val;
  reg         stq_1_bits_uop_fp_single;
  reg         stq_1_bits_uop_xcpt_pf_if;
  reg         stq_1_bits_uop_xcpt_ae_if;
  reg         stq_1_bits_uop_xcpt_ma_if;
  reg         stq_1_bits_uop_bp_debug_if;
  reg         stq_1_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_1_bits_uop_debug_fsrc;
  reg  [1:0]  stq_1_bits_uop_debug_tsrc;
  reg         stq_1_bits_addr_valid;
  reg  [39:0] stq_1_bits_addr_bits;
  reg         stq_1_bits_addr_is_virtual;
  reg         stq_1_bits_data_valid;
  reg  [63:0] stq_1_bits_data_bits;
  reg         stq_1_bits_committed;
  reg         stq_1_bits_succeeded;
  reg         stq_2_valid;
  reg  [6:0]  stq_2_bits_uop_uopc;
  reg  [31:0] stq_2_bits_uop_inst;
  reg  [31:0] stq_2_bits_uop_debug_inst;
  reg         stq_2_bits_uop_is_rvc;
  reg  [39:0] stq_2_bits_uop_debug_pc;
  reg  [2:0]  stq_2_bits_uop_iq_type;
  reg  [9:0]  stq_2_bits_uop_fu_code;
  reg  [3:0]  stq_2_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_2_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_2_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_2_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_2_bits_uop_ctrl_op_fcn;
  reg         stq_2_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_2_bits_uop_ctrl_csr_cmd;
  reg         stq_2_bits_uop_ctrl_is_load;
  reg         stq_2_bits_uop_ctrl_is_sta;
  reg         stq_2_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_2_bits_uop_iw_state;
  reg         stq_2_bits_uop_iw_p1_poisoned;
  reg         stq_2_bits_uop_iw_p2_poisoned;
  reg         stq_2_bits_uop_is_br;
  reg         stq_2_bits_uop_is_jalr;
  reg         stq_2_bits_uop_is_jal;
  reg         stq_2_bits_uop_is_sfb;
  reg  [19:0] stq_2_bits_uop_br_mask;
  reg  [4:0]  stq_2_bits_uop_br_tag;
  reg  [5:0]  stq_2_bits_uop_ftq_idx;
  reg         stq_2_bits_uop_edge_inst;
  reg  [5:0]  stq_2_bits_uop_pc_lob;
  reg         stq_2_bits_uop_taken;
  reg  [19:0] stq_2_bits_uop_imm_packed;
  reg  [11:0] stq_2_bits_uop_csr_addr;
  reg  [6:0]  stq_2_bits_uop_rob_idx;
  reg  [4:0]  stq_2_bits_uop_ldq_idx;
  reg  [4:0]  stq_2_bits_uop_stq_idx;
  reg  [1:0]  stq_2_bits_uop_rxq_idx;
  reg  [6:0]  stq_2_bits_uop_pdst;
  reg  [6:0]  stq_2_bits_uop_prs1;
  reg  [6:0]  stq_2_bits_uop_prs2;
  reg  [6:0]  stq_2_bits_uop_prs3;
  reg  [5:0]  stq_2_bits_uop_ppred;
  reg         stq_2_bits_uop_prs1_busy;
  reg         stq_2_bits_uop_prs2_busy;
  reg         stq_2_bits_uop_prs3_busy;
  reg         stq_2_bits_uop_ppred_busy;
  reg  [6:0]  stq_2_bits_uop_stale_pdst;
  reg         stq_2_bits_uop_exception;
  reg  [63:0] stq_2_bits_uop_exc_cause;
  reg         stq_2_bits_uop_bypassable;
  reg  [4:0]  stq_2_bits_uop_mem_cmd;
  reg  [1:0]  stq_2_bits_uop_mem_size;
  reg         stq_2_bits_uop_mem_signed;
  reg         stq_2_bits_uop_is_fence;
  reg         stq_2_bits_uop_is_fencei;
  reg         stq_2_bits_uop_is_amo;
  reg         stq_2_bits_uop_uses_ldq;
  reg         stq_2_bits_uop_uses_stq;
  reg         stq_2_bits_uop_is_sys_pc2epc;
  reg         stq_2_bits_uop_is_unique;
  reg         stq_2_bits_uop_flush_on_commit;
  reg         stq_2_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_2_bits_uop_ldst;
  reg  [5:0]  stq_2_bits_uop_lrs1;
  reg  [5:0]  stq_2_bits_uop_lrs2;
  reg  [5:0]  stq_2_bits_uop_lrs3;
  reg         stq_2_bits_uop_ldst_val;
  reg  [1:0]  stq_2_bits_uop_dst_rtype;
  reg  [1:0]  stq_2_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_2_bits_uop_lrs2_rtype;
  reg         stq_2_bits_uop_frs3_en;
  reg         stq_2_bits_uop_fp_val;
  reg         stq_2_bits_uop_fp_single;
  reg         stq_2_bits_uop_xcpt_pf_if;
  reg         stq_2_bits_uop_xcpt_ae_if;
  reg         stq_2_bits_uop_xcpt_ma_if;
  reg         stq_2_bits_uop_bp_debug_if;
  reg         stq_2_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_2_bits_uop_debug_fsrc;
  reg  [1:0]  stq_2_bits_uop_debug_tsrc;
  reg         stq_2_bits_addr_valid;
  reg  [39:0] stq_2_bits_addr_bits;
  reg         stq_2_bits_addr_is_virtual;
  reg         stq_2_bits_data_valid;
  reg  [63:0] stq_2_bits_data_bits;
  reg         stq_2_bits_committed;
  reg         stq_2_bits_succeeded;
  reg         stq_3_valid;
  reg  [6:0]  stq_3_bits_uop_uopc;
  reg  [31:0] stq_3_bits_uop_inst;
  reg  [31:0] stq_3_bits_uop_debug_inst;
  reg         stq_3_bits_uop_is_rvc;
  reg  [39:0] stq_3_bits_uop_debug_pc;
  reg  [2:0]  stq_3_bits_uop_iq_type;
  reg  [9:0]  stq_3_bits_uop_fu_code;
  reg  [3:0]  stq_3_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_3_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_3_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_3_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_3_bits_uop_ctrl_op_fcn;
  reg         stq_3_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_3_bits_uop_ctrl_csr_cmd;
  reg         stq_3_bits_uop_ctrl_is_load;
  reg         stq_3_bits_uop_ctrl_is_sta;
  reg         stq_3_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_3_bits_uop_iw_state;
  reg         stq_3_bits_uop_iw_p1_poisoned;
  reg         stq_3_bits_uop_iw_p2_poisoned;
  reg         stq_3_bits_uop_is_br;
  reg         stq_3_bits_uop_is_jalr;
  reg         stq_3_bits_uop_is_jal;
  reg         stq_3_bits_uop_is_sfb;
  reg  [19:0] stq_3_bits_uop_br_mask;
  reg  [4:0]  stq_3_bits_uop_br_tag;
  reg  [5:0]  stq_3_bits_uop_ftq_idx;
  reg         stq_3_bits_uop_edge_inst;
  reg  [5:0]  stq_3_bits_uop_pc_lob;
  reg         stq_3_bits_uop_taken;
  reg  [19:0] stq_3_bits_uop_imm_packed;
  reg  [11:0] stq_3_bits_uop_csr_addr;
  reg  [6:0]  stq_3_bits_uop_rob_idx;
  reg  [4:0]  stq_3_bits_uop_ldq_idx;
  reg  [4:0]  stq_3_bits_uop_stq_idx;
  reg  [1:0]  stq_3_bits_uop_rxq_idx;
  reg  [6:0]  stq_3_bits_uop_pdst;
  reg  [6:0]  stq_3_bits_uop_prs1;
  reg  [6:0]  stq_3_bits_uop_prs2;
  reg  [6:0]  stq_3_bits_uop_prs3;
  reg  [5:0]  stq_3_bits_uop_ppred;
  reg         stq_3_bits_uop_prs1_busy;
  reg         stq_3_bits_uop_prs2_busy;
  reg         stq_3_bits_uop_prs3_busy;
  reg         stq_3_bits_uop_ppred_busy;
  reg  [6:0]  stq_3_bits_uop_stale_pdst;
  reg         stq_3_bits_uop_exception;
  reg  [63:0] stq_3_bits_uop_exc_cause;
  reg         stq_3_bits_uop_bypassable;
  reg  [4:0]  stq_3_bits_uop_mem_cmd;
  reg  [1:0]  stq_3_bits_uop_mem_size;
  reg         stq_3_bits_uop_mem_signed;
  reg         stq_3_bits_uop_is_fence;
  reg         stq_3_bits_uop_is_fencei;
  reg         stq_3_bits_uop_is_amo;
  reg         stq_3_bits_uop_uses_ldq;
  reg         stq_3_bits_uop_uses_stq;
  reg         stq_3_bits_uop_is_sys_pc2epc;
  reg         stq_3_bits_uop_is_unique;
  reg         stq_3_bits_uop_flush_on_commit;
  reg         stq_3_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_3_bits_uop_ldst;
  reg  [5:0]  stq_3_bits_uop_lrs1;
  reg  [5:0]  stq_3_bits_uop_lrs2;
  reg  [5:0]  stq_3_bits_uop_lrs3;
  reg         stq_3_bits_uop_ldst_val;
  reg  [1:0]  stq_3_bits_uop_dst_rtype;
  reg  [1:0]  stq_3_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_3_bits_uop_lrs2_rtype;
  reg         stq_3_bits_uop_frs3_en;
  reg         stq_3_bits_uop_fp_val;
  reg         stq_3_bits_uop_fp_single;
  reg         stq_3_bits_uop_xcpt_pf_if;
  reg         stq_3_bits_uop_xcpt_ae_if;
  reg         stq_3_bits_uop_xcpt_ma_if;
  reg         stq_3_bits_uop_bp_debug_if;
  reg         stq_3_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_3_bits_uop_debug_fsrc;
  reg  [1:0]  stq_3_bits_uop_debug_tsrc;
  reg         stq_3_bits_addr_valid;
  reg  [39:0] stq_3_bits_addr_bits;
  reg         stq_3_bits_addr_is_virtual;
  reg         stq_3_bits_data_valid;
  reg  [63:0] stq_3_bits_data_bits;
  reg         stq_3_bits_committed;
  reg         stq_3_bits_succeeded;
  reg         stq_4_valid;
  reg  [6:0]  stq_4_bits_uop_uopc;
  reg  [31:0] stq_4_bits_uop_inst;
  reg  [31:0] stq_4_bits_uop_debug_inst;
  reg         stq_4_bits_uop_is_rvc;
  reg  [39:0] stq_4_bits_uop_debug_pc;
  reg  [2:0]  stq_4_bits_uop_iq_type;
  reg  [9:0]  stq_4_bits_uop_fu_code;
  reg  [3:0]  stq_4_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_4_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_4_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_4_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_4_bits_uop_ctrl_op_fcn;
  reg         stq_4_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_4_bits_uop_ctrl_csr_cmd;
  reg         stq_4_bits_uop_ctrl_is_load;
  reg         stq_4_bits_uop_ctrl_is_sta;
  reg         stq_4_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_4_bits_uop_iw_state;
  reg         stq_4_bits_uop_iw_p1_poisoned;
  reg         stq_4_bits_uop_iw_p2_poisoned;
  reg         stq_4_bits_uop_is_br;
  reg         stq_4_bits_uop_is_jalr;
  reg         stq_4_bits_uop_is_jal;
  reg         stq_4_bits_uop_is_sfb;
  reg  [19:0] stq_4_bits_uop_br_mask;
  reg  [4:0]  stq_4_bits_uop_br_tag;
  reg  [5:0]  stq_4_bits_uop_ftq_idx;
  reg         stq_4_bits_uop_edge_inst;
  reg  [5:0]  stq_4_bits_uop_pc_lob;
  reg         stq_4_bits_uop_taken;
  reg  [19:0] stq_4_bits_uop_imm_packed;
  reg  [11:0] stq_4_bits_uop_csr_addr;
  reg  [6:0]  stq_4_bits_uop_rob_idx;
  reg  [4:0]  stq_4_bits_uop_ldq_idx;
  reg  [4:0]  stq_4_bits_uop_stq_idx;
  reg  [1:0]  stq_4_bits_uop_rxq_idx;
  reg  [6:0]  stq_4_bits_uop_pdst;
  reg  [6:0]  stq_4_bits_uop_prs1;
  reg  [6:0]  stq_4_bits_uop_prs2;
  reg  [6:0]  stq_4_bits_uop_prs3;
  reg  [5:0]  stq_4_bits_uop_ppred;
  reg         stq_4_bits_uop_prs1_busy;
  reg         stq_4_bits_uop_prs2_busy;
  reg         stq_4_bits_uop_prs3_busy;
  reg         stq_4_bits_uop_ppred_busy;
  reg  [6:0]  stq_4_bits_uop_stale_pdst;
  reg         stq_4_bits_uop_exception;
  reg  [63:0] stq_4_bits_uop_exc_cause;
  reg         stq_4_bits_uop_bypassable;
  reg  [4:0]  stq_4_bits_uop_mem_cmd;
  reg  [1:0]  stq_4_bits_uop_mem_size;
  reg         stq_4_bits_uop_mem_signed;
  reg         stq_4_bits_uop_is_fence;
  reg         stq_4_bits_uop_is_fencei;
  reg         stq_4_bits_uop_is_amo;
  reg         stq_4_bits_uop_uses_ldq;
  reg         stq_4_bits_uop_uses_stq;
  reg         stq_4_bits_uop_is_sys_pc2epc;
  reg         stq_4_bits_uop_is_unique;
  reg         stq_4_bits_uop_flush_on_commit;
  reg         stq_4_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_4_bits_uop_ldst;
  reg  [5:0]  stq_4_bits_uop_lrs1;
  reg  [5:0]  stq_4_bits_uop_lrs2;
  reg  [5:0]  stq_4_bits_uop_lrs3;
  reg         stq_4_bits_uop_ldst_val;
  reg  [1:0]  stq_4_bits_uop_dst_rtype;
  reg  [1:0]  stq_4_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_4_bits_uop_lrs2_rtype;
  reg         stq_4_bits_uop_frs3_en;
  reg         stq_4_bits_uop_fp_val;
  reg         stq_4_bits_uop_fp_single;
  reg         stq_4_bits_uop_xcpt_pf_if;
  reg         stq_4_bits_uop_xcpt_ae_if;
  reg         stq_4_bits_uop_xcpt_ma_if;
  reg         stq_4_bits_uop_bp_debug_if;
  reg         stq_4_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_4_bits_uop_debug_fsrc;
  reg  [1:0]  stq_4_bits_uop_debug_tsrc;
  reg         stq_4_bits_addr_valid;
  reg  [39:0] stq_4_bits_addr_bits;
  reg         stq_4_bits_addr_is_virtual;
  reg         stq_4_bits_data_valid;
  reg  [63:0] stq_4_bits_data_bits;
  reg         stq_4_bits_committed;
  reg         stq_4_bits_succeeded;
  reg         stq_5_valid;
  reg  [6:0]  stq_5_bits_uop_uopc;
  reg  [31:0] stq_5_bits_uop_inst;
  reg  [31:0] stq_5_bits_uop_debug_inst;
  reg         stq_5_bits_uop_is_rvc;
  reg  [39:0] stq_5_bits_uop_debug_pc;
  reg  [2:0]  stq_5_bits_uop_iq_type;
  reg  [9:0]  stq_5_bits_uop_fu_code;
  reg  [3:0]  stq_5_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_5_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_5_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_5_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_5_bits_uop_ctrl_op_fcn;
  reg         stq_5_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_5_bits_uop_ctrl_csr_cmd;
  reg         stq_5_bits_uop_ctrl_is_load;
  reg         stq_5_bits_uop_ctrl_is_sta;
  reg         stq_5_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_5_bits_uop_iw_state;
  reg         stq_5_bits_uop_iw_p1_poisoned;
  reg         stq_5_bits_uop_iw_p2_poisoned;
  reg         stq_5_bits_uop_is_br;
  reg         stq_5_bits_uop_is_jalr;
  reg         stq_5_bits_uop_is_jal;
  reg         stq_5_bits_uop_is_sfb;
  reg  [19:0] stq_5_bits_uop_br_mask;
  reg  [4:0]  stq_5_bits_uop_br_tag;
  reg  [5:0]  stq_5_bits_uop_ftq_idx;
  reg         stq_5_bits_uop_edge_inst;
  reg  [5:0]  stq_5_bits_uop_pc_lob;
  reg         stq_5_bits_uop_taken;
  reg  [19:0] stq_5_bits_uop_imm_packed;
  reg  [11:0] stq_5_bits_uop_csr_addr;
  reg  [6:0]  stq_5_bits_uop_rob_idx;
  reg  [4:0]  stq_5_bits_uop_ldq_idx;
  reg  [4:0]  stq_5_bits_uop_stq_idx;
  reg  [1:0]  stq_5_bits_uop_rxq_idx;
  reg  [6:0]  stq_5_bits_uop_pdst;
  reg  [6:0]  stq_5_bits_uop_prs1;
  reg  [6:0]  stq_5_bits_uop_prs2;
  reg  [6:0]  stq_5_bits_uop_prs3;
  reg  [5:0]  stq_5_bits_uop_ppred;
  reg         stq_5_bits_uop_prs1_busy;
  reg         stq_5_bits_uop_prs2_busy;
  reg         stq_5_bits_uop_prs3_busy;
  reg         stq_5_bits_uop_ppred_busy;
  reg  [6:0]  stq_5_bits_uop_stale_pdst;
  reg         stq_5_bits_uop_exception;
  reg  [63:0] stq_5_bits_uop_exc_cause;
  reg         stq_5_bits_uop_bypassable;
  reg  [4:0]  stq_5_bits_uop_mem_cmd;
  reg  [1:0]  stq_5_bits_uop_mem_size;
  reg         stq_5_bits_uop_mem_signed;
  reg         stq_5_bits_uop_is_fence;
  reg         stq_5_bits_uop_is_fencei;
  reg         stq_5_bits_uop_is_amo;
  reg         stq_5_bits_uop_uses_ldq;
  reg         stq_5_bits_uop_uses_stq;
  reg         stq_5_bits_uop_is_sys_pc2epc;
  reg         stq_5_bits_uop_is_unique;
  reg         stq_5_bits_uop_flush_on_commit;
  reg         stq_5_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_5_bits_uop_ldst;
  reg  [5:0]  stq_5_bits_uop_lrs1;
  reg  [5:0]  stq_5_bits_uop_lrs2;
  reg  [5:0]  stq_5_bits_uop_lrs3;
  reg         stq_5_bits_uop_ldst_val;
  reg  [1:0]  stq_5_bits_uop_dst_rtype;
  reg  [1:0]  stq_5_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_5_bits_uop_lrs2_rtype;
  reg         stq_5_bits_uop_frs3_en;
  reg         stq_5_bits_uop_fp_val;
  reg         stq_5_bits_uop_fp_single;
  reg         stq_5_bits_uop_xcpt_pf_if;
  reg         stq_5_bits_uop_xcpt_ae_if;
  reg         stq_5_bits_uop_xcpt_ma_if;
  reg         stq_5_bits_uop_bp_debug_if;
  reg         stq_5_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_5_bits_uop_debug_fsrc;
  reg  [1:0]  stq_5_bits_uop_debug_tsrc;
  reg         stq_5_bits_addr_valid;
  reg  [39:0] stq_5_bits_addr_bits;
  reg         stq_5_bits_addr_is_virtual;
  reg         stq_5_bits_data_valid;
  reg  [63:0] stq_5_bits_data_bits;
  reg         stq_5_bits_committed;
  reg         stq_5_bits_succeeded;
  reg         stq_6_valid;
  reg  [6:0]  stq_6_bits_uop_uopc;
  reg  [31:0] stq_6_bits_uop_inst;
  reg  [31:0] stq_6_bits_uop_debug_inst;
  reg         stq_6_bits_uop_is_rvc;
  reg  [39:0] stq_6_bits_uop_debug_pc;
  reg  [2:0]  stq_6_bits_uop_iq_type;
  reg  [9:0]  stq_6_bits_uop_fu_code;
  reg  [3:0]  stq_6_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_6_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_6_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_6_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_6_bits_uop_ctrl_op_fcn;
  reg         stq_6_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_6_bits_uop_ctrl_csr_cmd;
  reg         stq_6_bits_uop_ctrl_is_load;
  reg         stq_6_bits_uop_ctrl_is_sta;
  reg         stq_6_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_6_bits_uop_iw_state;
  reg         stq_6_bits_uop_iw_p1_poisoned;
  reg         stq_6_bits_uop_iw_p2_poisoned;
  reg         stq_6_bits_uop_is_br;
  reg         stq_6_bits_uop_is_jalr;
  reg         stq_6_bits_uop_is_jal;
  reg         stq_6_bits_uop_is_sfb;
  reg  [19:0] stq_6_bits_uop_br_mask;
  reg  [4:0]  stq_6_bits_uop_br_tag;
  reg  [5:0]  stq_6_bits_uop_ftq_idx;
  reg         stq_6_bits_uop_edge_inst;
  reg  [5:0]  stq_6_bits_uop_pc_lob;
  reg         stq_6_bits_uop_taken;
  reg  [19:0] stq_6_bits_uop_imm_packed;
  reg  [11:0] stq_6_bits_uop_csr_addr;
  reg  [6:0]  stq_6_bits_uop_rob_idx;
  reg  [4:0]  stq_6_bits_uop_ldq_idx;
  reg  [4:0]  stq_6_bits_uop_stq_idx;
  reg  [1:0]  stq_6_bits_uop_rxq_idx;
  reg  [6:0]  stq_6_bits_uop_pdst;
  reg  [6:0]  stq_6_bits_uop_prs1;
  reg  [6:0]  stq_6_bits_uop_prs2;
  reg  [6:0]  stq_6_bits_uop_prs3;
  reg  [5:0]  stq_6_bits_uop_ppred;
  reg         stq_6_bits_uop_prs1_busy;
  reg         stq_6_bits_uop_prs2_busy;
  reg         stq_6_bits_uop_prs3_busy;
  reg         stq_6_bits_uop_ppred_busy;
  reg  [6:0]  stq_6_bits_uop_stale_pdst;
  reg         stq_6_bits_uop_exception;
  reg  [63:0] stq_6_bits_uop_exc_cause;
  reg         stq_6_bits_uop_bypassable;
  reg  [4:0]  stq_6_bits_uop_mem_cmd;
  reg  [1:0]  stq_6_bits_uop_mem_size;
  reg         stq_6_bits_uop_mem_signed;
  reg         stq_6_bits_uop_is_fence;
  reg         stq_6_bits_uop_is_fencei;
  reg         stq_6_bits_uop_is_amo;
  reg         stq_6_bits_uop_uses_ldq;
  reg         stq_6_bits_uop_uses_stq;
  reg         stq_6_bits_uop_is_sys_pc2epc;
  reg         stq_6_bits_uop_is_unique;
  reg         stq_6_bits_uop_flush_on_commit;
  reg         stq_6_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_6_bits_uop_ldst;
  reg  [5:0]  stq_6_bits_uop_lrs1;
  reg  [5:0]  stq_6_bits_uop_lrs2;
  reg  [5:0]  stq_6_bits_uop_lrs3;
  reg         stq_6_bits_uop_ldst_val;
  reg  [1:0]  stq_6_bits_uop_dst_rtype;
  reg  [1:0]  stq_6_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_6_bits_uop_lrs2_rtype;
  reg         stq_6_bits_uop_frs3_en;
  reg         stq_6_bits_uop_fp_val;
  reg         stq_6_bits_uop_fp_single;
  reg         stq_6_bits_uop_xcpt_pf_if;
  reg         stq_6_bits_uop_xcpt_ae_if;
  reg         stq_6_bits_uop_xcpt_ma_if;
  reg         stq_6_bits_uop_bp_debug_if;
  reg         stq_6_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_6_bits_uop_debug_fsrc;
  reg  [1:0]  stq_6_bits_uop_debug_tsrc;
  reg         stq_6_bits_addr_valid;
  reg  [39:0] stq_6_bits_addr_bits;
  reg         stq_6_bits_addr_is_virtual;
  reg         stq_6_bits_data_valid;
  reg  [63:0] stq_6_bits_data_bits;
  reg         stq_6_bits_committed;
  reg         stq_6_bits_succeeded;
  reg         stq_7_valid;
  reg  [6:0]  stq_7_bits_uop_uopc;
  reg  [31:0] stq_7_bits_uop_inst;
  reg  [31:0] stq_7_bits_uop_debug_inst;
  reg         stq_7_bits_uop_is_rvc;
  reg  [39:0] stq_7_bits_uop_debug_pc;
  reg  [2:0]  stq_7_bits_uop_iq_type;
  reg  [9:0]  stq_7_bits_uop_fu_code;
  reg  [3:0]  stq_7_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_7_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_7_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_7_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_7_bits_uop_ctrl_op_fcn;
  reg         stq_7_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_7_bits_uop_ctrl_csr_cmd;
  reg         stq_7_bits_uop_ctrl_is_load;
  reg         stq_7_bits_uop_ctrl_is_sta;
  reg         stq_7_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_7_bits_uop_iw_state;
  reg         stq_7_bits_uop_iw_p1_poisoned;
  reg         stq_7_bits_uop_iw_p2_poisoned;
  reg         stq_7_bits_uop_is_br;
  reg         stq_7_bits_uop_is_jalr;
  reg         stq_7_bits_uop_is_jal;
  reg         stq_7_bits_uop_is_sfb;
  reg  [19:0] stq_7_bits_uop_br_mask;
  reg  [4:0]  stq_7_bits_uop_br_tag;
  reg  [5:0]  stq_7_bits_uop_ftq_idx;
  reg         stq_7_bits_uop_edge_inst;
  reg  [5:0]  stq_7_bits_uop_pc_lob;
  reg         stq_7_bits_uop_taken;
  reg  [19:0] stq_7_bits_uop_imm_packed;
  reg  [11:0] stq_7_bits_uop_csr_addr;
  reg  [6:0]  stq_7_bits_uop_rob_idx;
  reg  [4:0]  stq_7_bits_uop_ldq_idx;
  reg  [4:0]  stq_7_bits_uop_stq_idx;
  reg  [1:0]  stq_7_bits_uop_rxq_idx;
  reg  [6:0]  stq_7_bits_uop_pdst;
  reg  [6:0]  stq_7_bits_uop_prs1;
  reg  [6:0]  stq_7_bits_uop_prs2;
  reg  [6:0]  stq_7_bits_uop_prs3;
  reg  [5:0]  stq_7_bits_uop_ppred;
  reg         stq_7_bits_uop_prs1_busy;
  reg         stq_7_bits_uop_prs2_busy;
  reg         stq_7_bits_uop_prs3_busy;
  reg         stq_7_bits_uop_ppred_busy;
  reg  [6:0]  stq_7_bits_uop_stale_pdst;
  reg         stq_7_bits_uop_exception;
  reg  [63:0] stq_7_bits_uop_exc_cause;
  reg         stq_7_bits_uop_bypassable;
  reg  [4:0]  stq_7_bits_uop_mem_cmd;
  reg  [1:0]  stq_7_bits_uop_mem_size;
  reg         stq_7_bits_uop_mem_signed;
  reg         stq_7_bits_uop_is_fence;
  reg         stq_7_bits_uop_is_fencei;
  reg         stq_7_bits_uop_is_amo;
  reg         stq_7_bits_uop_uses_ldq;
  reg         stq_7_bits_uop_uses_stq;
  reg         stq_7_bits_uop_is_sys_pc2epc;
  reg         stq_7_bits_uop_is_unique;
  reg         stq_7_bits_uop_flush_on_commit;
  reg         stq_7_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_7_bits_uop_ldst;
  reg  [5:0]  stq_7_bits_uop_lrs1;
  reg  [5:0]  stq_7_bits_uop_lrs2;
  reg  [5:0]  stq_7_bits_uop_lrs3;
  reg         stq_7_bits_uop_ldst_val;
  reg  [1:0]  stq_7_bits_uop_dst_rtype;
  reg  [1:0]  stq_7_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_7_bits_uop_lrs2_rtype;
  reg         stq_7_bits_uop_frs3_en;
  reg         stq_7_bits_uop_fp_val;
  reg         stq_7_bits_uop_fp_single;
  reg         stq_7_bits_uop_xcpt_pf_if;
  reg         stq_7_bits_uop_xcpt_ae_if;
  reg         stq_7_bits_uop_xcpt_ma_if;
  reg         stq_7_bits_uop_bp_debug_if;
  reg         stq_7_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_7_bits_uop_debug_fsrc;
  reg  [1:0]  stq_7_bits_uop_debug_tsrc;
  reg         stq_7_bits_addr_valid;
  reg  [39:0] stq_7_bits_addr_bits;
  reg         stq_7_bits_addr_is_virtual;
  reg         stq_7_bits_data_valid;
  reg  [63:0] stq_7_bits_data_bits;
  reg         stq_7_bits_committed;
  reg         stq_7_bits_succeeded;
  reg         stq_8_valid;
  reg  [6:0]  stq_8_bits_uop_uopc;
  reg  [31:0] stq_8_bits_uop_inst;
  reg  [31:0] stq_8_bits_uop_debug_inst;
  reg         stq_8_bits_uop_is_rvc;
  reg  [39:0] stq_8_bits_uop_debug_pc;
  reg  [2:0]  stq_8_bits_uop_iq_type;
  reg  [9:0]  stq_8_bits_uop_fu_code;
  reg  [3:0]  stq_8_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_8_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_8_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_8_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_8_bits_uop_ctrl_op_fcn;
  reg         stq_8_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_8_bits_uop_ctrl_csr_cmd;
  reg         stq_8_bits_uop_ctrl_is_load;
  reg         stq_8_bits_uop_ctrl_is_sta;
  reg         stq_8_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_8_bits_uop_iw_state;
  reg         stq_8_bits_uop_iw_p1_poisoned;
  reg         stq_8_bits_uop_iw_p2_poisoned;
  reg         stq_8_bits_uop_is_br;
  reg         stq_8_bits_uop_is_jalr;
  reg         stq_8_bits_uop_is_jal;
  reg         stq_8_bits_uop_is_sfb;
  reg  [19:0] stq_8_bits_uop_br_mask;
  reg  [4:0]  stq_8_bits_uop_br_tag;
  reg  [5:0]  stq_8_bits_uop_ftq_idx;
  reg         stq_8_bits_uop_edge_inst;
  reg  [5:0]  stq_8_bits_uop_pc_lob;
  reg         stq_8_bits_uop_taken;
  reg  [19:0] stq_8_bits_uop_imm_packed;
  reg  [11:0] stq_8_bits_uop_csr_addr;
  reg  [6:0]  stq_8_bits_uop_rob_idx;
  reg  [4:0]  stq_8_bits_uop_ldq_idx;
  reg  [4:0]  stq_8_bits_uop_stq_idx;
  reg  [1:0]  stq_8_bits_uop_rxq_idx;
  reg  [6:0]  stq_8_bits_uop_pdst;
  reg  [6:0]  stq_8_bits_uop_prs1;
  reg  [6:0]  stq_8_bits_uop_prs2;
  reg  [6:0]  stq_8_bits_uop_prs3;
  reg  [5:0]  stq_8_bits_uop_ppred;
  reg         stq_8_bits_uop_prs1_busy;
  reg         stq_8_bits_uop_prs2_busy;
  reg         stq_8_bits_uop_prs3_busy;
  reg         stq_8_bits_uop_ppred_busy;
  reg  [6:0]  stq_8_bits_uop_stale_pdst;
  reg         stq_8_bits_uop_exception;
  reg  [63:0] stq_8_bits_uop_exc_cause;
  reg         stq_8_bits_uop_bypassable;
  reg  [4:0]  stq_8_bits_uop_mem_cmd;
  reg  [1:0]  stq_8_bits_uop_mem_size;
  reg         stq_8_bits_uop_mem_signed;
  reg         stq_8_bits_uop_is_fence;
  reg         stq_8_bits_uop_is_fencei;
  reg         stq_8_bits_uop_is_amo;
  reg         stq_8_bits_uop_uses_ldq;
  reg         stq_8_bits_uop_uses_stq;
  reg         stq_8_bits_uop_is_sys_pc2epc;
  reg         stq_8_bits_uop_is_unique;
  reg         stq_8_bits_uop_flush_on_commit;
  reg         stq_8_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_8_bits_uop_ldst;
  reg  [5:0]  stq_8_bits_uop_lrs1;
  reg  [5:0]  stq_8_bits_uop_lrs2;
  reg  [5:0]  stq_8_bits_uop_lrs3;
  reg         stq_8_bits_uop_ldst_val;
  reg  [1:0]  stq_8_bits_uop_dst_rtype;
  reg  [1:0]  stq_8_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_8_bits_uop_lrs2_rtype;
  reg         stq_8_bits_uop_frs3_en;
  reg         stq_8_bits_uop_fp_val;
  reg         stq_8_bits_uop_fp_single;
  reg         stq_8_bits_uop_xcpt_pf_if;
  reg         stq_8_bits_uop_xcpt_ae_if;
  reg         stq_8_bits_uop_xcpt_ma_if;
  reg         stq_8_bits_uop_bp_debug_if;
  reg         stq_8_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_8_bits_uop_debug_fsrc;
  reg  [1:0]  stq_8_bits_uop_debug_tsrc;
  reg         stq_8_bits_addr_valid;
  reg  [39:0] stq_8_bits_addr_bits;
  reg         stq_8_bits_addr_is_virtual;
  reg         stq_8_bits_data_valid;
  reg  [63:0] stq_8_bits_data_bits;
  reg         stq_8_bits_committed;
  reg         stq_8_bits_succeeded;
  reg         stq_9_valid;
  reg  [6:0]  stq_9_bits_uop_uopc;
  reg  [31:0] stq_9_bits_uop_inst;
  reg  [31:0] stq_9_bits_uop_debug_inst;
  reg         stq_9_bits_uop_is_rvc;
  reg  [39:0] stq_9_bits_uop_debug_pc;
  reg  [2:0]  stq_9_bits_uop_iq_type;
  reg  [9:0]  stq_9_bits_uop_fu_code;
  reg  [3:0]  stq_9_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_9_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_9_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_9_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_9_bits_uop_ctrl_op_fcn;
  reg         stq_9_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_9_bits_uop_ctrl_csr_cmd;
  reg         stq_9_bits_uop_ctrl_is_load;
  reg         stq_9_bits_uop_ctrl_is_sta;
  reg         stq_9_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_9_bits_uop_iw_state;
  reg         stq_9_bits_uop_iw_p1_poisoned;
  reg         stq_9_bits_uop_iw_p2_poisoned;
  reg         stq_9_bits_uop_is_br;
  reg         stq_9_bits_uop_is_jalr;
  reg         stq_9_bits_uop_is_jal;
  reg         stq_9_bits_uop_is_sfb;
  reg  [19:0] stq_9_bits_uop_br_mask;
  reg  [4:0]  stq_9_bits_uop_br_tag;
  reg  [5:0]  stq_9_bits_uop_ftq_idx;
  reg         stq_9_bits_uop_edge_inst;
  reg  [5:0]  stq_9_bits_uop_pc_lob;
  reg         stq_9_bits_uop_taken;
  reg  [19:0] stq_9_bits_uop_imm_packed;
  reg  [11:0] stq_9_bits_uop_csr_addr;
  reg  [6:0]  stq_9_bits_uop_rob_idx;
  reg  [4:0]  stq_9_bits_uop_ldq_idx;
  reg  [4:0]  stq_9_bits_uop_stq_idx;
  reg  [1:0]  stq_9_bits_uop_rxq_idx;
  reg  [6:0]  stq_9_bits_uop_pdst;
  reg  [6:0]  stq_9_bits_uop_prs1;
  reg  [6:0]  stq_9_bits_uop_prs2;
  reg  [6:0]  stq_9_bits_uop_prs3;
  reg  [5:0]  stq_9_bits_uop_ppred;
  reg         stq_9_bits_uop_prs1_busy;
  reg         stq_9_bits_uop_prs2_busy;
  reg         stq_9_bits_uop_prs3_busy;
  reg         stq_9_bits_uop_ppred_busy;
  reg  [6:0]  stq_9_bits_uop_stale_pdst;
  reg         stq_9_bits_uop_exception;
  reg  [63:0] stq_9_bits_uop_exc_cause;
  reg         stq_9_bits_uop_bypassable;
  reg  [4:0]  stq_9_bits_uop_mem_cmd;
  reg  [1:0]  stq_9_bits_uop_mem_size;
  reg         stq_9_bits_uop_mem_signed;
  reg         stq_9_bits_uop_is_fence;
  reg         stq_9_bits_uop_is_fencei;
  reg         stq_9_bits_uop_is_amo;
  reg         stq_9_bits_uop_uses_ldq;
  reg         stq_9_bits_uop_uses_stq;
  reg         stq_9_bits_uop_is_sys_pc2epc;
  reg         stq_9_bits_uop_is_unique;
  reg         stq_9_bits_uop_flush_on_commit;
  reg         stq_9_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_9_bits_uop_ldst;
  reg  [5:0]  stq_9_bits_uop_lrs1;
  reg  [5:0]  stq_9_bits_uop_lrs2;
  reg  [5:0]  stq_9_bits_uop_lrs3;
  reg         stq_9_bits_uop_ldst_val;
  reg  [1:0]  stq_9_bits_uop_dst_rtype;
  reg  [1:0]  stq_9_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_9_bits_uop_lrs2_rtype;
  reg         stq_9_bits_uop_frs3_en;
  reg         stq_9_bits_uop_fp_val;
  reg         stq_9_bits_uop_fp_single;
  reg         stq_9_bits_uop_xcpt_pf_if;
  reg         stq_9_bits_uop_xcpt_ae_if;
  reg         stq_9_bits_uop_xcpt_ma_if;
  reg         stq_9_bits_uop_bp_debug_if;
  reg         stq_9_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_9_bits_uop_debug_fsrc;
  reg  [1:0]  stq_9_bits_uop_debug_tsrc;
  reg         stq_9_bits_addr_valid;
  reg  [39:0] stq_9_bits_addr_bits;
  reg         stq_9_bits_addr_is_virtual;
  reg         stq_9_bits_data_valid;
  reg  [63:0] stq_9_bits_data_bits;
  reg         stq_9_bits_committed;
  reg         stq_9_bits_succeeded;
  reg         stq_10_valid;
  reg  [6:0]  stq_10_bits_uop_uopc;
  reg  [31:0] stq_10_bits_uop_inst;
  reg  [31:0] stq_10_bits_uop_debug_inst;
  reg         stq_10_bits_uop_is_rvc;
  reg  [39:0] stq_10_bits_uop_debug_pc;
  reg  [2:0]  stq_10_bits_uop_iq_type;
  reg  [9:0]  stq_10_bits_uop_fu_code;
  reg  [3:0]  stq_10_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_10_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_10_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_10_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_10_bits_uop_ctrl_op_fcn;
  reg         stq_10_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_10_bits_uop_ctrl_csr_cmd;
  reg         stq_10_bits_uop_ctrl_is_load;
  reg         stq_10_bits_uop_ctrl_is_sta;
  reg         stq_10_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_10_bits_uop_iw_state;
  reg         stq_10_bits_uop_iw_p1_poisoned;
  reg         stq_10_bits_uop_iw_p2_poisoned;
  reg         stq_10_bits_uop_is_br;
  reg         stq_10_bits_uop_is_jalr;
  reg         stq_10_bits_uop_is_jal;
  reg         stq_10_bits_uop_is_sfb;
  reg  [19:0] stq_10_bits_uop_br_mask;
  reg  [4:0]  stq_10_bits_uop_br_tag;
  reg  [5:0]  stq_10_bits_uop_ftq_idx;
  reg         stq_10_bits_uop_edge_inst;
  reg  [5:0]  stq_10_bits_uop_pc_lob;
  reg         stq_10_bits_uop_taken;
  reg  [19:0] stq_10_bits_uop_imm_packed;
  reg  [11:0] stq_10_bits_uop_csr_addr;
  reg  [6:0]  stq_10_bits_uop_rob_idx;
  reg  [4:0]  stq_10_bits_uop_ldq_idx;
  reg  [4:0]  stq_10_bits_uop_stq_idx;
  reg  [1:0]  stq_10_bits_uop_rxq_idx;
  reg  [6:0]  stq_10_bits_uop_pdst;
  reg  [6:0]  stq_10_bits_uop_prs1;
  reg  [6:0]  stq_10_bits_uop_prs2;
  reg  [6:0]  stq_10_bits_uop_prs3;
  reg  [5:0]  stq_10_bits_uop_ppred;
  reg         stq_10_bits_uop_prs1_busy;
  reg         stq_10_bits_uop_prs2_busy;
  reg         stq_10_bits_uop_prs3_busy;
  reg         stq_10_bits_uop_ppred_busy;
  reg  [6:0]  stq_10_bits_uop_stale_pdst;
  reg         stq_10_bits_uop_exception;
  reg  [63:0] stq_10_bits_uop_exc_cause;
  reg         stq_10_bits_uop_bypassable;
  reg  [4:0]  stq_10_bits_uop_mem_cmd;
  reg  [1:0]  stq_10_bits_uop_mem_size;
  reg         stq_10_bits_uop_mem_signed;
  reg         stq_10_bits_uop_is_fence;
  reg         stq_10_bits_uop_is_fencei;
  reg         stq_10_bits_uop_is_amo;
  reg         stq_10_bits_uop_uses_ldq;
  reg         stq_10_bits_uop_uses_stq;
  reg         stq_10_bits_uop_is_sys_pc2epc;
  reg         stq_10_bits_uop_is_unique;
  reg         stq_10_bits_uop_flush_on_commit;
  reg         stq_10_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_10_bits_uop_ldst;
  reg  [5:0]  stq_10_bits_uop_lrs1;
  reg  [5:0]  stq_10_bits_uop_lrs2;
  reg  [5:0]  stq_10_bits_uop_lrs3;
  reg         stq_10_bits_uop_ldst_val;
  reg  [1:0]  stq_10_bits_uop_dst_rtype;
  reg  [1:0]  stq_10_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_10_bits_uop_lrs2_rtype;
  reg         stq_10_bits_uop_frs3_en;
  reg         stq_10_bits_uop_fp_val;
  reg         stq_10_bits_uop_fp_single;
  reg         stq_10_bits_uop_xcpt_pf_if;
  reg         stq_10_bits_uop_xcpt_ae_if;
  reg         stq_10_bits_uop_xcpt_ma_if;
  reg         stq_10_bits_uop_bp_debug_if;
  reg         stq_10_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_10_bits_uop_debug_fsrc;
  reg  [1:0]  stq_10_bits_uop_debug_tsrc;
  reg         stq_10_bits_addr_valid;
  reg  [39:0] stq_10_bits_addr_bits;
  reg         stq_10_bits_addr_is_virtual;
  reg         stq_10_bits_data_valid;
  reg  [63:0] stq_10_bits_data_bits;
  reg         stq_10_bits_committed;
  reg         stq_10_bits_succeeded;
  reg         stq_11_valid;
  reg  [6:0]  stq_11_bits_uop_uopc;
  reg  [31:0] stq_11_bits_uop_inst;
  reg  [31:0] stq_11_bits_uop_debug_inst;
  reg         stq_11_bits_uop_is_rvc;
  reg  [39:0] stq_11_bits_uop_debug_pc;
  reg  [2:0]  stq_11_bits_uop_iq_type;
  reg  [9:0]  stq_11_bits_uop_fu_code;
  reg  [3:0]  stq_11_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_11_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_11_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_11_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_11_bits_uop_ctrl_op_fcn;
  reg         stq_11_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_11_bits_uop_ctrl_csr_cmd;
  reg         stq_11_bits_uop_ctrl_is_load;
  reg         stq_11_bits_uop_ctrl_is_sta;
  reg         stq_11_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_11_bits_uop_iw_state;
  reg         stq_11_bits_uop_iw_p1_poisoned;
  reg         stq_11_bits_uop_iw_p2_poisoned;
  reg         stq_11_bits_uop_is_br;
  reg         stq_11_bits_uop_is_jalr;
  reg         stq_11_bits_uop_is_jal;
  reg         stq_11_bits_uop_is_sfb;
  reg  [19:0] stq_11_bits_uop_br_mask;
  reg  [4:0]  stq_11_bits_uop_br_tag;
  reg  [5:0]  stq_11_bits_uop_ftq_idx;
  reg         stq_11_bits_uop_edge_inst;
  reg  [5:0]  stq_11_bits_uop_pc_lob;
  reg         stq_11_bits_uop_taken;
  reg  [19:0] stq_11_bits_uop_imm_packed;
  reg  [11:0] stq_11_bits_uop_csr_addr;
  reg  [6:0]  stq_11_bits_uop_rob_idx;
  reg  [4:0]  stq_11_bits_uop_ldq_idx;
  reg  [4:0]  stq_11_bits_uop_stq_idx;
  reg  [1:0]  stq_11_bits_uop_rxq_idx;
  reg  [6:0]  stq_11_bits_uop_pdst;
  reg  [6:0]  stq_11_bits_uop_prs1;
  reg  [6:0]  stq_11_bits_uop_prs2;
  reg  [6:0]  stq_11_bits_uop_prs3;
  reg  [5:0]  stq_11_bits_uop_ppred;
  reg         stq_11_bits_uop_prs1_busy;
  reg         stq_11_bits_uop_prs2_busy;
  reg         stq_11_bits_uop_prs3_busy;
  reg         stq_11_bits_uop_ppred_busy;
  reg  [6:0]  stq_11_bits_uop_stale_pdst;
  reg         stq_11_bits_uop_exception;
  reg  [63:0] stq_11_bits_uop_exc_cause;
  reg         stq_11_bits_uop_bypassable;
  reg  [4:0]  stq_11_bits_uop_mem_cmd;
  reg  [1:0]  stq_11_bits_uop_mem_size;
  reg         stq_11_bits_uop_mem_signed;
  reg         stq_11_bits_uop_is_fence;
  reg         stq_11_bits_uop_is_fencei;
  reg         stq_11_bits_uop_is_amo;
  reg         stq_11_bits_uop_uses_ldq;
  reg         stq_11_bits_uop_uses_stq;
  reg         stq_11_bits_uop_is_sys_pc2epc;
  reg         stq_11_bits_uop_is_unique;
  reg         stq_11_bits_uop_flush_on_commit;
  reg         stq_11_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_11_bits_uop_ldst;
  reg  [5:0]  stq_11_bits_uop_lrs1;
  reg  [5:0]  stq_11_bits_uop_lrs2;
  reg  [5:0]  stq_11_bits_uop_lrs3;
  reg         stq_11_bits_uop_ldst_val;
  reg  [1:0]  stq_11_bits_uop_dst_rtype;
  reg  [1:0]  stq_11_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_11_bits_uop_lrs2_rtype;
  reg         stq_11_bits_uop_frs3_en;
  reg         stq_11_bits_uop_fp_val;
  reg         stq_11_bits_uop_fp_single;
  reg         stq_11_bits_uop_xcpt_pf_if;
  reg         stq_11_bits_uop_xcpt_ae_if;
  reg         stq_11_bits_uop_xcpt_ma_if;
  reg         stq_11_bits_uop_bp_debug_if;
  reg         stq_11_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_11_bits_uop_debug_fsrc;
  reg  [1:0]  stq_11_bits_uop_debug_tsrc;
  reg         stq_11_bits_addr_valid;
  reg  [39:0] stq_11_bits_addr_bits;
  reg         stq_11_bits_addr_is_virtual;
  reg         stq_11_bits_data_valid;
  reg  [63:0] stq_11_bits_data_bits;
  reg         stq_11_bits_committed;
  reg         stq_11_bits_succeeded;
  reg         stq_12_valid;
  reg  [6:0]  stq_12_bits_uop_uopc;
  reg  [31:0] stq_12_bits_uop_inst;
  reg  [31:0] stq_12_bits_uop_debug_inst;
  reg         stq_12_bits_uop_is_rvc;
  reg  [39:0] stq_12_bits_uop_debug_pc;
  reg  [2:0]  stq_12_bits_uop_iq_type;
  reg  [9:0]  stq_12_bits_uop_fu_code;
  reg  [3:0]  stq_12_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_12_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_12_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_12_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_12_bits_uop_ctrl_op_fcn;
  reg         stq_12_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_12_bits_uop_ctrl_csr_cmd;
  reg         stq_12_bits_uop_ctrl_is_load;
  reg         stq_12_bits_uop_ctrl_is_sta;
  reg         stq_12_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_12_bits_uop_iw_state;
  reg         stq_12_bits_uop_iw_p1_poisoned;
  reg         stq_12_bits_uop_iw_p2_poisoned;
  reg         stq_12_bits_uop_is_br;
  reg         stq_12_bits_uop_is_jalr;
  reg         stq_12_bits_uop_is_jal;
  reg         stq_12_bits_uop_is_sfb;
  reg  [19:0] stq_12_bits_uop_br_mask;
  reg  [4:0]  stq_12_bits_uop_br_tag;
  reg  [5:0]  stq_12_bits_uop_ftq_idx;
  reg         stq_12_bits_uop_edge_inst;
  reg  [5:0]  stq_12_bits_uop_pc_lob;
  reg         stq_12_bits_uop_taken;
  reg  [19:0] stq_12_bits_uop_imm_packed;
  reg  [11:0] stq_12_bits_uop_csr_addr;
  reg  [6:0]  stq_12_bits_uop_rob_idx;
  reg  [4:0]  stq_12_bits_uop_ldq_idx;
  reg  [4:0]  stq_12_bits_uop_stq_idx;
  reg  [1:0]  stq_12_bits_uop_rxq_idx;
  reg  [6:0]  stq_12_bits_uop_pdst;
  reg  [6:0]  stq_12_bits_uop_prs1;
  reg  [6:0]  stq_12_bits_uop_prs2;
  reg  [6:0]  stq_12_bits_uop_prs3;
  reg  [5:0]  stq_12_bits_uop_ppred;
  reg         stq_12_bits_uop_prs1_busy;
  reg         stq_12_bits_uop_prs2_busy;
  reg         stq_12_bits_uop_prs3_busy;
  reg         stq_12_bits_uop_ppred_busy;
  reg  [6:0]  stq_12_bits_uop_stale_pdst;
  reg         stq_12_bits_uop_exception;
  reg  [63:0] stq_12_bits_uop_exc_cause;
  reg         stq_12_bits_uop_bypassable;
  reg  [4:0]  stq_12_bits_uop_mem_cmd;
  reg  [1:0]  stq_12_bits_uop_mem_size;
  reg         stq_12_bits_uop_mem_signed;
  reg         stq_12_bits_uop_is_fence;
  reg         stq_12_bits_uop_is_fencei;
  reg         stq_12_bits_uop_is_amo;
  reg         stq_12_bits_uop_uses_ldq;
  reg         stq_12_bits_uop_uses_stq;
  reg         stq_12_bits_uop_is_sys_pc2epc;
  reg         stq_12_bits_uop_is_unique;
  reg         stq_12_bits_uop_flush_on_commit;
  reg         stq_12_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_12_bits_uop_ldst;
  reg  [5:0]  stq_12_bits_uop_lrs1;
  reg  [5:0]  stq_12_bits_uop_lrs2;
  reg  [5:0]  stq_12_bits_uop_lrs3;
  reg         stq_12_bits_uop_ldst_val;
  reg  [1:0]  stq_12_bits_uop_dst_rtype;
  reg  [1:0]  stq_12_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_12_bits_uop_lrs2_rtype;
  reg         stq_12_bits_uop_frs3_en;
  reg         stq_12_bits_uop_fp_val;
  reg         stq_12_bits_uop_fp_single;
  reg         stq_12_bits_uop_xcpt_pf_if;
  reg         stq_12_bits_uop_xcpt_ae_if;
  reg         stq_12_bits_uop_xcpt_ma_if;
  reg         stq_12_bits_uop_bp_debug_if;
  reg         stq_12_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_12_bits_uop_debug_fsrc;
  reg  [1:0]  stq_12_bits_uop_debug_tsrc;
  reg         stq_12_bits_addr_valid;
  reg  [39:0] stq_12_bits_addr_bits;
  reg         stq_12_bits_addr_is_virtual;
  reg         stq_12_bits_data_valid;
  reg  [63:0] stq_12_bits_data_bits;
  reg         stq_12_bits_committed;
  reg         stq_12_bits_succeeded;
  reg         stq_13_valid;
  reg  [6:0]  stq_13_bits_uop_uopc;
  reg  [31:0] stq_13_bits_uop_inst;
  reg  [31:0] stq_13_bits_uop_debug_inst;
  reg         stq_13_bits_uop_is_rvc;
  reg  [39:0] stq_13_bits_uop_debug_pc;
  reg  [2:0]  stq_13_bits_uop_iq_type;
  reg  [9:0]  stq_13_bits_uop_fu_code;
  reg  [3:0]  stq_13_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_13_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_13_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_13_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_13_bits_uop_ctrl_op_fcn;
  reg         stq_13_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_13_bits_uop_ctrl_csr_cmd;
  reg         stq_13_bits_uop_ctrl_is_load;
  reg         stq_13_bits_uop_ctrl_is_sta;
  reg         stq_13_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_13_bits_uop_iw_state;
  reg         stq_13_bits_uop_iw_p1_poisoned;
  reg         stq_13_bits_uop_iw_p2_poisoned;
  reg         stq_13_bits_uop_is_br;
  reg         stq_13_bits_uop_is_jalr;
  reg         stq_13_bits_uop_is_jal;
  reg         stq_13_bits_uop_is_sfb;
  reg  [19:0] stq_13_bits_uop_br_mask;
  reg  [4:0]  stq_13_bits_uop_br_tag;
  reg  [5:0]  stq_13_bits_uop_ftq_idx;
  reg         stq_13_bits_uop_edge_inst;
  reg  [5:0]  stq_13_bits_uop_pc_lob;
  reg         stq_13_bits_uop_taken;
  reg  [19:0] stq_13_bits_uop_imm_packed;
  reg  [11:0] stq_13_bits_uop_csr_addr;
  reg  [6:0]  stq_13_bits_uop_rob_idx;
  reg  [4:0]  stq_13_bits_uop_ldq_idx;
  reg  [4:0]  stq_13_bits_uop_stq_idx;
  reg  [1:0]  stq_13_bits_uop_rxq_idx;
  reg  [6:0]  stq_13_bits_uop_pdst;
  reg  [6:0]  stq_13_bits_uop_prs1;
  reg  [6:0]  stq_13_bits_uop_prs2;
  reg  [6:0]  stq_13_bits_uop_prs3;
  reg  [5:0]  stq_13_bits_uop_ppred;
  reg         stq_13_bits_uop_prs1_busy;
  reg         stq_13_bits_uop_prs2_busy;
  reg         stq_13_bits_uop_prs3_busy;
  reg         stq_13_bits_uop_ppred_busy;
  reg  [6:0]  stq_13_bits_uop_stale_pdst;
  reg         stq_13_bits_uop_exception;
  reg  [63:0] stq_13_bits_uop_exc_cause;
  reg         stq_13_bits_uop_bypassable;
  reg  [4:0]  stq_13_bits_uop_mem_cmd;
  reg  [1:0]  stq_13_bits_uop_mem_size;
  reg         stq_13_bits_uop_mem_signed;
  reg         stq_13_bits_uop_is_fence;
  reg         stq_13_bits_uop_is_fencei;
  reg         stq_13_bits_uop_is_amo;
  reg         stq_13_bits_uop_uses_ldq;
  reg         stq_13_bits_uop_uses_stq;
  reg         stq_13_bits_uop_is_sys_pc2epc;
  reg         stq_13_bits_uop_is_unique;
  reg         stq_13_bits_uop_flush_on_commit;
  reg         stq_13_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_13_bits_uop_ldst;
  reg  [5:0]  stq_13_bits_uop_lrs1;
  reg  [5:0]  stq_13_bits_uop_lrs2;
  reg  [5:0]  stq_13_bits_uop_lrs3;
  reg         stq_13_bits_uop_ldst_val;
  reg  [1:0]  stq_13_bits_uop_dst_rtype;
  reg  [1:0]  stq_13_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_13_bits_uop_lrs2_rtype;
  reg         stq_13_bits_uop_frs3_en;
  reg         stq_13_bits_uop_fp_val;
  reg         stq_13_bits_uop_fp_single;
  reg         stq_13_bits_uop_xcpt_pf_if;
  reg         stq_13_bits_uop_xcpt_ae_if;
  reg         stq_13_bits_uop_xcpt_ma_if;
  reg         stq_13_bits_uop_bp_debug_if;
  reg         stq_13_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_13_bits_uop_debug_fsrc;
  reg  [1:0]  stq_13_bits_uop_debug_tsrc;
  reg         stq_13_bits_addr_valid;
  reg  [39:0] stq_13_bits_addr_bits;
  reg         stq_13_bits_addr_is_virtual;
  reg         stq_13_bits_data_valid;
  reg  [63:0] stq_13_bits_data_bits;
  reg         stq_13_bits_committed;
  reg         stq_13_bits_succeeded;
  reg         stq_14_valid;
  reg  [6:0]  stq_14_bits_uop_uopc;
  reg  [31:0] stq_14_bits_uop_inst;
  reg  [31:0] stq_14_bits_uop_debug_inst;
  reg         stq_14_bits_uop_is_rvc;
  reg  [39:0] stq_14_bits_uop_debug_pc;
  reg  [2:0]  stq_14_bits_uop_iq_type;
  reg  [9:0]  stq_14_bits_uop_fu_code;
  reg  [3:0]  stq_14_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_14_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_14_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_14_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_14_bits_uop_ctrl_op_fcn;
  reg         stq_14_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_14_bits_uop_ctrl_csr_cmd;
  reg         stq_14_bits_uop_ctrl_is_load;
  reg         stq_14_bits_uop_ctrl_is_sta;
  reg         stq_14_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_14_bits_uop_iw_state;
  reg         stq_14_bits_uop_iw_p1_poisoned;
  reg         stq_14_bits_uop_iw_p2_poisoned;
  reg         stq_14_bits_uop_is_br;
  reg         stq_14_bits_uop_is_jalr;
  reg         stq_14_bits_uop_is_jal;
  reg         stq_14_bits_uop_is_sfb;
  reg  [19:0] stq_14_bits_uop_br_mask;
  reg  [4:0]  stq_14_bits_uop_br_tag;
  reg  [5:0]  stq_14_bits_uop_ftq_idx;
  reg         stq_14_bits_uop_edge_inst;
  reg  [5:0]  stq_14_bits_uop_pc_lob;
  reg         stq_14_bits_uop_taken;
  reg  [19:0] stq_14_bits_uop_imm_packed;
  reg  [11:0] stq_14_bits_uop_csr_addr;
  reg  [6:0]  stq_14_bits_uop_rob_idx;
  reg  [4:0]  stq_14_bits_uop_ldq_idx;
  reg  [4:0]  stq_14_bits_uop_stq_idx;
  reg  [1:0]  stq_14_bits_uop_rxq_idx;
  reg  [6:0]  stq_14_bits_uop_pdst;
  reg  [6:0]  stq_14_bits_uop_prs1;
  reg  [6:0]  stq_14_bits_uop_prs2;
  reg  [6:0]  stq_14_bits_uop_prs3;
  reg  [5:0]  stq_14_bits_uop_ppred;
  reg         stq_14_bits_uop_prs1_busy;
  reg         stq_14_bits_uop_prs2_busy;
  reg         stq_14_bits_uop_prs3_busy;
  reg         stq_14_bits_uop_ppred_busy;
  reg  [6:0]  stq_14_bits_uop_stale_pdst;
  reg         stq_14_bits_uop_exception;
  reg  [63:0] stq_14_bits_uop_exc_cause;
  reg         stq_14_bits_uop_bypassable;
  reg  [4:0]  stq_14_bits_uop_mem_cmd;
  reg  [1:0]  stq_14_bits_uop_mem_size;
  reg         stq_14_bits_uop_mem_signed;
  reg         stq_14_bits_uop_is_fence;
  reg         stq_14_bits_uop_is_fencei;
  reg         stq_14_bits_uop_is_amo;
  reg         stq_14_bits_uop_uses_ldq;
  reg         stq_14_bits_uop_uses_stq;
  reg         stq_14_bits_uop_is_sys_pc2epc;
  reg         stq_14_bits_uop_is_unique;
  reg         stq_14_bits_uop_flush_on_commit;
  reg         stq_14_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_14_bits_uop_ldst;
  reg  [5:0]  stq_14_bits_uop_lrs1;
  reg  [5:0]  stq_14_bits_uop_lrs2;
  reg  [5:0]  stq_14_bits_uop_lrs3;
  reg         stq_14_bits_uop_ldst_val;
  reg  [1:0]  stq_14_bits_uop_dst_rtype;
  reg  [1:0]  stq_14_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_14_bits_uop_lrs2_rtype;
  reg         stq_14_bits_uop_frs3_en;
  reg         stq_14_bits_uop_fp_val;
  reg         stq_14_bits_uop_fp_single;
  reg         stq_14_bits_uop_xcpt_pf_if;
  reg         stq_14_bits_uop_xcpt_ae_if;
  reg         stq_14_bits_uop_xcpt_ma_if;
  reg         stq_14_bits_uop_bp_debug_if;
  reg         stq_14_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_14_bits_uop_debug_fsrc;
  reg  [1:0]  stq_14_bits_uop_debug_tsrc;
  reg         stq_14_bits_addr_valid;
  reg  [39:0] stq_14_bits_addr_bits;
  reg         stq_14_bits_addr_is_virtual;
  reg         stq_14_bits_data_valid;
  reg  [63:0] stq_14_bits_data_bits;
  reg         stq_14_bits_committed;
  reg         stq_14_bits_succeeded;
  reg         stq_15_valid;
  reg  [6:0]  stq_15_bits_uop_uopc;
  reg  [31:0] stq_15_bits_uop_inst;
  reg  [31:0] stq_15_bits_uop_debug_inst;
  reg         stq_15_bits_uop_is_rvc;
  reg  [39:0] stq_15_bits_uop_debug_pc;
  reg  [2:0]  stq_15_bits_uop_iq_type;
  reg  [9:0]  stq_15_bits_uop_fu_code;
  reg  [3:0]  stq_15_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_15_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_15_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_15_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_15_bits_uop_ctrl_op_fcn;
  reg         stq_15_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_15_bits_uop_ctrl_csr_cmd;
  reg         stq_15_bits_uop_ctrl_is_load;
  reg         stq_15_bits_uop_ctrl_is_sta;
  reg         stq_15_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_15_bits_uop_iw_state;
  reg         stq_15_bits_uop_iw_p1_poisoned;
  reg         stq_15_bits_uop_iw_p2_poisoned;
  reg         stq_15_bits_uop_is_br;
  reg         stq_15_bits_uop_is_jalr;
  reg         stq_15_bits_uop_is_jal;
  reg         stq_15_bits_uop_is_sfb;
  reg  [19:0] stq_15_bits_uop_br_mask;
  reg  [4:0]  stq_15_bits_uop_br_tag;
  reg  [5:0]  stq_15_bits_uop_ftq_idx;
  reg         stq_15_bits_uop_edge_inst;
  reg  [5:0]  stq_15_bits_uop_pc_lob;
  reg         stq_15_bits_uop_taken;
  reg  [19:0] stq_15_bits_uop_imm_packed;
  reg  [11:0] stq_15_bits_uop_csr_addr;
  reg  [6:0]  stq_15_bits_uop_rob_idx;
  reg  [4:0]  stq_15_bits_uop_ldq_idx;
  reg  [4:0]  stq_15_bits_uop_stq_idx;
  reg  [1:0]  stq_15_bits_uop_rxq_idx;
  reg  [6:0]  stq_15_bits_uop_pdst;
  reg  [6:0]  stq_15_bits_uop_prs1;
  reg  [6:0]  stq_15_bits_uop_prs2;
  reg  [6:0]  stq_15_bits_uop_prs3;
  reg  [5:0]  stq_15_bits_uop_ppred;
  reg         stq_15_bits_uop_prs1_busy;
  reg         stq_15_bits_uop_prs2_busy;
  reg         stq_15_bits_uop_prs3_busy;
  reg         stq_15_bits_uop_ppred_busy;
  reg  [6:0]  stq_15_bits_uop_stale_pdst;
  reg         stq_15_bits_uop_exception;
  reg  [63:0] stq_15_bits_uop_exc_cause;
  reg         stq_15_bits_uop_bypassable;
  reg  [4:0]  stq_15_bits_uop_mem_cmd;
  reg  [1:0]  stq_15_bits_uop_mem_size;
  reg         stq_15_bits_uop_mem_signed;
  reg         stq_15_bits_uop_is_fence;
  reg         stq_15_bits_uop_is_fencei;
  reg         stq_15_bits_uop_is_amo;
  reg         stq_15_bits_uop_uses_ldq;
  reg         stq_15_bits_uop_uses_stq;
  reg         stq_15_bits_uop_is_sys_pc2epc;
  reg         stq_15_bits_uop_is_unique;
  reg         stq_15_bits_uop_flush_on_commit;
  reg         stq_15_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_15_bits_uop_ldst;
  reg  [5:0]  stq_15_bits_uop_lrs1;
  reg  [5:0]  stq_15_bits_uop_lrs2;
  reg  [5:0]  stq_15_bits_uop_lrs3;
  reg         stq_15_bits_uop_ldst_val;
  reg  [1:0]  stq_15_bits_uop_dst_rtype;
  reg  [1:0]  stq_15_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_15_bits_uop_lrs2_rtype;
  reg         stq_15_bits_uop_frs3_en;
  reg         stq_15_bits_uop_fp_val;
  reg         stq_15_bits_uop_fp_single;
  reg         stq_15_bits_uop_xcpt_pf_if;
  reg         stq_15_bits_uop_xcpt_ae_if;
  reg         stq_15_bits_uop_xcpt_ma_if;
  reg         stq_15_bits_uop_bp_debug_if;
  reg         stq_15_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_15_bits_uop_debug_fsrc;
  reg  [1:0]  stq_15_bits_uop_debug_tsrc;
  reg         stq_15_bits_addr_valid;
  reg  [39:0] stq_15_bits_addr_bits;
  reg         stq_15_bits_addr_is_virtual;
  reg         stq_15_bits_data_valid;
  reg  [63:0] stq_15_bits_data_bits;
  reg         stq_15_bits_committed;
  reg         stq_15_bits_succeeded;
  reg         stq_16_valid;
  reg  [6:0]  stq_16_bits_uop_uopc;
  reg  [31:0] stq_16_bits_uop_inst;
  reg  [31:0] stq_16_bits_uop_debug_inst;
  reg         stq_16_bits_uop_is_rvc;
  reg  [39:0] stq_16_bits_uop_debug_pc;
  reg  [2:0]  stq_16_bits_uop_iq_type;
  reg  [9:0]  stq_16_bits_uop_fu_code;
  reg  [3:0]  stq_16_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_16_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_16_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_16_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_16_bits_uop_ctrl_op_fcn;
  reg         stq_16_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_16_bits_uop_ctrl_csr_cmd;
  reg         stq_16_bits_uop_ctrl_is_load;
  reg         stq_16_bits_uop_ctrl_is_sta;
  reg         stq_16_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_16_bits_uop_iw_state;
  reg         stq_16_bits_uop_iw_p1_poisoned;
  reg         stq_16_bits_uop_iw_p2_poisoned;
  reg         stq_16_bits_uop_is_br;
  reg         stq_16_bits_uop_is_jalr;
  reg         stq_16_bits_uop_is_jal;
  reg         stq_16_bits_uop_is_sfb;
  reg  [19:0] stq_16_bits_uop_br_mask;
  reg  [4:0]  stq_16_bits_uop_br_tag;
  reg  [5:0]  stq_16_bits_uop_ftq_idx;
  reg         stq_16_bits_uop_edge_inst;
  reg  [5:0]  stq_16_bits_uop_pc_lob;
  reg         stq_16_bits_uop_taken;
  reg  [19:0] stq_16_bits_uop_imm_packed;
  reg  [11:0] stq_16_bits_uop_csr_addr;
  reg  [6:0]  stq_16_bits_uop_rob_idx;
  reg  [4:0]  stq_16_bits_uop_ldq_idx;
  reg  [4:0]  stq_16_bits_uop_stq_idx;
  reg  [1:0]  stq_16_bits_uop_rxq_idx;
  reg  [6:0]  stq_16_bits_uop_pdst;
  reg  [6:0]  stq_16_bits_uop_prs1;
  reg  [6:0]  stq_16_bits_uop_prs2;
  reg  [6:0]  stq_16_bits_uop_prs3;
  reg  [5:0]  stq_16_bits_uop_ppred;
  reg         stq_16_bits_uop_prs1_busy;
  reg         stq_16_bits_uop_prs2_busy;
  reg         stq_16_bits_uop_prs3_busy;
  reg         stq_16_bits_uop_ppred_busy;
  reg  [6:0]  stq_16_bits_uop_stale_pdst;
  reg         stq_16_bits_uop_exception;
  reg  [63:0] stq_16_bits_uop_exc_cause;
  reg         stq_16_bits_uop_bypassable;
  reg  [4:0]  stq_16_bits_uop_mem_cmd;
  reg  [1:0]  stq_16_bits_uop_mem_size;
  reg         stq_16_bits_uop_mem_signed;
  reg         stq_16_bits_uop_is_fence;
  reg         stq_16_bits_uop_is_fencei;
  reg         stq_16_bits_uop_is_amo;
  reg         stq_16_bits_uop_uses_ldq;
  reg         stq_16_bits_uop_uses_stq;
  reg         stq_16_bits_uop_is_sys_pc2epc;
  reg         stq_16_bits_uop_is_unique;
  reg         stq_16_bits_uop_flush_on_commit;
  reg         stq_16_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_16_bits_uop_ldst;
  reg  [5:0]  stq_16_bits_uop_lrs1;
  reg  [5:0]  stq_16_bits_uop_lrs2;
  reg  [5:0]  stq_16_bits_uop_lrs3;
  reg         stq_16_bits_uop_ldst_val;
  reg  [1:0]  stq_16_bits_uop_dst_rtype;
  reg  [1:0]  stq_16_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_16_bits_uop_lrs2_rtype;
  reg         stq_16_bits_uop_frs3_en;
  reg         stq_16_bits_uop_fp_val;
  reg         stq_16_bits_uop_fp_single;
  reg         stq_16_bits_uop_xcpt_pf_if;
  reg         stq_16_bits_uop_xcpt_ae_if;
  reg         stq_16_bits_uop_xcpt_ma_if;
  reg         stq_16_bits_uop_bp_debug_if;
  reg         stq_16_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_16_bits_uop_debug_fsrc;
  reg  [1:0]  stq_16_bits_uop_debug_tsrc;
  reg         stq_16_bits_addr_valid;
  reg  [39:0] stq_16_bits_addr_bits;
  reg         stq_16_bits_addr_is_virtual;
  reg         stq_16_bits_data_valid;
  reg  [63:0] stq_16_bits_data_bits;
  reg         stq_16_bits_committed;
  reg         stq_16_bits_succeeded;
  reg         stq_17_valid;
  reg  [6:0]  stq_17_bits_uop_uopc;
  reg  [31:0] stq_17_bits_uop_inst;
  reg  [31:0] stq_17_bits_uop_debug_inst;
  reg         stq_17_bits_uop_is_rvc;
  reg  [39:0] stq_17_bits_uop_debug_pc;
  reg  [2:0]  stq_17_bits_uop_iq_type;
  reg  [9:0]  stq_17_bits_uop_fu_code;
  reg  [3:0]  stq_17_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_17_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_17_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_17_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_17_bits_uop_ctrl_op_fcn;
  reg         stq_17_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_17_bits_uop_ctrl_csr_cmd;
  reg         stq_17_bits_uop_ctrl_is_load;
  reg         stq_17_bits_uop_ctrl_is_sta;
  reg         stq_17_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_17_bits_uop_iw_state;
  reg         stq_17_bits_uop_iw_p1_poisoned;
  reg         stq_17_bits_uop_iw_p2_poisoned;
  reg         stq_17_bits_uop_is_br;
  reg         stq_17_bits_uop_is_jalr;
  reg         stq_17_bits_uop_is_jal;
  reg         stq_17_bits_uop_is_sfb;
  reg  [19:0] stq_17_bits_uop_br_mask;
  reg  [4:0]  stq_17_bits_uop_br_tag;
  reg  [5:0]  stq_17_bits_uop_ftq_idx;
  reg         stq_17_bits_uop_edge_inst;
  reg  [5:0]  stq_17_bits_uop_pc_lob;
  reg         stq_17_bits_uop_taken;
  reg  [19:0] stq_17_bits_uop_imm_packed;
  reg  [11:0] stq_17_bits_uop_csr_addr;
  reg  [6:0]  stq_17_bits_uop_rob_idx;
  reg  [4:0]  stq_17_bits_uop_ldq_idx;
  reg  [4:0]  stq_17_bits_uop_stq_idx;
  reg  [1:0]  stq_17_bits_uop_rxq_idx;
  reg  [6:0]  stq_17_bits_uop_pdst;
  reg  [6:0]  stq_17_bits_uop_prs1;
  reg  [6:0]  stq_17_bits_uop_prs2;
  reg  [6:0]  stq_17_bits_uop_prs3;
  reg  [5:0]  stq_17_bits_uop_ppred;
  reg         stq_17_bits_uop_prs1_busy;
  reg         stq_17_bits_uop_prs2_busy;
  reg         stq_17_bits_uop_prs3_busy;
  reg         stq_17_bits_uop_ppred_busy;
  reg  [6:0]  stq_17_bits_uop_stale_pdst;
  reg         stq_17_bits_uop_exception;
  reg  [63:0] stq_17_bits_uop_exc_cause;
  reg         stq_17_bits_uop_bypassable;
  reg  [4:0]  stq_17_bits_uop_mem_cmd;
  reg  [1:0]  stq_17_bits_uop_mem_size;
  reg         stq_17_bits_uop_mem_signed;
  reg         stq_17_bits_uop_is_fence;
  reg         stq_17_bits_uop_is_fencei;
  reg         stq_17_bits_uop_is_amo;
  reg         stq_17_bits_uop_uses_ldq;
  reg         stq_17_bits_uop_uses_stq;
  reg         stq_17_bits_uop_is_sys_pc2epc;
  reg         stq_17_bits_uop_is_unique;
  reg         stq_17_bits_uop_flush_on_commit;
  reg         stq_17_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_17_bits_uop_ldst;
  reg  [5:0]  stq_17_bits_uop_lrs1;
  reg  [5:0]  stq_17_bits_uop_lrs2;
  reg  [5:0]  stq_17_bits_uop_lrs3;
  reg         stq_17_bits_uop_ldst_val;
  reg  [1:0]  stq_17_bits_uop_dst_rtype;
  reg  [1:0]  stq_17_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_17_bits_uop_lrs2_rtype;
  reg         stq_17_bits_uop_frs3_en;
  reg         stq_17_bits_uop_fp_val;
  reg         stq_17_bits_uop_fp_single;
  reg         stq_17_bits_uop_xcpt_pf_if;
  reg         stq_17_bits_uop_xcpt_ae_if;
  reg         stq_17_bits_uop_xcpt_ma_if;
  reg         stq_17_bits_uop_bp_debug_if;
  reg         stq_17_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_17_bits_uop_debug_fsrc;
  reg  [1:0]  stq_17_bits_uop_debug_tsrc;
  reg         stq_17_bits_addr_valid;
  reg  [39:0] stq_17_bits_addr_bits;
  reg         stq_17_bits_addr_is_virtual;
  reg         stq_17_bits_data_valid;
  reg  [63:0] stq_17_bits_data_bits;
  reg         stq_17_bits_committed;
  reg         stq_17_bits_succeeded;
  reg         stq_18_valid;
  reg  [6:0]  stq_18_bits_uop_uopc;
  reg  [31:0] stq_18_bits_uop_inst;
  reg  [31:0] stq_18_bits_uop_debug_inst;
  reg         stq_18_bits_uop_is_rvc;
  reg  [39:0] stq_18_bits_uop_debug_pc;
  reg  [2:0]  stq_18_bits_uop_iq_type;
  reg  [9:0]  stq_18_bits_uop_fu_code;
  reg  [3:0]  stq_18_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_18_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_18_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_18_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_18_bits_uop_ctrl_op_fcn;
  reg         stq_18_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_18_bits_uop_ctrl_csr_cmd;
  reg         stq_18_bits_uop_ctrl_is_load;
  reg         stq_18_bits_uop_ctrl_is_sta;
  reg         stq_18_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_18_bits_uop_iw_state;
  reg         stq_18_bits_uop_iw_p1_poisoned;
  reg         stq_18_bits_uop_iw_p2_poisoned;
  reg         stq_18_bits_uop_is_br;
  reg         stq_18_bits_uop_is_jalr;
  reg         stq_18_bits_uop_is_jal;
  reg         stq_18_bits_uop_is_sfb;
  reg  [19:0] stq_18_bits_uop_br_mask;
  reg  [4:0]  stq_18_bits_uop_br_tag;
  reg  [5:0]  stq_18_bits_uop_ftq_idx;
  reg         stq_18_bits_uop_edge_inst;
  reg  [5:0]  stq_18_bits_uop_pc_lob;
  reg         stq_18_bits_uop_taken;
  reg  [19:0] stq_18_bits_uop_imm_packed;
  reg  [11:0] stq_18_bits_uop_csr_addr;
  reg  [6:0]  stq_18_bits_uop_rob_idx;
  reg  [4:0]  stq_18_bits_uop_ldq_idx;
  reg  [4:0]  stq_18_bits_uop_stq_idx;
  reg  [1:0]  stq_18_bits_uop_rxq_idx;
  reg  [6:0]  stq_18_bits_uop_pdst;
  reg  [6:0]  stq_18_bits_uop_prs1;
  reg  [6:0]  stq_18_bits_uop_prs2;
  reg  [6:0]  stq_18_bits_uop_prs3;
  reg  [5:0]  stq_18_bits_uop_ppred;
  reg         stq_18_bits_uop_prs1_busy;
  reg         stq_18_bits_uop_prs2_busy;
  reg         stq_18_bits_uop_prs3_busy;
  reg         stq_18_bits_uop_ppred_busy;
  reg  [6:0]  stq_18_bits_uop_stale_pdst;
  reg         stq_18_bits_uop_exception;
  reg  [63:0] stq_18_bits_uop_exc_cause;
  reg         stq_18_bits_uop_bypassable;
  reg  [4:0]  stq_18_bits_uop_mem_cmd;
  reg  [1:0]  stq_18_bits_uop_mem_size;
  reg         stq_18_bits_uop_mem_signed;
  reg         stq_18_bits_uop_is_fence;
  reg         stq_18_bits_uop_is_fencei;
  reg         stq_18_bits_uop_is_amo;
  reg         stq_18_bits_uop_uses_ldq;
  reg         stq_18_bits_uop_uses_stq;
  reg         stq_18_bits_uop_is_sys_pc2epc;
  reg         stq_18_bits_uop_is_unique;
  reg         stq_18_bits_uop_flush_on_commit;
  reg         stq_18_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_18_bits_uop_ldst;
  reg  [5:0]  stq_18_bits_uop_lrs1;
  reg  [5:0]  stq_18_bits_uop_lrs2;
  reg  [5:0]  stq_18_bits_uop_lrs3;
  reg         stq_18_bits_uop_ldst_val;
  reg  [1:0]  stq_18_bits_uop_dst_rtype;
  reg  [1:0]  stq_18_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_18_bits_uop_lrs2_rtype;
  reg         stq_18_bits_uop_frs3_en;
  reg         stq_18_bits_uop_fp_val;
  reg         stq_18_bits_uop_fp_single;
  reg         stq_18_bits_uop_xcpt_pf_if;
  reg         stq_18_bits_uop_xcpt_ae_if;
  reg         stq_18_bits_uop_xcpt_ma_if;
  reg         stq_18_bits_uop_bp_debug_if;
  reg         stq_18_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_18_bits_uop_debug_fsrc;
  reg  [1:0]  stq_18_bits_uop_debug_tsrc;
  reg         stq_18_bits_addr_valid;
  reg  [39:0] stq_18_bits_addr_bits;
  reg         stq_18_bits_addr_is_virtual;
  reg         stq_18_bits_data_valid;
  reg  [63:0] stq_18_bits_data_bits;
  reg         stq_18_bits_committed;
  reg         stq_18_bits_succeeded;
  reg         stq_19_valid;
  reg  [6:0]  stq_19_bits_uop_uopc;
  reg  [31:0] stq_19_bits_uop_inst;
  reg  [31:0] stq_19_bits_uop_debug_inst;
  reg         stq_19_bits_uop_is_rvc;
  reg  [39:0] stq_19_bits_uop_debug_pc;
  reg  [2:0]  stq_19_bits_uop_iq_type;
  reg  [9:0]  stq_19_bits_uop_fu_code;
  reg  [3:0]  stq_19_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_19_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_19_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_19_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_19_bits_uop_ctrl_op_fcn;
  reg         stq_19_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_19_bits_uop_ctrl_csr_cmd;
  reg         stq_19_bits_uop_ctrl_is_load;
  reg         stq_19_bits_uop_ctrl_is_sta;
  reg         stq_19_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_19_bits_uop_iw_state;
  reg         stq_19_bits_uop_iw_p1_poisoned;
  reg         stq_19_bits_uop_iw_p2_poisoned;
  reg         stq_19_bits_uop_is_br;
  reg         stq_19_bits_uop_is_jalr;
  reg         stq_19_bits_uop_is_jal;
  reg         stq_19_bits_uop_is_sfb;
  reg  [19:0] stq_19_bits_uop_br_mask;
  reg  [4:0]  stq_19_bits_uop_br_tag;
  reg  [5:0]  stq_19_bits_uop_ftq_idx;
  reg         stq_19_bits_uop_edge_inst;
  reg  [5:0]  stq_19_bits_uop_pc_lob;
  reg         stq_19_bits_uop_taken;
  reg  [19:0] stq_19_bits_uop_imm_packed;
  reg  [11:0] stq_19_bits_uop_csr_addr;
  reg  [6:0]  stq_19_bits_uop_rob_idx;
  reg  [4:0]  stq_19_bits_uop_ldq_idx;
  reg  [4:0]  stq_19_bits_uop_stq_idx;
  reg  [1:0]  stq_19_bits_uop_rxq_idx;
  reg  [6:0]  stq_19_bits_uop_pdst;
  reg  [6:0]  stq_19_bits_uop_prs1;
  reg  [6:0]  stq_19_bits_uop_prs2;
  reg  [6:0]  stq_19_bits_uop_prs3;
  reg  [5:0]  stq_19_bits_uop_ppred;
  reg         stq_19_bits_uop_prs1_busy;
  reg         stq_19_bits_uop_prs2_busy;
  reg         stq_19_bits_uop_prs3_busy;
  reg         stq_19_bits_uop_ppred_busy;
  reg  [6:0]  stq_19_bits_uop_stale_pdst;
  reg         stq_19_bits_uop_exception;
  reg  [63:0] stq_19_bits_uop_exc_cause;
  reg         stq_19_bits_uop_bypassable;
  reg  [4:0]  stq_19_bits_uop_mem_cmd;
  reg  [1:0]  stq_19_bits_uop_mem_size;
  reg         stq_19_bits_uop_mem_signed;
  reg         stq_19_bits_uop_is_fence;
  reg         stq_19_bits_uop_is_fencei;
  reg         stq_19_bits_uop_is_amo;
  reg         stq_19_bits_uop_uses_ldq;
  reg         stq_19_bits_uop_uses_stq;
  reg         stq_19_bits_uop_is_sys_pc2epc;
  reg         stq_19_bits_uop_is_unique;
  reg         stq_19_bits_uop_flush_on_commit;
  reg         stq_19_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_19_bits_uop_ldst;
  reg  [5:0]  stq_19_bits_uop_lrs1;
  reg  [5:0]  stq_19_bits_uop_lrs2;
  reg  [5:0]  stq_19_bits_uop_lrs3;
  reg         stq_19_bits_uop_ldst_val;
  reg  [1:0]  stq_19_bits_uop_dst_rtype;
  reg  [1:0]  stq_19_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_19_bits_uop_lrs2_rtype;
  reg         stq_19_bits_uop_frs3_en;
  reg         stq_19_bits_uop_fp_val;
  reg         stq_19_bits_uop_fp_single;
  reg         stq_19_bits_uop_xcpt_pf_if;
  reg         stq_19_bits_uop_xcpt_ae_if;
  reg         stq_19_bits_uop_xcpt_ma_if;
  reg         stq_19_bits_uop_bp_debug_if;
  reg         stq_19_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_19_bits_uop_debug_fsrc;
  reg  [1:0]  stq_19_bits_uop_debug_tsrc;
  reg         stq_19_bits_addr_valid;
  reg  [39:0] stq_19_bits_addr_bits;
  reg         stq_19_bits_addr_is_virtual;
  reg         stq_19_bits_data_valid;
  reg  [63:0] stq_19_bits_data_bits;
  reg         stq_19_bits_committed;
  reg         stq_19_bits_succeeded;
  reg         stq_20_valid;
  reg  [6:0]  stq_20_bits_uop_uopc;
  reg  [31:0] stq_20_bits_uop_inst;
  reg  [31:0] stq_20_bits_uop_debug_inst;
  reg         stq_20_bits_uop_is_rvc;
  reg  [39:0] stq_20_bits_uop_debug_pc;
  reg  [2:0]  stq_20_bits_uop_iq_type;
  reg  [9:0]  stq_20_bits_uop_fu_code;
  reg  [3:0]  stq_20_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_20_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_20_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_20_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_20_bits_uop_ctrl_op_fcn;
  reg         stq_20_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_20_bits_uop_ctrl_csr_cmd;
  reg         stq_20_bits_uop_ctrl_is_load;
  reg         stq_20_bits_uop_ctrl_is_sta;
  reg         stq_20_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_20_bits_uop_iw_state;
  reg         stq_20_bits_uop_iw_p1_poisoned;
  reg         stq_20_bits_uop_iw_p2_poisoned;
  reg         stq_20_bits_uop_is_br;
  reg         stq_20_bits_uop_is_jalr;
  reg         stq_20_bits_uop_is_jal;
  reg         stq_20_bits_uop_is_sfb;
  reg  [19:0] stq_20_bits_uop_br_mask;
  reg  [4:0]  stq_20_bits_uop_br_tag;
  reg  [5:0]  stq_20_bits_uop_ftq_idx;
  reg         stq_20_bits_uop_edge_inst;
  reg  [5:0]  stq_20_bits_uop_pc_lob;
  reg         stq_20_bits_uop_taken;
  reg  [19:0] stq_20_bits_uop_imm_packed;
  reg  [11:0] stq_20_bits_uop_csr_addr;
  reg  [6:0]  stq_20_bits_uop_rob_idx;
  reg  [4:0]  stq_20_bits_uop_ldq_idx;
  reg  [4:0]  stq_20_bits_uop_stq_idx;
  reg  [1:0]  stq_20_bits_uop_rxq_idx;
  reg  [6:0]  stq_20_bits_uop_pdst;
  reg  [6:0]  stq_20_bits_uop_prs1;
  reg  [6:0]  stq_20_bits_uop_prs2;
  reg  [6:0]  stq_20_bits_uop_prs3;
  reg  [5:0]  stq_20_bits_uop_ppred;
  reg         stq_20_bits_uop_prs1_busy;
  reg         stq_20_bits_uop_prs2_busy;
  reg         stq_20_bits_uop_prs3_busy;
  reg         stq_20_bits_uop_ppred_busy;
  reg  [6:0]  stq_20_bits_uop_stale_pdst;
  reg         stq_20_bits_uop_exception;
  reg  [63:0] stq_20_bits_uop_exc_cause;
  reg         stq_20_bits_uop_bypassable;
  reg  [4:0]  stq_20_bits_uop_mem_cmd;
  reg  [1:0]  stq_20_bits_uop_mem_size;
  reg         stq_20_bits_uop_mem_signed;
  reg         stq_20_bits_uop_is_fence;
  reg         stq_20_bits_uop_is_fencei;
  reg         stq_20_bits_uop_is_amo;
  reg         stq_20_bits_uop_uses_ldq;
  reg         stq_20_bits_uop_uses_stq;
  reg         stq_20_bits_uop_is_sys_pc2epc;
  reg         stq_20_bits_uop_is_unique;
  reg         stq_20_bits_uop_flush_on_commit;
  reg         stq_20_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_20_bits_uop_ldst;
  reg  [5:0]  stq_20_bits_uop_lrs1;
  reg  [5:0]  stq_20_bits_uop_lrs2;
  reg  [5:0]  stq_20_bits_uop_lrs3;
  reg         stq_20_bits_uop_ldst_val;
  reg  [1:0]  stq_20_bits_uop_dst_rtype;
  reg  [1:0]  stq_20_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_20_bits_uop_lrs2_rtype;
  reg         stq_20_bits_uop_frs3_en;
  reg         stq_20_bits_uop_fp_val;
  reg         stq_20_bits_uop_fp_single;
  reg         stq_20_bits_uop_xcpt_pf_if;
  reg         stq_20_bits_uop_xcpt_ae_if;
  reg         stq_20_bits_uop_xcpt_ma_if;
  reg         stq_20_bits_uop_bp_debug_if;
  reg         stq_20_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_20_bits_uop_debug_fsrc;
  reg  [1:0]  stq_20_bits_uop_debug_tsrc;
  reg         stq_20_bits_addr_valid;
  reg  [39:0] stq_20_bits_addr_bits;
  reg         stq_20_bits_addr_is_virtual;
  reg         stq_20_bits_data_valid;
  reg  [63:0] stq_20_bits_data_bits;
  reg         stq_20_bits_committed;
  reg         stq_20_bits_succeeded;
  reg         stq_21_valid;
  reg  [6:0]  stq_21_bits_uop_uopc;
  reg  [31:0] stq_21_bits_uop_inst;
  reg  [31:0] stq_21_bits_uop_debug_inst;
  reg         stq_21_bits_uop_is_rvc;
  reg  [39:0] stq_21_bits_uop_debug_pc;
  reg  [2:0]  stq_21_bits_uop_iq_type;
  reg  [9:0]  stq_21_bits_uop_fu_code;
  reg  [3:0]  stq_21_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_21_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_21_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_21_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_21_bits_uop_ctrl_op_fcn;
  reg         stq_21_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_21_bits_uop_ctrl_csr_cmd;
  reg         stq_21_bits_uop_ctrl_is_load;
  reg         stq_21_bits_uop_ctrl_is_sta;
  reg         stq_21_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_21_bits_uop_iw_state;
  reg         stq_21_bits_uop_iw_p1_poisoned;
  reg         stq_21_bits_uop_iw_p2_poisoned;
  reg         stq_21_bits_uop_is_br;
  reg         stq_21_bits_uop_is_jalr;
  reg         stq_21_bits_uop_is_jal;
  reg         stq_21_bits_uop_is_sfb;
  reg  [19:0] stq_21_bits_uop_br_mask;
  reg  [4:0]  stq_21_bits_uop_br_tag;
  reg  [5:0]  stq_21_bits_uop_ftq_idx;
  reg         stq_21_bits_uop_edge_inst;
  reg  [5:0]  stq_21_bits_uop_pc_lob;
  reg         stq_21_bits_uop_taken;
  reg  [19:0] stq_21_bits_uop_imm_packed;
  reg  [11:0] stq_21_bits_uop_csr_addr;
  reg  [6:0]  stq_21_bits_uop_rob_idx;
  reg  [4:0]  stq_21_bits_uop_ldq_idx;
  reg  [4:0]  stq_21_bits_uop_stq_idx;
  reg  [1:0]  stq_21_bits_uop_rxq_idx;
  reg  [6:0]  stq_21_bits_uop_pdst;
  reg  [6:0]  stq_21_bits_uop_prs1;
  reg  [6:0]  stq_21_bits_uop_prs2;
  reg  [6:0]  stq_21_bits_uop_prs3;
  reg  [5:0]  stq_21_bits_uop_ppred;
  reg         stq_21_bits_uop_prs1_busy;
  reg         stq_21_bits_uop_prs2_busy;
  reg         stq_21_bits_uop_prs3_busy;
  reg         stq_21_bits_uop_ppred_busy;
  reg  [6:0]  stq_21_bits_uop_stale_pdst;
  reg         stq_21_bits_uop_exception;
  reg  [63:0] stq_21_bits_uop_exc_cause;
  reg         stq_21_bits_uop_bypassable;
  reg  [4:0]  stq_21_bits_uop_mem_cmd;
  reg  [1:0]  stq_21_bits_uop_mem_size;
  reg         stq_21_bits_uop_mem_signed;
  reg         stq_21_bits_uop_is_fence;
  reg         stq_21_bits_uop_is_fencei;
  reg         stq_21_bits_uop_is_amo;
  reg         stq_21_bits_uop_uses_ldq;
  reg         stq_21_bits_uop_uses_stq;
  reg         stq_21_bits_uop_is_sys_pc2epc;
  reg         stq_21_bits_uop_is_unique;
  reg         stq_21_bits_uop_flush_on_commit;
  reg         stq_21_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_21_bits_uop_ldst;
  reg  [5:0]  stq_21_bits_uop_lrs1;
  reg  [5:0]  stq_21_bits_uop_lrs2;
  reg  [5:0]  stq_21_bits_uop_lrs3;
  reg         stq_21_bits_uop_ldst_val;
  reg  [1:0]  stq_21_bits_uop_dst_rtype;
  reg  [1:0]  stq_21_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_21_bits_uop_lrs2_rtype;
  reg         stq_21_bits_uop_frs3_en;
  reg         stq_21_bits_uop_fp_val;
  reg         stq_21_bits_uop_fp_single;
  reg         stq_21_bits_uop_xcpt_pf_if;
  reg         stq_21_bits_uop_xcpt_ae_if;
  reg         stq_21_bits_uop_xcpt_ma_if;
  reg         stq_21_bits_uop_bp_debug_if;
  reg         stq_21_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_21_bits_uop_debug_fsrc;
  reg  [1:0]  stq_21_bits_uop_debug_tsrc;
  reg         stq_21_bits_addr_valid;
  reg  [39:0] stq_21_bits_addr_bits;
  reg         stq_21_bits_addr_is_virtual;
  reg         stq_21_bits_data_valid;
  reg  [63:0] stq_21_bits_data_bits;
  reg         stq_21_bits_committed;
  reg         stq_21_bits_succeeded;
  reg         stq_22_valid;
  reg  [6:0]  stq_22_bits_uop_uopc;
  reg  [31:0] stq_22_bits_uop_inst;
  reg  [31:0] stq_22_bits_uop_debug_inst;
  reg         stq_22_bits_uop_is_rvc;
  reg  [39:0] stq_22_bits_uop_debug_pc;
  reg  [2:0]  stq_22_bits_uop_iq_type;
  reg  [9:0]  stq_22_bits_uop_fu_code;
  reg  [3:0]  stq_22_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_22_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_22_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_22_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_22_bits_uop_ctrl_op_fcn;
  reg         stq_22_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_22_bits_uop_ctrl_csr_cmd;
  reg         stq_22_bits_uop_ctrl_is_load;
  reg         stq_22_bits_uop_ctrl_is_sta;
  reg         stq_22_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_22_bits_uop_iw_state;
  reg         stq_22_bits_uop_iw_p1_poisoned;
  reg         stq_22_bits_uop_iw_p2_poisoned;
  reg         stq_22_bits_uop_is_br;
  reg         stq_22_bits_uop_is_jalr;
  reg         stq_22_bits_uop_is_jal;
  reg         stq_22_bits_uop_is_sfb;
  reg  [19:0] stq_22_bits_uop_br_mask;
  reg  [4:0]  stq_22_bits_uop_br_tag;
  reg  [5:0]  stq_22_bits_uop_ftq_idx;
  reg         stq_22_bits_uop_edge_inst;
  reg  [5:0]  stq_22_bits_uop_pc_lob;
  reg         stq_22_bits_uop_taken;
  reg  [19:0] stq_22_bits_uop_imm_packed;
  reg  [11:0] stq_22_bits_uop_csr_addr;
  reg  [6:0]  stq_22_bits_uop_rob_idx;
  reg  [4:0]  stq_22_bits_uop_ldq_idx;
  reg  [4:0]  stq_22_bits_uop_stq_idx;
  reg  [1:0]  stq_22_bits_uop_rxq_idx;
  reg  [6:0]  stq_22_bits_uop_pdst;
  reg  [6:0]  stq_22_bits_uop_prs1;
  reg  [6:0]  stq_22_bits_uop_prs2;
  reg  [6:0]  stq_22_bits_uop_prs3;
  reg  [5:0]  stq_22_bits_uop_ppred;
  reg         stq_22_bits_uop_prs1_busy;
  reg         stq_22_bits_uop_prs2_busy;
  reg         stq_22_bits_uop_prs3_busy;
  reg         stq_22_bits_uop_ppred_busy;
  reg  [6:0]  stq_22_bits_uop_stale_pdst;
  reg         stq_22_bits_uop_exception;
  reg  [63:0] stq_22_bits_uop_exc_cause;
  reg         stq_22_bits_uop_bypassable;
  reg  [4:0]  stq_22_bits_uop_mem_cmd;
  reg  [1:0]  stq_22_bits_uop_mem_size;
  reg         stq_22_bits_uop_mem_signed;
  reg         stq_22_bits_uop_is_fence;
  reg         stq_22_bits_uop_is_fencei;
  reg         stq_22_bits_uop_is_amo;
  reg         stq_22_bits_uop_uses_ldq;
  reg         stq_22_bits_uop_uses_stq;
  reg         stq_22_bits_uop_is_sys_pc2epc;
  reg         stq_22_bits_uop_is_unique;
  reg         stq_22_bits_uop_flush_on_commit;
  reg         stq_22_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_22_bits_uop_ldst;
  reg  [5:0]  stq_22_bits_uop_lrs1;
  reg  [5:0]  stq_22_bits_uop_lrs2;
  reg  [5:0]  stq_22_bits_uop_lrs3;
  reg         stq_22_bits_uop_ldst_val;
  reg  [1:0]  stq_22_bits_uop_dst_rtype;
  reg  [1:0]  stq_22_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_22_bits_uop_lrs2_rtype;
  reg         stq_22_bits_uop_frs3_en;
  reg         stq_22_bits_uop_fp_val;
  reg         stq_22_bits_uop_fp_single;
  reg         stq_22_bits_uop_xcpt_pf_if;
  reg         stq_22_bits_uop_xcpt_ae_if;
  reg         stq_22_bits_uop_xcpt_ma_if;
  reg         stq_22_bits_uop_bp_debug_if;
  reg         stq_22_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_22_bits_uop_debug_fsrc;
  reg  [1:0]  stq_22_bits_uop_debug_tsrc;
  reg         stq_22_bits_addr_valid;
  reg  [39:0] stq_22_bits_addr_bits;
  reg         stq_22_bits_addr_is_virtual;
  reg         stq_22_bits_data_valid;
  reg  [63:0] stq_22_bits_data_bits;
  reg         stq_22_bits_committed;
  reg         stq_22_bits_succeeded;
  reg         stq_23_valid;
  reg  [6:0]  stq_23_bits_uop_uopc;
  reg  [31:0] stq_23_bits_uop_inst;
  reg  [31:0] stq_23_bits_uop_debug_inst;
  reg         stq_23_bits_uop_is_rvc;
  reg  [39:0] stq_23_bits_uop_debug_pc;
  reg  [2:0]  stq_23_bits_uop_iq_type;
  reg  [9:0]  stq_23_bits_uop_fu_code;
  reg  [3:0]  stq_23_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_23_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_23_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_23_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_23_bits_uop_ctrl_op_fcn;
  reg         stq_23_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_23_bits_uop_ctrl_csr_cmd;
  reg         stq_23_bits_uop_ctrl_is_load;
  reg         stq_23_bits_uop_ctrl_is_sta;
  reg         stq_23_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_23_bits_uop_iw_state;
  reg         stq_23_bits_uop_iw_p1_poisoned;
  reg         stq_23_bits_uop_iw_p2_poisoned;
  reg         stq_23_bits_uop_is_br;
  reg         stq_23_bits_uop_is_jalr;
  reg         stq_23_bits_uop_is_jal;
  reg         stq_23_bits_uop_is_sfb;
  reg  [19:0] stq_23_bits_uop_br_mask;
  reg  [4:0]  stq_23_bits_uop_br_tag;
  reg  [5:0]  stq_23_bits_uop_ftq_idx;
  reg         stq_23_bits_uop_edge_inst;
  reg  [5:0]  stq_23_bits_uop_pc_lob;
  reg         stq_23_bits_uop_taken;
  reg  [19:0] stq_23_bits_uop_imm_packed;
  reg  [11:0] stq_23_bits_uop_csr_addr;
  reg  [6:0]  stq_23_bits_uop_rob_idx;
  reg  [4:0]  stq_23_bits_uop_ldq_idx;
  reg  [4:0]  stq_23_bits_uop_stq_idx;
  reg  [1:0]  stq_23_bits_uop_rxq_idx;
  reg  [6:0]  stq_23_bits_uop_pdst;
  reg  [6:0]  stq_23_bits_uop_prs1;
  reg  [6:0]  stq_23_bits_uop_prs2;
  reg  [6:0]  stq_23_bits_uop_prs3;
  reg  [5:0]  stq_23_bits_uop_ppred;
  reg         stq_23_bits_uop_prs1_busy;
  reg         stq_23_bits_uop_prs2_busy;
  reg         stq_23_bits_uop_prs3_busy;
  reg         stq_23_bits_uop_ppred_busy;
  reg  [6:0]  stq_23_bits_uop_stale_pdst;
  reg         stq_23_bits_uop_exception;
  reg  [63:0] stq_23_bits_uop_exc_cause;
  reg         stq_23_bits_uop_bypassable;
  reg  [4:0]  stq_23_bits_uop_mem_cmd;
  reg  [1:0]  stq_23_bits_uop_mem_size;
  reg         stq_23_bits_uop_mem_signed;
  reg         stq_23_bits_uop_is_fence;
  reg         stq_23_bits_uop_is_fencei;
  reg         stq_23_bits_uop_is_amo;
  reg         stq_23_bits_uop_uses_ldq;
  reg         stq_23_bits_uop_uses_stq;
  reg         stq_23_bits_uop_is_sys_pc2epc;
  reg         stq_23_bits_uop_is_unique;
  reg         stq_23_bits_uop_flush_on_commit;
  reg         stq_23_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_23_bits_uop_ldst;
  reg  [5:0]  stq_23_bits_uop_lrs1;
  reg  [5:0]  stq_23_bits_uop_lrs2;
  reg  [5:0]  stq_23_bits_uop_lrs3;
  reg         stq_23_bits_uop_ldst_val;
  reg  [1:0]  stq_23_bits_uop_dst_rtype;
  reg  [1:0]  stq_23_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_23_bits_uop_lrs2_rtype;
  reg         stq_23_bits_uop_frs3_en;
  reg         stq_23_bits_uop_fp_val;
  reg         stq_23_bits_uop_fp_single;
  reg         stq_23_bits_uop_xcpt_pf_if;
  reg         stq_23_bits_uop_xcpt_ae_if;
  reg         stq_23_bits_uop_xcpt_ma_if;
  reg         stq_23_bits_uop_bp_debug_if;
  reg         stq_23_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_23_bits_uop_debug_fsrc;
  reg  [1:0]  stq_23_bits_uop_debug_tsrc;
  reg         stq_23_bits_addr_valid;
  reg  [39:0] stq_23_bits_addr_bits;
  reg         stq_23_bits_addr_is_virtual;
  reg         stq_23_bits_data_valid;
  reg  [63:0] stq_23_bits_data_bits;
  reg         stq_23_bits_committed;
  reg         stq_23_bits_succeeded;
  reg         stq_24_valid;
  reg  [6:0]  stq_24_bits_uop_uopc;
  reg  [31:0] stq_24_bits_uop_inst;
  reg  [31:0] stq_24_bits_uop_debug_inst;
  reg         stq_24_bits_uop_is_rvc;
  reg  [39:0] stq_24_bits_uop_debug_pc;
  reg  [2:0]  stq_24_bits_uop_iq_type;
  reg  [9:0]  stq_24_bits_uop_fu_code;
  reg  [3:0]  stq_24_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_24_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_24_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_24_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_24_bits_uop_ctrl_op_fcn;
  reg         stq_24_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_24_bits_uop_ctrl_csr_cmd;
  reg         stq_24_bits_uop_ctrl_is_load;
  reg         stq_24_bits_uop_ctrl_is_sta;
  reg         stq_24_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_24_bits_uop_iw_state;
  reg         stq_24_bits_uop_iw_p1_poisoned;
  reg         stq_24_bits_uop_iw_p2_poisoned;
  reg         stq_24_bits_uop_is_br;
  reg         stq_24_bits_uop_is_jalr;
  reg         stq_24_bits_uop_is_jal;
  reg         stq_24_bits_uop_is_sfb;
  reg  [19:0] stq_24_bits_uop_br_mask;
  reg  [4:0]  stq_24_bits_uop_br_tag;
  reg  [5:0]  stq_24_bits_uop_ftq_idx;
  reg         stq_24_bits_uop_edge_inst;
  reg  [5:0]  stq_24_bits_uop_pc_lob;
  reg         stq_24_bits_uop_taken;
  reg  [19:0] stq_24_bits_uop_imm_packed;
  reg  [11:0] stq_24_bits_uop_csr_addr;
  reg  [6:0]  stq_24_bits_uop_rob_idx;
  reg  [4:0]  stq_24_bits_uop_ldq_idx;
  reg  [4:0]  stq_24_bits_uop_stq_idx;
  reg  [1:0]  stq_24_bits_uop_rxq_idx;
  reg  [6:0]  stq_24_bits_uop_pdst;
  reg  [6:0]  stq_24_bits_uop_prs1;
  reg  [6:0]  stq_24_bits_uop_prs2;
  reg  [6:0]  stq_24_bits_uop_prs3;
  reg  [5:0]  stq_24_bits_uop_ppred;
  reg         stq_24_bits_uop_prs1_busy;
  reg         stq_24_bits_uop_prs2_busy;
  reg         stq_24_bits_uop_prs3_busy;
  reg         stq_24_bits_uop_ppred_busy;
  reg  [6:0]  stq_24_bits_uop_stale_pdst;
  reg         stq_24_bits_uop_exception;
  reg  [63:0] stq_24_bits_uop_exc_cause;
  reg         stq_24_bits_uop_bypassable;
  reg  [4:0]  stq_24_bits_uop_mem_cmd;
  reg  [1:0]  stq_24_bits_uop_mem_size;
  reg         stq_24_bits_uop_mem_signed;
  reg         stq_24_bits_uop_is_fence;
  reg         stq_24_bits_uop_is_fencei;
  reg         stq_24_bits_uop_is_amo;
  reg         stq_24_bits_uop_uses_ldq;
  reg         stq_24_bits_uop_uses_stq;
  reg         stq_24_bits_uop_is_sys_pc2epc;
  reg         stq_24_bits_uop_is_unique;
  reg         stq_24_bits_uop_flush_on_commit;
  reg         stq_24_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_24_bits_uop_ldst;
  reg  [5:0]  stq_24_bits_uop_lrs1;
  reg  [5:0]  stq_24_bits_uop_lrs2;
  reg  [5:0]  stq_24_bits_uop_lrs3;
  reg         stq_24_bits_uop_ldst_val;
  reg  [1:0]  stq_24_bits_uop_dst_rtype;
  reg  [1:0]  stq_24_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_24_bits_uop_lrs2_rtype;
  reg         stq_24_bits_uop_frs3_en;
  reg         stq_24_bits_uop_fp_val;
  reg         stq_24_bits_uop_fp_single;
  reg         stq_24_bits_uop_xcpt_pf_if;
  reg         stq_24_bits_uop_xcpt_ae_if;
  reg         stq_24_bits_uop_xcpt_ma_if;
  reg         stq_24_bits_uop_bp_debug_if;
  reg         stq_24_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_24_bits_uop_debug_fsrc;
  reg  [1:0]  stq_24_bits_uop_debug_tsrc;
  reg         stq_24_bits_addr_valid;
  reg  [39:0] stq_24_bits_addr_bits;
  reg         stq_24_bits_addr_is_virtual;
  reg         stq_24_bits_data_valid;
  reg  [63:0] stq_24_bits_data_bits;
  reg         stq_24_bits_committed;
  reg         stq_24_bits_succeeded;
  reg         stq_25_valid;
  reg  [6:0]  stq_25_bits_uop_uopc;
  reg  [31:0] stq_25_bits_uop_inst;
  reg  [31:0] stq_25_bits_uop_debug_inst;
  reg         stq_25_bits_uop_is_rvc;
  reg  [39:0] stq_25_bits_uop_debug_pc;
  reg  [2:0]  stq_25_bits_uop_iq_type;
  reg  [9:0]  stq_25_bits_uop_fu_code;
  reg  [3:0]  stq_25_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_25_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_25_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_25_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_25_bits_uop_ctrl_op_fcn;
  reg         stq_25_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_25_bits_uop_ctrl_csr_cmd;
  reg         stq_25_bits_uop_ctrl_is_load;
  reg         stq_25_bits_uop_ctrl_is_sta;
  reg         stq_25_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_25_bits_uop_iw_state;
  reg         stq_25_bits_uop_iw_p1_poisoned;
  reg         stq_25_bits_uop_iw_p2_poisoned;
  reg         stq_25_bits_uop_is_br;
  reg         stq_25_bits_uop_is_jalr;
  reg         stq_25_bits_uop_is_jal;
  reg         stq_25_bits_uop_is_sfb;
  reg  [19:0] stq_25_bits_uop_br_mask;
  reg  [4:0]  stq_25_bits_uop_br_tag;
  reg  [5:0]  stq_25_bits_uop_ftq_idx;
  reg         stq_25_bits_uop_edge_inst;
  reg  [5:0]  stq_25_bits_uop_pc_lob;
  reg         stq_25_bits_uop_taken;
  reg  [19:0] stq_25_bits_uop_imm_packed;
  reg  [11:0] stq_25_bits_uop_csr_addr;
  reg  [6:0]  stq_25_bits_uop_rob_idx;
  reg  [4:0]  stq_25_bits_uop_ldq_idx;
  reg  [4:0]  stq_25_bits_uop_stq_idx;
  reg  [1:0]  stq_25_bits_uop_rxq_idx;
  reg  [6:0]  stq_25_bits_uop_pdst;
  reg  [6:0]  stq_25_bits_uop_prs1;
  reg  [6:0]  stq_25_bits_uop_prs2;
  reg  [6:0]  stq_25_bits_uop_prs3;
  reg  [5:0]  stq_25_bits_uop_ppred;
  reg         stq_25_bits_uop_prs1_busy;
  reg         stq_25_bits_uop_prs2_busy;
  reg         stq_25_bits_uop_prs3_busy;
  reg         stq_25_bits_uop_ppred_busy;
  reg  [6:0]  stq_25_bits_uop_stale_pdst;
  reg         stq_25_bits_uop_exception;
  reg  [63:0] stq_25_bits_uop_exc_cause;
  reg         stq_25_bits_uop_bypassable;
  reg  [4:0]  stq_25_bits_uop_mem_cmd;
  reg  [1:0]  stq_25_bits_uop_mem_size;
  reg         stq_25_bits_uop_mem_signed;
  reg         stq_25_bits_uop_is_fence;
  reg         stq_25_bits_uop_is_fencei;
  reg         stq_25_bits_uop_is_amo;
  reg         stq_25_bits_uop_uses_ldq;
  reg         stq_25_bits_uop_uses_stq;
  reg         stq_25_bits_uop_is_sys_pc2epc;
  reg         stq_25_bits_uop_is_unique;
  reg         stq_25_bits_uop_flush_on_commit;
  reg         stq_25_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_25_bits_uop_ldst;
  reg  [5:0]  stq_25_bits_uop_lrs1;
  reg  [5:0]  stq_25_bits_uop_lrs2;
  reg  [5:0]  stq_25_bits_uop_lrs3;
  reg         stq_25_bits_uop_ldst_val;
  reg  [1:0]  stq_25_bits_uop_dst_rtype;
  reg  [1:0]  stq_25_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_25_bits_uop_lrs2_rtype;
  reg         stq_25_bits_uop_frs3_en;
  reg         stq_25_bits_uop_fp_val;
  reg         stq_25_bits_uop_fp_single;
  reg         stq_25_bits_uop_xcpt_pf_if;
  reg         stq_25_bits_uop_xcpt_ae_if;
  reg         stq_25_bits_uop_xcpt_ma_if;
  reg         stq_25_bits_uop_bp_debug_if;
  reg         stq_25_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_25_bits_uop_debug_fsrc;
  reg  [1:0]  stq_25_bits_uop_debug_tsrc;
  reg         stq_25_bits_addr_valid;
  reg  [39:0] stq_25_bits_addr_bits;
  reg         stq_25_bits_addr_is_virtual;
  reg         stq_25_bits_data_valid;
  reg  [63:0] stq_25_bits_data_bits;
  reg         stq_25_bits_committed;
  reg         stq_25_bits_succeeded;
  reg         stq_26_valid;
  reg  [6:0]  stq_26_bits_uop_uopc;
  reg  [31:0] stq_26_bits_uop_inst;
  reg  [31:0] stq_26_bits_uop_debug_inst;
  reg         stq_26_bits_uop_is_rvc;
  reg  [39:0] stq_26_bits_uop_debug_pc;
  reg  [2:0]  stq_26_bits_uop_iq_type;
  reg  [9:0]  stq_26_bits_uop_fu_code;
  reg  [3:0]  stq_26_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_26_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_26_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_26_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_26_bits_uop_ctrl_op_fcn;
  reg         stq_26_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_26_bits_uop_ctrl_csr_cmd;
  reg         stq_26_bits_uop_ctrl_is_load;
  reg         stq_26_bits_uop_ctrl_is_sta;
  reg         stq_26_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_26_bits_uop_iw_state;
  reg         stq_26_bits_uop_iw_p1_poisoned;
  reg         stq_26_bits_uop_iw_p2_poisoned;
  reg         stq_26_bits_uop_is_br;
  reg         stq_26_bits_uop_is_jalr;
  reg         stq_26_bits_uop_is_jal;
  reg         stq_26_bits_uop_is_sfb;
  reg  [19:0] stq_26_bits_uop_br_mask;
  reg  [4:0]  stq_26_bits_uop_br_tag;
  reg  [5:0]  stq_26_bits_uop_ftq_idx;
  reg         stq_26_bits_uop_edge_inst;
  reg  [5:0]  stq_26_bits_uop_pc_lob;
  reg         stq_26_bits_uop_taken;
  reg  [19:0] stq_26_bits_uop_imm_packed;
  reg  [11:0] stq_26_bits_uop_csr_addr;
  reg  [6:0]  stq_26_bits_uop_rob_idx;
  reg  [4:0]  stq_26_bits_uop_ldq_idx;
  reg  [4:0]  stq_26_bits_uop_stq_idx;
  reg  [1:0]  stq_26_bits_uop_rxq_idx;
  reg  [6:0]  stq_26_bits_uop_pdst;
  reg  [6:0]  stq_26_bits_uop_prs1;
  reg  [6:0]  stq_26_bits_uop_prs2;
  reg  [6:0]  stq_26_bits_uop_prs3;
  reg  [5:0]  stq_26_bits_uop_ppred;
  reg         stq_26_bits_uop_prs1_busy;
  reg         stq_26_bits_uop_prs2_busy;
  reg         stq_26_bits_uop_prs3_busy;
  reg         stq_26_bits_uop_ppred_busy;
  reg  [6:0]  stq_26_bits_uop_stale_pdst;
  reg         stq_26_bits_uop_exception;
  reg  [63:0] stq_26_bits_uop_exc_cause;
  reg         stq_26_bits_uop_bypassable;
  reg  [4:0]  stq_26_bits_uop_mem_cmd;
  reg  [1:0]  stq_26_bits_uop_mem_size;
  reg         stq_26_bits_uop_mem_signed;
  reg         stq_26_bits_uop_is_fence;
  reg         stq_26_bits_uop_is_fencei;
  reg         stq_26_bits_uop_is_amo;
  reg         stq_26_bits_uop_uses_ldq;
  reg         stq_26_bits_uop_uses_stq;
  reg         stq_26_bits_uop_is_sys_pc2epc;
  reg         stq_26_bits_uop_is_unique;
  reg         stq_26_bits_uop_flush_on_commit;
  reg         stq_26_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_26_bits_uop_ldst;
  reg  [5:0]  stq_26_bits_uop_lrs1;
  reg  [5:0]  stq_26_bits_uop_lrs2;
  reg  [5:0]  stq_26_bits_uop_lrs3;
  reg         stq_26_bits_uop_ldst_val;
  reg  [1:0]  stq_26_bits_uop_dst_rtype;
  reg  [1:0]  stq_26_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_26_bits_uop_lrs2_rtype;
  reg         stq_26_bits_uop_frs3_en;
  reg         stq_26_bits_uop_fp_val;
  reg         stq_26_bits_uop_fp_single;
  reg         stq_26_bits_uop_xcpt_pf_if;
  reg         stq_26_bits_uop_xcpt_ae_if;
  reg         stq_26_bits_uop_xcpt_ma_if;
  reg         stq_26_bits_uop_bp_debug_if;
  reg         stq_26_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_26_bits_uop_debug_fsrc;
  reg  [1:0]  stq_26_bits_uop_debug_tsrc;
  reg         stq_26_bits_addr_valid;
  reg  [39:0] stq_26_bits_addr_bits;
  reg         stq_26_bits_addr_is_virtual;
  reg         stq_26_bits_data_valid;
  reg  [63:0] stq_26_bits_data_bits;
  reg         stq_26_bits_committed;
  reg         stq_26_bits_succeeded;
  reg         stq_27_valid;
  reg  [6:0]  stq_27_bits_uop_uopc;
  reg  [31:0] stq_27_bits_uop_inst;
  reg  [31:0] stq_27_bits_uop_debug_inst;
  reg         stq_27_bits_uop_is_rvc;
  reg  [39:0] stq_27_bits_uop_debug_pc;
  reg  [2:0]  stq_27_bits_uop_iq_type;
  reg  [9:0]  stq_27_bits_uop_fu_code;
  reg  [3:0]  stq_27_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_27_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_27_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_27_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_27_bits_uop_ctrl_op_fcn;
  reg         stq_27_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_27_bits_uop_ctrl_csr_cmd;
  reg         stq_27_bits_uop_ctrl_is_load;
  reg         stq_27_bits_uop_ctrl_is_sta;
  reg         stq_27_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_27_bits_uop_iw_state;
  reg         stq_27_bits_uop_iw_p1_poisoned;
  reg         stq_27_bits_uop_iw_p2_poisoned;
  reg         stq_27_bits_uop_is_br;
  reg         stq_27_bits_uop_is_jalr;
  reg         stq_27_bits_uop_is_jal;
  reg         stq_27_bits_uop_is_sfb;
  reg  [19:0] stq_27_bits_uop_br_mask;
  reg  [4:0]  stq_27_bits_uop_br_tag;
  reg  [5:0]  stq_27_bits_uop_ftq_idx;
  reg         stq_27_bits_uop_edge_inst;
  reg  [5:0]  stq_27_bits_uop_pc_lob;
  reg         stq_27_bits_uop_taken;
  reg  [19:0] stq_27_bits_uop_imm_packed;
  reg  [11:0] stq_27_bits_uop_csr_addr;
  reg  [6:0]  stq_27_bits_uop_rob_idx;
  reg  [4:0]  stq_27_bits_uop_ldq_idx;
  reg  [4:0]  stq_27_bits_uop_stq_idx;
  reg  [1:0]  stq_27_bits_uop_rxq_idx;
  reg  [6:0]  stq_27_bits_uop_pdst;
  reg  [6:0]  stq_27_bits_uop_prs1;
  reg  [6:0]  stq_27_bits_uop_prs2;
  reg  [6:0]  stq_27_bits_uop_prs3;
  reg  [5:0]  stq_27_bits_uop_ppred;
  reg         stq_27_bits_uop_prs1_busy;
  reg         stq_27_bits_uop_prs2_busy;
  reg         stq_27_bits_uop_prs3_busy;
  reg         stq_27_bits_uop_ppred_busy;
  reg  [6:0]  stq_27_bits_uop_stale_pdst;
  reg         stq_27_bits_uop_exception;
  reg  [63:0] stq_27_bits_uop_exc_cause;
  reg         stq_27_bits_uop_bypassable;
  reg  [4:0]  stq_27_bits_uop_mem_cmd;
  reg  [1:0]  stq_27_bits_uop_mem_size;
  reg         stq_27_bits_uop_mem_signed;
  reg         stq_27_bits_uop_is_fence;
  reg         stq_27_bits_uop_is_fencei;
  reg         stq_27_bits_uop_is_amo;
  reg         stq_27_bits_uop_uses_ldq;
  reg         stq_27_bits_uop_uses_stq;
  reg         stq_27_bits_uop_is_sys_pc2epc;
  reg         stq_27_bits_uop_is_unique;
  reg         stq_27_bits_uop_flush_on_commit;
  reg         stq_27_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_27_bits_uop_ldst;
  reg  [5:0]  stq_27_bits_uop_lrs1;
  reg  [5:0]  stq_27_bits_uop_lrs2;
  reg  [5:0]  stq_27_bits_uop_lrs3;
  reg         stq_27_bits_uop_ldst_val;
  reg  [1:0]  stq_27_bits_uop_dst_rtype;
  reg  [1:0]  stq_27_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_27_bits_uop_lrs2_rtype;
  reg         stq_27_bits_uop_frs3_en;
  reg         stq_27_bits_uop_fp_val;
  reg         stq_27_bits_uop_fp_single;
  reg         stq_27_bits_uop_xcpt_pf_if;
  reg         stq_27_bits_uop_xcpt_ae_if;
  reg         stq_27_bits_uop_xcpt_ma_if;
  reg         stq_27_bits_uop_bp_debug_if;
  reg         stq_27_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_27_bits_uop_debug_fsrc;
  reg  [1:0]  stq_27_bits_uop_debug_tsrc;
  reg         stq_27_bits_addr_valid;
  reg  [39:0] stq_27_bits_addr_bits;
  reg         stq_27_bits_addr_is_virtual;
  reg         stq_27_bits_data_valid;
  reg  [63:0] stq_27_bits_data_bits;
  reg         stq_27_bits_committed;
  reg         stq_27_bits_succeeded;
  reg         stq_28_valid;
  reg  [6:0]  stq_28_bits_uop_uopc;
  reg  [31:0] stq_28_bits_uop_inst;
  reg  [31:0] stq_28_bits_uop_debug_inst;
  reg         stq_28_bits_uop_is_rvc;
  reg  [39:0] stq_28_bits_uop_debug_pc;
  reg  [2:0]  stq_28_bits_uop_iq_type;
  reg  [9:0]  stq_28_bits_uop_fu_code;
  reg  [3:0]  stq_28_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_28_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_28_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_28_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_28_bits_uop_ctrl_op_fcn;
  reg         stq_28_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_28_bits_uop_ctrl_csr_cmd;
  reg         stq_28_bits_uop_ctrl_is_load;
  reg         stq_28_bits_uop_ctrl_is_sta;
  reg         stq_28_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_28_bits_uop_iw_state;
  reg         stq_28_bits_uop_iw_p1_poisoned;
  reg         stq_28_bits_uop_iw_p2_poisoned;
  reg         stq_28_bits_uop_is_br;
  reg         stq_28_bits_uop_is_jalr;
  reg         stq_28_bits_uop_is_jal;
  reg         stq_28_bits_uop_is_sfb;
  reg  [19:0] stq_28_bits_uop_br_mask;
  reg  [4:0]  stq_28_bits_uop_br_tag;
  reg  [5:0]  stq_28_bits_uop_ftq_idx;
  reg         stq_28_bits_uop_edge_inst;
  reg  [5:0]  stq_28_bits_uop_pc_lob;
  reg         stq_28_bits_uop_taken;
  reg  [19:0] stq_28_bits_uop_imm_packed;
  reg  [11:0] stq_28_bits_uop_csr_addr;
  reg  [6:0]  stq_28_bits_uop_rob_idx;
  reg  [4:0]  stq_28_bits_uop_ldq_idx;
  reg  [4:0]  stq_28_bits_uop_stq_idx;
  reg  [1:0]  stq_28_bits_uop_rxq_idx;
  reg  [6:0]  stq_28_bits_uop_pdst;
  reg  [6:0]  stq_28_bits_uop_prs1;
  reg  [6:0]  stq_28_bits_uop_prs2;
  reg  [6:0]  stq_28_bits_uop_prs3;
  reg  [5:0]  stq_28_bits_uop_ppred;
  reg         stq_28_bits_uop_prs1_busy;
  reg         stq_28_bits_uop_prs2_busy;
  reg         stq_28_bits_uop_prs3_busy;
  reg         stq_28_bits_uop_ppred_busy;
  reg  [6:0]  stq_28_bits_uop_stale_pdst;
  reg         stq_28_bits_uop_exception;
  reg  [63:0] stq_28_bits_uop_exc_cause;
  reg         stq_28_bits_uop_bypassable;
  reg  [4:0]  stq_28_bits_uop_mem_cmd;
  reg  [1:0]  stq_28_bits_uop_mem_size;
  reg         stq_28_bits_uop_mem_signed;
  reg         stq_28_bits_uop_is_fence;
  reg         stq_28_bits_uop_is_fencei;
  reg         stq_28_bits_uop_is_amo;
  reg         stq_28_bits_uop_uses_ldq;
  reg         stq_28_bits_uop_uses_stq;
  reg         stq_28_bits_uop_is_sys_pc2epc;
  reg         stq_28_bits_uop_is_unique;
  reg         stq_28_bits_uop_flush_on_commit;
  reg         stq_28_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_28_bits_uop_ldst;
  reg  [5:0]  stq_28_bits_uop_lrs1;
  reg  [5:0]  stq_28_bits_uop_lrs2;
  reg  [5:0]  stq_28_bits_uop_lrs3;
  reg         stq_28_bits_uop_ldst_val;
  reg  [1:0]  stq_28_bits_uop_dst_rtype;
  reg  [1:0]  stq_28_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_28_bits_uop_lrs2_rtype;
  reg         stq_28_bits_uop_frs3_en;
  reg         stq_28_bits_uop_fp_val;
  reg         stq_28_bits_uop_fp_single;
  reg         stq_28_bits_uop_xcpt_pf_if;
  reg         stq_28_bits_uop_xcpt_ae_if;
  reg         stq_28_bits_uop_xcpt_ma_if;
  reg         stq_28_bits_uop_bp_debug_if;
  reg         stq_28_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_28_bits_uop_debug_fsrc;
  reg  [1:0]  stq_28_bits_uop_debug_tsrc;
  reg         stq_28_bits_addr_valid;
  reg  [39:0] stq_28_bits_addr_bits;
  reg         stq_28_bits_addr_is_virtual;
  reg         stq_28_bits_data_valid;
  reg  [63:0] stq_28_bits_data_bits;
  reg         stq_28_bits_committed;
  reg         stq_28_bits_succeeded;
  reg         stq_29_valid;
  reg  [6:0]  stq_29_bits_uop_uopc;
  reg  [31:0] stq_29_bits_uop_inst;
  reg  [31:0] stq_29_bits_uop_debug_inst;
  reg         stq_29_bits_uop_is_rvc;
  reg  [39:0] stq_29_bits_uop_debug_pc;
  reg  [2:0]  stq_29_bits_uop_iq_type;
  reg  [9:0]  stq_29_bits_uop_fu_code;
  reg  [3:0]  stq_29_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_29_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_29_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_29_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_29_bits_uop_ctrl_op_fcn;
  reg         stq_29_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_29_bits_uop_ctrl_csr_cmd;
  reg         stq_29_bits_uop_ctrl_is_load;
  reg         stq_29_bits_uop_ctrl_is_sta;
  reg         stq_29_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_29_bits_uop_iw_state;
  reg         stq_29_bits_uop_iw_p1_poisoned;
  reg         stq_29_bits_uop_iw_p2_poisoned;
  reg         stq_29_bits_uop_is_br;
  reg         stq_29_bits_uop_is_jalr;
  reg         stq_29_bits_uop_is_jal;
  reg         stq_29_bits_uop_is_sfb;
  reg  [19:0] stq_29_bits_uop_br_mask;
  reg  [4:0]  stq_29_bits_uop_br_tag;
  reg  [5:0]  stq_29_bits_uop_ftq_idx;
  reg         stq_29_bits_uop_edge_inst;
  reg  [5:0]  stq_29_bits_uop_pc_lob;
  reg         stq_29_bits_uop_taken;
  reg  [19:0] stq_29_bits_uop_imm_packed;
  reg  [11:0] stq_29_bits_uop_csr_addr;
  reg  [6:0]  stq_29_bits_uop_rob_idx;
  reg  [4:0]  stq_29_bits_uop_ldq_idx;
  reg  [4:0]  stq_29_bits_uop_stq_idx;
  reg  [1:0]  stq_29_bits_uop_rxq_idx;
  reg  [6:0]  stq_29_bits_uop_pdst;
  reg  [6:0]  stq_29_bits_uop_prs1;
  reg  [6:0]  stq_29_bits_uop_prs2;
  reg  [6:0]  stq_29_bits_uop_prs3;
  reg  [5:0]  stq_29_bits_uop_ppred;
  reg         stq_29_bits_uop_prs1_busy;
  reg         stq_29_bits_uop_prs2_busy;
  reg         stq_29_bits_uop_prs3_busy;
  reg         stq_29_bits_uop_ppred_busy;
  reg  [6:0]  stq_29_bits_uop_stale_pdst;
  reg         stq_29_bits_uop_exception;
  reg  [63:0] stq_29_bits_uop_exc_cause;
  reg         stq_29_bits_uop_bypassable;
  reg  [4:0]  stq_29_bits_uop_mem_cmd;
  reg  [1:0]  stq_29_bits_uop_mem_size;
  reg         stq_29_bits_uop_mem_signed;
  reg         stq_29_bits_uop_is_fence;
  reg         stq_29_bits_uop_is_fencei;
  reg         stq_29_bits_uop_is_amo;
  reg         stq_29_bits_uop_uses_ldq;
  reg         stq_29_bits_uop_uses_stq;
  reg         stq_29_bits_uop_is_sys_pc2epc;
  reg         stq_29_bits_uop_is_unique;
  reg         stq_29_bits_uop_flush_on_commit;
  reg         stq_29_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_29_bits_uop_ldst;
  reg  [5:0]  stq_29_bits_uop_lrs1;
  reg  [5:0]  stq_29_bits_uop_lrs2;
  reg  [5:0]  stq_29_bits_uop_lrs3;
  reg         stq_29_bits_uop_ldst_val;
  reg  [1:0]  stq_29_bits_uop_dst_rtype;
  reg  [1:0]  stq_29_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_29_bits_uop_lrs2_rtype;
  reg         stq_29_bits_uop_frs3_en;
  reg         stq_29_bits_uop_fp_val;
  reg         stq_29_bits_uop_fp_single;
  reg         stq_29_bits_uop_xcpt_pf_if;
  reg         stq_29_bits_uop_xcpt_ae_if;
  reg         stq_29_bits_uop_xcpt_ma_if;
  reg         stq_29_bits_uop_bp_debug_if;
  reg         stq_29_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_29_bits_uop_debug_fsrc;
  reg  [1:0]  stq_29_bits_uop_debug_tsrc;
  reg         stq_29_bits_addr_valid;
  reg  [39:0] stq_29_bits_addr_bits;
  reg         stq_29_bits_addr_is_virtual;
  reg         stq_29_bits_data_valid;
  reg  [63:0] stq_29_bits_data_bits;
  reg         stq_29_bits_committed;
  reg         stq_29_bits_succeeded;
  reg         stq_30_valid;
  reg  [6:0]  stq_30_bits_uop_uopc;
  reg  [31:0] stq_30_bits_uop_inst;
  reg  [31:0] stq_30_bits_uop_debug_inst;
  reg         stq_30_bits_uop_is_rvc;
  reg  [39:0] stq_30_bits_uop_debug_pc;
  reg  [2:0]  stq_30_bits_uop_iq_type;
  reg  [9:0]  stq_30_bits_uop_fu_code;
  reg  [3:0]  stq_30_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_30_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_30_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_30_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_30_bits_uop_ctrl_op_fcn;
  reg         stq_30_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_30_bits_uop_ctrl_csr_cmd;
  reg         stq_30_bits_uop_ctrl_is_load;
  reg         stq_30_bits_uop_ctrl_is_sta;
  reg         stq_30_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_30_bits_uop_iw_state;
  reg         stq_30_bits_uop_iw_p1_poisoned;
  reg         stq_30_bits_uop_iw_p2_poisoned;
  reg         stq_30_bits_uop_is_br;
  reg         stq_30_bits_uop_is_jalr;
  reg         stq_30_bits_uop_is_jal;
  reg         stq_30_bits_uop_is_sfb;
  reg  [19:0] stq_30_bits_uop_br_mask;
  reg  [4:0]  stq_30_bits_uop_br_tag;
  reg  [5:0]  stq_30_bits_uop_ftq_idx;
  reg         stq_30_bits_uop_edge_inst;
  reg  [5:0]  stq_30_bits_uop_pc_lob;
  reg         stq_30_bits_uop_taken;
  reg  [19:0] stq_30_bits_uop_imm_packed;
  reg  [11:0] stq_30_bits_uop_csr_addr;
  reg  [6:0]  stq_30_bits_uop_rob_idx;
  reg  [4:0]  stq_30_bits_uop_ldq_idx;
  reg  [4:0]  stq_30_bits_uop_stq_idx;
  reg  [1:0]  stq_30_bits_uop_rxq_idx;
  reg  [6:0]  stq_30_bits_uop_pdst;
  reg  [6:0]  stq_30_bits_uop_prs1;
  reg  [6:0]  stq_30_bits_uop_prs2;
  reg  [6:0]  stq_30_bits_uop_prs3;
  reg  [5:0]  stq_30_bits_uop_ppred;
  reg         stq_30_bits_uop_prs1_busy;
  reg         stq_30_bits_uop_prs2_busy;
  reg         stq_30_bits_uop_prs3_busy;
  reg         stq_30_bits_uop_ppred_busy;
  reg  [6:0]  stq_30_bits_uop_stale_pdst;
  reg         stq_30_bits_uop_exception;
  reg  [63:0] stq_30_bits_uop_exc_cause;
  reg         stq_30_bits_uop_bypassable;
  reg  [4:0]  stq_30_bits_uop_mem_cmd;
  reg  [1:0]  stq_30_bits_uop_mem_size;
  reg         stq_30_bits_uop_mem_signed;
  reg         stq_30_bits_uop_is_fence;
  reg         stq_30_bits_uop_is_fencei;
  reg         stq_30_bits_uop_is_amo;
  reg         stq_30_bits_uop_uses_ldq;
  reg         stq_30_bits_uop_uses_stq;
  reg         stq_30_bits_uop_is_sys_pc2epc;
  reg         stq_30_bits_uop_is_unique;
  reg         stq_30_bits_uop_flush_on_commit;
  reg         stq_30_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_30_bits_uop_ldst;
  reg  [5:0]  stq_30_bits_uop_lrs1;
  reg  [5:0]  stq_30_bits_uop_lrs2;
  reg  [5:0]  stq_30_bits_uop_lrs3;
  reg         stq_30_bits_uop_ldst_val;
  reg  [1:0]  stq_30_bits_uop_dst_rtype;
  reg  [1:0]  stq_30_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_30_bits_uop_lrs2_rtype;
  reg         stq_30_bits_uop_frs3_en;
  reg         stq_30_bits_uop_fp_val;
  reg         stq_30_bits_uop_fp_single;
  reg         stq_30_bits_uop_xcpt_pf_if;
  reg         stq_30_bits_uop_xcpt_ae_if;
  reg         stq_30_bits_uop_xcpt_ma_if;
  reg         stq_30_bits_uop_bp_debug_if;
  reg         stq_30_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_30_bits_uop_debug_fsrc;
  reg  [1:0]  stq_30_bits_uop_debug_tsrc;
  reg         stq_30_bits_addr_valid;
  reg  [39:0] stq_30_bits_addr_bits;
  reg         stq_30_bits_addr_is_virtual;
  reg         stq_30_bits_data_valid;
  reg  [63:0] stq_30_bits_data_bits;
  reg         stq_30_bits_committed;
  reg         stq_30_bits_succeeded;
  reg         stq_31_valid;
  reg  [6:0]  stq_31_bits_uop_uopc;
  reg  [31:0] stq_31_bits_uop_inst;
  reg  [31:0] stq_31_bits_uop_debug_inst;
  reg         stq_31_bits_uop_is_rvc;
  reg  [39:0] stq_31_bits_uop_debug_pc;
  reg  [2:0]  stq_31_bits_uop_iq_type;
  reg  [9:0]  stq_31_bits_uop_fu_code;
  reg  [3:0]  stq_31_bits_uop_ctrl_br_type;
  reg  [1:0]  stq_31_bits_uop_ctrl_op1_sel;
  reg  [2:0]  stq_31_bits_uop_ctrl_op2_sel;
  reg  [2:0]  stq_31_bits_uop_ctrl_imm_sel;
  reg  [3:0]  stq_31_bits_uop_ctrl_op_fcn;
  reg         stq_31_bits_uop_ctrl_fcn_dw;
  reg  [2:0]  stq_31_bits_uop_ctrl_csr_cmd;
  reg         stq_31_bits_uop_ctrl_is_load;
  reg         stq_31_bits_uop_ctrl_is_sta;
  reg         stq_31_bits_uop_ctrl_is_std;
  reg  [1:0]  stq_31_bits_uop_iw_state;
  reg         stq_31_bits_uop_iw_p1_poisoned;
  reg         stq_31_bits_uop_iw_p2_poisoned;
  reg         stq_31_bits_uop_is_br;
  reg         stq_31_bits_uop_is_jalr;
  reg         stq_31_bits_uop_is_jal;
  reg         stq_31_bits_uop_is_sfb;
  reg  [19:0] stq_31_bits_uop_br_mask;
  reg  [4:0]  stq_31_bits_uop_br_tag;
  reg  [5:0]  stq_31_bits_uop_ftq_idx;
  reg         stq_31_bits_uop_edge_inst;
  reg  [5:0]  stq_31_bits_uop_pc_lob;
  reg         stq_31_bits_uop_taken;
  reg  [19:0] stq_31_bits_uop_imm_packed;
  reg  [11:0] stq_31_bits_uop_csr_addr;
  reg  [6:0]  stq_31_bits_uop_rob_idx;
  reg  [4:0]  stq_31_bits_uop_ldq_idx;
  reg  [4:0]  stq_31_bits_uop_stq_idx;
  reg  [1:0]  stq_31_bits_uop_rxq_idx;
  reg  [6:0]  stq_31_bits_uop_pdst;
  reg  [6:0]  stq_31_bits_uop_prs1;
  reg  [6:0]  stq_31_bits_uop_prs2;
  reg  [6:0]  stq_31_bits_uop_prs3;
  reg  [5:0]  stq_31_bits_uop_ppred;
  reg         stq_31_bits_uop_prs1_busy;
  reg         stq_31_bits_uop_prs2_busy;
  reg         stq_31_bits_uop_prs3_busy;
  reg         stq_31_bits_uop_ppred_busy;
  reg  [6:0]  stq_31_bits_uop_stale_pdst;
  reg         stq_31_bits_uop_exception;
  reg  [63:0] stq_31_bits_uop_exc_cause;
  reg         stq_31_bits_uop_bypassable;
  reg  [4:0]  stq_31_bits_uop_mem_cmd;
  reg  [1:0]  stq_31_bits_uop_mem_size;
  reg         stq_31_bits_uop_mem_signed;
  reg         stq_31_bits_uop_is_fence;
  reg         stq_31_bits_uop_is_fencei;
  reg         stq_31_bits_uop_is_amo;
  reg         stq_31_bits_uop_uses_ldq;
  reg         stq_31_bits_uop_uses_stq;
  reg         stq_31_bits_uop_is_sys_pc2epc;
  reg         stq_31_bits_uop_is_unique;
  reg         stq_31_bits_uop_flush_on_commit;
  reg         stq_31_bits_uop_ldst_is_rs1;
  reg  [5:0]  stq_31_bits_uop_ldst;
  reg  [5:0]  stq_31_bits_uop_lrs1;
  reg  [5:0]  stq_31_bits_uop_lrs2;
  reg  [5:0]  stq_31_bits_uop_lrs3;
  reg         stq_31_bits_uop_ldst_val;
  reg  [1:0]  stq_31_bits_uop_dst_rtype;
  reg  [1:0]  stq_31_bits_uop_lrs1_rtype;
  reg  [1:0]  stq_31_bits_uop_lrs2_rtype;
  reg         stq_31_bits_uop_frs3_en;
  reg         stq_31_bits_uop_fp_val;
  reg         stq_31_bits_uop_fp_single;
  reg         stq_31_bits_uop_xcpt_pf_if;
  reg         stq_31_bits_uop_xcpt_ae_if;
  reg         stq_31_bits_uop_xcpt_ma_if;
  reg         stq_31_bits_uop_bp_debug_if;
  reg         stq_31_bits_uop_bp_xcpt_if;
  reg  [1:0]  stq_31_bits_uop_debug_fsrc;
  reg  [1:0]  stq_31_bits_uop_debug_tsrc;
  reg         stq_31_bits_addr_valid;
  reg  [39:0] stq_31_bits_addr_bits;
  reg         stq_31_bits_addr_is_virtual;
  reg         stq_31_bits_data_valid;
  reg  [63:0] stq_31_bits_data_bits;
  reg         stq_31_bits_committed;
  reg         stq_31_bits_succeeded;
  reg  [4:0]  ldq_head;
  reg  [4:0]  ldq_tail;
  reg  [4:0]  stq_head;
  reg  [4:0]  stq_tail;
  reg  [4:0]  stq_commit_head;
  reg  [4:0]  stq_execute_head;
  reg         casez_tmp;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp = stq_0_valid;
      5'b00001:
        casez_tmp = stq_1_valid;
      5'b00010:
        casez_tmp = stq_2_valid;
      5'b00011:
        casez_tmp = stq_3_valid;
      5'b00100:
        casez_tmp = stq_4_valid;
      5'b00101:
        casez_tmp = stq_5_valid;
      5'b00110:
        casez_tmp = stq_6_valid;
      5'b00111:
        casez_tmp = stq_7_valid;
      5'b01000:
        casez_tmp = stq_8_valid;
      5'b01001:
        casez_tmp = stq_9_valid;
      5'b01010:
        casez_tmp = stq_10_valid;
      5'b01011:
        casez_tmp = stq_11_valid;
      5'b01100:
        casez_tmp = stq_12_valid;
      5'b01101:
        casez_tmp = stq_13_valid;
      5'b01110:
        casez_tmp = stq_14_valid;
      5'b01111:
        casez_tmp = stq_15_valid;
      5'b10000:
        casez_tmp = stq_16_valid;
      5'b10001:
        casez_tmp = stq_17_valid;
      5'b10010:
        casez_tmp = stq_18_valid;
      5'b10011:
        casez_tmp = stq_19_valid;
      5'b10100:
        casez_tmp = stq_20_valid;
      5'b10101:
        casez_tmp = stq_21_valid;
      5'b10110:
        casez_tmp = stq_22_valid;
      5'b10111:
        casez_tmp = stq_23_valid;
      5'b11000:
        casez_tmp = stq_24_valid;
      5'b11001:
        casez_tmp = stq_25_valid;
      5'b11010:
        casez_tmp = stq_26_valid;
      5'b11011:
        casez_tmp = stq_27_valid;
      5'b11100:
        casez_tmp = stq_28_valid;
      5'b11101:
        casez_tmp = stq_29_valid;
      5'b11110:
        casez_tmp = stq_30_valid;
      default:
        casez_tmp = stq_31_valid;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_0;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_0 = stq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_0 = stq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_0 = stq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_0 = stq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_0 = stq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_0 = stq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_0 = stq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_0 = stq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_0 = stq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_0 = stq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_0 = stq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_0 = stq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_0 = stq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_0 = stq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_0 = stq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_0 = stq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_0 = stq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_0 = stq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_0 = stq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_0 = stq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_0 = stq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_0 = stq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_0 = stq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_0 = stq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_0 = stq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_0 = stq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_0 = stq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_0 = stq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_0 = stq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_0 = stq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_0 = stq_30_bits_uop_uopc;
      default:
        casez_tmp_0 = stq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_1;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_1 = stq_0_bits_uop_inst;
      5'b00001:
        casez_tmp_1 = stq_1_bits_uop_inst;
      5'b00010:
        casez_tmp_1 = stq_2_bits_uop_inst;
      5'b00011:
        casez_tmp_1 = stq_3_bits_uop_inst;
      5'b00100:
        casez_tmp_1 = stq_4_bits_uop_inst;
      5'b00101:
        casez_tmp_1 = stq_5_bits_uop_inst;
      5'b00110:
        casez_tmp_1 = stq_6_bits_uop_inst;
      5'b00111:
        casez_tmp_1 = stq_7_bits_uop_inst;
      5'b01000:
        casez_tmp_1 = stq_8_bits_uop_inst;
      5'b01001:
        casez_tmp_1 = stq_9_bits_uop_inst;
      5'b01010:
        casez_tmp_1 = stq_10_bits_uop_inst;
      5'b01011:
        casez_tmp_1 = stq_11_bits_uop_inst;
      5'b01100:
        casez_tmp_1 = stq_12_bits_uop_inst;
      5'b01101:
        casez_tmp_1 = stq_13_bits_uop_inst;
      5'b01110:
        casez_tmp_1 = stq_14_bits_uop_inst;
      5'b01111:
        casez_tmp_1 = stq_15_bits_uop_inst;
      5'b10000:
        casez_tmp_1 = stq_16_bits_uop_inst;
      5'b10001:
        casez_tmp_1 = stq_17_bits_uop_inst;
      5'b10010:
        casez_tmp_1 = stq_18_bits_uop_inst;
      5'b10011:
        casez_tmp_1 = stq_19_bits_uop_inst;
      5'b10100:
        casez_tmp_1 = stq_20_bits_uop_inst;
      5'b10101:
        casez_tmp_1 = stq_21_bits_uop_inst;
      5'b10110:
        casez_tmp_1 = stq_22_bits_uop_inst;
      5'b10111:
        casez_tmp_1 = stq_23_bits_uop_inst;
      5'b11000:
        casez_tmp_1 = stq_24_bits_uop_inst;
      5'b11001:
        casez_tmp_1 = stq_25_bits_uop_inst;
      5'b11010:
        casez_tmp_1 = stq_26_bits_uop_inst;
      5'b11011:
        casez_tmp_1 = stq_27_bits_uop_inst;
      5'b11100:
        casez_tmp_1 = stq_28_bits_uop_inst;
      5'b11101:
        casez_tmp_1 = stq_29_bits_uop_inst;
      5'b11110:
        casez_tmp_1 = stq_30_bits_uop_inst;
      default:
        casez_tmp_1 = stq_31_bits_uop_inst;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_2;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_2 = stq_0_bits_uop_debug_inst;
      5'b00001:
        casez_tmp_2 = stq_1_bits_uop_debug_inst;
      5'b00010:
        casez_tmp_2 = stq_2_bits_uop_debug_inst;
      5'b00011:
        casez_tmp_2 = stq_3_bits_uop_debug_inst;
      5'b00100:
        casez_tmp_2 = stq_4_bits_uop_debug_inst;
      5'b00101:
        casez_tmp_2 = stq_5_bits_uop_debug_inst;
      5'b00110:
        casez_tmp_2 = stq_6_bits_uop_debug_inst;
      5'b00111:
        casez_tmp_2 = stq_7_bits_uop_debug_inst;
      5'b01000:
        casez_tmp_2 = stq_8_bits_uop_debug_inst;
      5'b01001:
        casez_tmp_2 = stq_9_bits_uop_debug_inst;
      5'b01010:
        casez_tmp_2 = stq_10_bits_uop_debug_inst;
      5'b01011:
        casez_tmp_2 = stq_11_bits_uop_debug_inst;
      5'b01100:
        casez_tmp_2 = stq_12_bits_uop_debug_inst;
      5'b01101:
        casez_tmp_2 = stq_13_bits_uop_debug_inst;
      5'b01110:
        casez_tmp_2 = stq_14_bits_uop_debug_inst;
      5'b01111:
        casez_tmp_2 = stq_15_bits_uop_debug_inst;
      5'b10000:
        casez_tmp_2 = stq_16_bits_uop_debug_inst;
      5'b10001:
        casez_tmp_2 = stq_17_bits_uop_debug_inst;
      5'b10010:
        casez_tmp_2 = stq_18_bits_uop_debug_inst;
      5'b10011:
        casez_tmp_2 = stq_19_bits_uop_debug_inst;
      5'b10100:
        casez_tmp_2 = stq_20_bits_uop_debug_inst;
      5'b10101:
        casez_tmp_2 = stq_21_bits_uop_debug_inst;
      5'b10110:
        casez_tmp_2 = stq_22_bits_uop_debug_inst;
      5'b10111:
        casez_tmp_2 = stq_23_bits_uop_debug_inst;
      5'b11000:
        casez_tmp_2 = stq_24_bits_uop_debug_inst;
      5'b11001:
        casez_tmp_2 = stq_25_bits_uop_debug_inst;
      5'b11010:
        casez_tmp_2 = stq_26_bits_uop_debug_inst;
      5'b11011:
        casez_tmp_2 = stq_27_bits_uop_debug_inst;
      5'b11100:
        casez_tmp_2 = stq_28_bits_uop_debug_inst;
      5'b11101:
        casez_tmp_2 = stq_29_bits_uop_debug_inst;
      5'b11110:
        casez_tmp_2 = stq_30_bits_uop_debug_inst;
      default:
        casez_tmp_2 = stq_31_bits_uop_debug_inst;
    endcase
  end // always @(*)
  reg         casez_tmp_3;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_3 = stq_0_bits_uop_is_rvc;
      5'b00001:
        casez_tmp_3 = stq_1_bits_uop_is_rvc;
      5'b00010:
        casez_tmp_3 = stq_2_bits_uop_is_rvc;
      5'b00011:
        casez_tmp_3 = stq_3_bits_uop_is_rvc;
      5'b00100:
        casez_tmp_3 = stq_4_bits_uop_is_rvc;
      5'b00101:
        casez_tmp_3 = stq_5_bits_uop_is_rvc;
      5'b00110:
        casez_tmp_3 = stq_6_bits_uop_is_rvc;
      5'b00111:
        casez_tmp_3 = stq_7_bits_uop_is_rvc;
      5'b01000:
        casez_tmp_3 = stq_8_bits_uop_is_rvc;
      5'b01001:
        casez_tmp_3 = stq_9_bits_uop_is_rvc;
      5'b01010:
        casez_tmp_3 = stq_10_bits_uop_is_rvc;
      5'b01011:
        casez_tmp_3 = stq_11_bits_uop_is_rvc;
      5'b01100:
        casez_tmp_3 = stq_12_bits_uop_is_rvc;
      5'b01101:
        casez_tmp_3 = stq_13_bits_uop_is_rvc;
      5'b01110:
        casez_tmp_3 = stq_14_bits_uop_is_rvc;
      5'b01111:
        casez_tmp_3 = stq_15_bits_uop_is_rvc;
      5'b10000:
        casez_tmp_3 = stq_16_bits_uop_is_rvc;
      5'b10001:
        casez_tmp_3 = stq_17_bits_uop_is_rvc;
      5'b10010:
        casez_tmp_3 = stq_18_bits_uop_is_rvc;
      5'b10011:
        casez_tmp_3 = stq_19_bits_uop_is_rvc;
      5'b10100:
        casez_tmp_3 = stq_20_bits_uop_is_rvc;
      5'b10101:
        casez_tmp_3 = stq_21_bits_uop_is_rvc;
      5'b10110:
        casez_tmp_3 = stq_22_bits_uop_is_rvc;
      5'b10111:
        casez_tmp_3 = stq_23_bits_uop_is_rvc;
      5'b11000:
        casez_tmp_3 = stq_24_bits_uop_is_rvc;
      5'b11001:
        casez_tmp_3 = stq_25_bits_uop_is_rvc;
      5'b11010:
        casez_tmp_3 = stq_26_bits_uop_is_rvc;
      5'b11011:
        casez_tmp_3 = stq_27_bits_uop_is_rvc;
      5'b11100:
        casez_tmp_3 = stq_28_bits_uop_is_rvc;
      5'b11101:
        casez_tmp_3 = stq_29_bits_uop_is_rvc;
      5'b11110:
        casez_tmp_3 = stq_30_bits_uop_is_rvc;
      default:
        casez_tmp_3 = stq_31_bits_uop_is_rvc;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_4;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_4 = stq_0_bits_uop_debug_pc;
      5'b00001:
        casez_tmp_4 = stq_1_bits_uop_debug_pc;
      5'b00010:
        casez_tmp_4 = stq_2_bits_uop_debug_pc;
      5'b00011:
        casez_tmp_4 = stq_3_bits_uop_debug_pc;
      5'b00100:
        casez_tmp_4 = stq_4_bits_uop_debug_pc;
      5'b00101:
        casez_tmp_4 = stq_5_bits_uop_debug_pc;
      5'b00110:
        casez_tmp_4 = stq_6_bits_uop_debug_pc;
      5'b00111:
        casez_tmp_4 = stq_7_bits_uop_debug_pc;
      5'b01000:
        casez_tmp_4 = stq_8_bits_uop_debug_pc;
      5'b01001:
        casez_tmp_4 = stq_9_bits_uop_debug_pc;
      5'b01010:
        casez_tmp_4 = stq_10_bits_uop_debug_pc;
      5'b01011:
        casez_tmp_4 = stq_11_bits_uop_debug_pc;
      5'b01100:
        casez_tmp_4 = stq_12_bits_uop_debug_pc;
      5'b01101:
        casez_tmp_4 = stq_13_bits_uop_debug_pc;
      5'b01110:
        casez_tmp_4 = stq_14_bits_uop_debug_pc;
      5'b01111:
        casez_tmp_4 = stq_15_bits_uop_debug_pc;
      5'b10000:
        casez_tmp_4 = stq_16_bits_uop_debug_pc;
      5'b10001:
        casez_tmp_4 = stq_17_bits_uop_debug_pc;
      5'b10010:
        casez_tmp_4 = stq_18_bits_uop_debug_pc;
      5'b10011:
        casez_tmp_4 = stq_19_bits_uop_debug_pc;
      5'b10100:
        casez_tmp_4 = stq_20_bits_uop_debug_pc;
      5'b10101:
        casez_tmp_4 = stq_21_bits_uop_debug_pc;
      5'b10110:
        casez_tmp_4 = stq_22_bits_uop_debug_pc;
      5'b10111:
        casez_tmp_4 = stq_23_bits_uop_debug_pc;
      5'b11000:
        casez_tmp_4 = stq_24_bits_uop_debug_pc;
      5'b11001:
        casez_tmp_4 = stq_25_bits_uop_debug_pc;
      5'b11010:
        casez_tmp_4 = stq_26_bits_uop_debug_pc;
      5'b11011:
        casez_tmp_4 = stq_27_bits_uop_debug_pc;
      5'b11100:
        casez_tmp_4 = stq_28_bits_uop_debug_pc;
      5'b11101:
        casez_tmp_4 = stq_29_bits_uop_debug_pc;
      5'b11110:
        casez_tmp_4 = stq_30_bits_uop_debug_pc;
      default:
        casez_tmp_4 = stq_31_bits_uop_debug_pc;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_5;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_5 = stq_0_bits_uop_iq_type;
      5'b00001:
        casez_tmp_5 = stq_1_bits_uop_iq_type;
      5'b00010:
        casez_tmp_5 = stq_2_bits_uop_iq_type;
      5'b00011:
        casez_tmp_5 = stq_3_bits_uop_iq_type;
      5'b00100:
        casez_tmp_5 = stq_4_bits_uop_iq_type;
      5'b00101:
        casez_tmp_5 = stq_5_bits_uop_iq_type;
      5'b00110:
        casez_tmp_5 = stq_6_bits_uop_iq_type;
      5'b00111:
        casez_tmp_5 = stq_7_bits_uop_iq_type;
      5'b01000:
        casez_tmp_5 = stq_8_bits_uop_iq_type;
      5'b01001:
        casez_tmp_5 = stq_9_bits_uop_iq_type;
      5'b01010:
        casez_tmp_5 = stq_10_bits_uop_iq_type;
      5'b01011:
        casez_tmp_5 = stq_11_bits_uop_iq_type;
      5'b01100:
        casez_tmp_5 = stq_12_bits_uop_iq_type;
      5'b01101:
        casez_tmp_5 = stq_13_bits_uop_iq_type;
      5'b01110:
        casez_tmp_5 = stq_14_bits_uop_iq_type;
      5'b01111:
        casez_tmp_5 = stq_15_bits_uop_iq_type;
      5'b10000:
        casez_tmp_5 = stq_16_bits_uop_iq_type;
      5'b10001:
        casez_tmp_5 = stq_17_bits_uop_iq_type;
      5'b10010:
        casez_tmp_5 = stq_18_bits_uop_iq_type;
      5'b10011:
        casez_tmp_5 = stq_19_bits_uop_iq_type;
      5'b10100:
        casez_tmp_5 = stq_20_bits_uop_iq_type;
      5'b10101:
        casez_tmp_5 = stq_21_bits_uop_iq_type;
      5'b10110:
        casez_tmp_5 = stq_22_bits_uop_iq_type;
      5'b10111:
        casez_tmp_5 = stq_23_bits_uop_iq_type;
      5'b11000:
        casez_tmp_5 = stq_24_bits_uop_iq_type;
      5'b11001:
        casez_tmp_5 = stq_25_bits_uop_iq_type;
      5'b11010:
        casez_tmp_5 = stq_26_bits_uop_iq_type;
      5'b11011:
        casez_tmp_5 = stq_27_bits_uop_iq_type;
      5'b11100:
        casez_tmp_5 = stq_28_bits_uop_iq_type;
      5'b11101:
        casez_tmp_5 = stq_29_bits_uop_iq_type;
      5'b11110:
        casez_tmp_5 = stq_30_bits_uop_iq_type;
      default:
        casez_tmp_5 = stq_31_bits_uop_iq_type;
    endcase
  end // always @(*)
  reg  [9:0]  casez_tmp_6;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_6 = stq_0_bits_uop_fu_code;
      5'b00001:
        casez_tmp_6 = stq_1_bits_uop_fu_code;
      5'b00010:
        casez_tmp_6 = stq_2_bits_uop_fu_code;
      5'b00011:
        casez_tmp_6 = stq_3_bits_uop_fu_code;
      5'b00100:
        casez_tmp_6 = stq_4_bits_uop_fu_code;
      5'b00101:
        casez_tmp_6 = stq_5_bits_uop_fu_code;
      5'b00110:
        casez_tmp_6 = stq_6_bits_uop_fu_code;
      5'b00111:
        casez_tmp_6 = stq_7_bits_uop_fu_code;
      5'b01000:
        casez_tmp_6 = stq_8_bits_uop_fu_code;
      5'b01001:
        casez_tmp_6 = stq_9_bits_uop_fu_code;
      5'b01010:
        casez_tmp_6 = stq_10_bits_uop_fu_code;
      5'b01011:
        casez_tmp_6 = stq_11_bits_uop_fu_code;
      5'b01100:
        casez_tmp_6 = stq_12_bits_uop_fu_code;
      5'b01101:
        casez_tmp_6 = stq_13_bits_uop_fu_code;
      5'b01110:
        casez_tmp_6 = stq_14_bits_uop_fu_code;
      5'b01111:
        casez_tmp_6 = stq_15_bits_uop_fu_code;
      5'b10000:
        casez_tmp_6 = stq_16_bits_uop_fu_code;
      5'b10001:
        casez_tmp_6 = stq_17_bits_uop_fu_code;
      5'b10010:
        casez_tmp_6 = stq_18_bits_uop_fu_code;
      5'b10011:
        casez_tmp_6 = stq_19_bits_uop_fu_code;
      5'b10100:
        casez_tmp_6 = stq_20_bits_uop_fu_code;
      5'b10101:
        casez_tmp_6 = stq_21_bits_uop_fu_code;
      5'b10110:
        casez_tmp_6 = stq_22_bits_uop_fu_code;
      5'b10111:
        casez_tmp_6 = stq_23_bits_uop_fu_code;
      5'b11000:
        casez_tmp_6 = stq_24_bits_uop_fu_code;
      5'b11001:
        casez_tmp_6 = stq_25_bits_uop_fu_code;
      5'b11010:
        casez_tmp_6 = stq_26_bits_uop_fu_code;
      5'b11011:
        casez_tmp_6 = stq_27_bits_uop_fu_code;
      5'b11100:
        casez_tmp_6 = stq_28_bits_uop_fu_code;
      5'b11101:
        casez_tmp_6 = stq_29_bits_uop_fu_code;
      5'b11110:
        casez_tmp_6 = stq_30_bits_uop_fu_code;
      default:
        casez_tmp_6 = stq_31_bits_uop_fu_code;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_7;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_7 = stq_0_bits_uop_ctrl_br_type;
      5'b00001:
        casez_tmp_7 = stq_1_bits_uop_ctrl_br_type;
      5'b00010:
        casez_tmp_7 = stq_2_bits_uop_ctrl_br_type;
      5'b00011:
        casez_tmp_7 = stq_3_bits_uop_ctrl_br_type;
      5'b00100:
        casez_tmp_7 = stq_4_bits_uop_ctrl_br_type;
      5'b00101:
        casez_tmp_7 = stq_5_bits_uop_ctrl_br_type;
      5'b00110:
        casez_tmp_7 = stq_6_bits_uop_ctrl_br_type;
      5'b00111:
        casez_tmp_7 = stq_7_bits_uop_ctrl_br_type;
      5'b01000:
        casez_tmp_7 = stq_8_bits_uop_ctrl_br_type;
      5'b01001:
        casez_tmp_7 = stq_9_bits_uop_ctrl_br_type;
      5'b01010:
        casez_tmp_7 = stq_10_bits_uop_ctrl_br_type;
      5'b01011:
        casez_tmp_7 = stq_11_bits_uop_ctrl_br_type;
      5'b01100:
        casez_tmp_7 = stq_12_bits_uop_ctrl_br_type;
      5'b01101:
        casez_tmp_7 = stq_13_bits_uop_ctrl_br_type;
      5'b01110:
        casez_tmp_7 = stq_14_bits_uop_ctrl_br_type;
      5'b01111:
        casez_tmp_7 = stq_15_bits_uop_ctrl_br_type;
      5'b10000:
        casez_tmp_7 = stq_16_bits_uop_ctrl_br_type;
      5'b10001:
        casez_tmp_7 = stq_17_bits_uop_ctrl_br_type;
      5'b10010:
        casez_tmp_7 = stq_18_bits_uop_ctrl_br_type;
      5'b10011:
        casez_tmp_7 = stq_19_bits_uop_ctrl_br_type;
      5'b10100:
        casez_tmp_7 = stq_20_bits_uop_ctrl_br_type;
      5'b10101:
        casez_tmp_7 = stq_21_bits_uop_ctrl_br_type;
      5'b10110:
        casez_tmp_7 = stq_22_bits_uop_ctrl_br_type;
      5'b10111:
        casez_tmp_7 = stq_23_bits_uop_ctrl_br_type;
      5'b11000:
        casez_tmp_7 = stq_24_bits_uop_ctrl_br_type;
      5'b11001:
        casez_tmp_7 = stq_25_bits_uop_ctrl_br_type;
      5'b11010:
        casez_tmp_7 = stq_26_bits_uop_ctrl_br_type;
      5'b11011:
        casez_tmp_7 = stq_27_bits_uop_ctrl_br_type;
      5'b11100:
        casez_tmp_7 = stq_28_bits_uop_ctrl_br_type;
      5'b11101:
        casez_tmp_7 = stq_29_bits_uop_ctrl_br_type;
      5'b11110:
        casez_tmp_7 = stq_30_bits_uop_ctrl_br_type;
      default:
        casez_tmp_7 = stq_31_bits_uop_ctrl_br_type;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_8;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_8 = stq_0_bits_uop_ctrl_op1_sel;
      5'b00001:
        casez_tmp_8 = stq_1_bits_uop_ctrl_op1_sel;
      5'b00010:
        casez_tmp_8 = stq_2_bits_uop_ctrl_op1_sel;
      5'b00011:
        casez_tmp_8 = stq_3_bits_uop_ctrl_op1_sel;
      5'b00100:
        casez_tmp_8 = stq_4_bits_uop_ctrl_op1_sel;
      5'b00101:
        casez_tmp_8 = stq_5_bits_uop_ctrl_op1_sel;
      5'b00110:
        casez_tmp_8 = stq_6_bits_uop_ctrl_op1_sel;
      5'b00111:
        casez_tmp_8 = stq_7_bits_uop_ctrl_op1_sel;
      5'b01000:
        casez_tmp_8 = stq_8_bits_uop_ctrl_op1_sel;
      5'b01001:
        casez_tmp_8 = stq_9_bits_uop_ctrl_op1_sel;
      5'b01010:
        casez_tmp_8 = stq_10_bits_uop_ctrl_op1_sel;
      5'b01011:
        casez_tmp_8 = stq_11_bits_uop_ctrl_op1_sel;
      5'b01100:
        casez_tmp_8 = stq_12_bits_uop_ctrl_op1_sel;
      5'b01101:
        casez_tmp_8 = stq_13_bits_uop_ctrl_op1_sel;
      5'b01110:
        casez_tmp_8 = stq_14_bits_uop_ctrl_op1_sel;
      5'b01111:
        casez_tmp_8 = stq_15_bits_uop_ctrl_op1_sel;
      5'b10000:
        casez_tmp_8 = stq_16_bits_uop_ctrl_op1_sel;
      5'b10001:
        casez_tmp_8 = stq_17_bits_uop_ctrl_op1_sel;
      5'b10010:
        casez_tmp_8 = stq_18_bits_uop_ctrl_op1_sel;
      5'b10011:
        casez_tmp_8 = stq_19_bits_uop_ctrl_op1_sel;
      5'b10100:
        casez_tmp_8 = stq_20_bits_uop_ctrl_op1_sel;
      5'b10101:
        casez_tmp_8 = stq_21_bits_uop_ctrl_op1_sel;
      5'b10110:
        casez_tmp_8 = stq_22_bits_uop_ctrl_op1_sel;
      5'b10111:
        casez_tmp_8 = stq_23_bits_uop_ctrl_op1_sel;
      5'b11000:
        casez_tmp_8 = stq_24_bits_uop_ctrl_op1_sel;
      5'b11001:
        casez_tmp_8 = stq_25_bits_uop_ctrl_op1_sel;
      5'b11010:
        casez_tmp_8 = stq_26_bits_uop_ctrl_op1_sel;
      5'b11011:
        casez_tmp_8 = stq_27_bits_uop_ctrl_op1_sel;
      5'b11100:
        casez_tmp_8 = stq_28_bits_uop_ctrl_op1_sel;
      5'b11101:
        casez_tmp_8 = stq_29_bits_uop_ctrl_op1_sel;
      5'b11110:
        casez_tmp_8 = stq_30_bits_uop_ctrl_op1_sel;
      default:
        casez_tmp_8 = stq_31_bits_uop_ctrl_op1_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_9;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_9 = stq_0_bits_uop_ctrl_op2_sel;
      5'b00001:
        casez_tmp_9 = stq_1_bits_uop_ctrl_op2_sel;
      5'b00010:
        casez_tmp_9 = stq_2_bits_uop_ctrl_op2_sel;
      5'b00011:
        casez_tmp_9 = stq_3_bits_uop_ctrl_op2_sel;
      5'b00100:
        casez_tmp_9 = stq_4_bits_uop_ctrl_op2_sel;
      5'b00101:
        casez_tmp_9 = stq_5_bits_uop_ctrl_op2_sel;
      5'b00110:
        casez_tmp_9 = stq_6_bits_uop_ctrl_op2_sel;
      5'b00111:
        casez_tmp_9 = stq_7_bits_uop_ctrl_op2_sel;
      5'b01000:
        casez_tmp_9 = stq_8_bits_uop_ctrl_op2_sel;
      5'b01001:
        casez_tmp_9 = stq_9_bits_uop_ctrl_op2_sel;
      5'b01010:
        casez_tmp_9 = stq_10_bits_uop_ctrl_op2_sel;
      5'b01011:
        casez_tmp_9 = stq_11_bits_uop_ctrl_op2_sel;
      5'b01100:
        casez_tmp_9 = stq_12_bits_uop_ctrl_op2_sel;
      5'b01101:
        casez_tmp_9 = stq_13_bits_uop_ctrl_op2_sel;
      5'b01110:
        casez_tmp_9 = stq_14_bits_uop_ctrl_op2_sel;
      5'b01111:
        casez_tmp_9 = stq_15_bits_uop_ctrl_op2_sel;
      5'b10000:
        casez_tmp_9 = stq_16_bits_uop_ctrl_op2_sel;
      5'b10001:
        casez_tmp_9 = stq_17_bits_uop_ctrl_op2_sel;
      5'b10010:
        casez_tmp_9 = stq_18_bits_uop_ctrl_op2_sel;
      5'b10011:
        casez_tmp_9 = stq_19_bits_uop_ctrl_op2_sel;
      5'b10100:
        casez_tmp_9 = stq_20_bits_uop_ctrl_op2_sel;
      5'b10101:
        casez_tmp_9 = stq_21_bits_uop_ctrl_op2_sel;
      5'b10110:
        casez_tmp_9 = stq_22_bits_uop_ctrl_op2_sel;
      5'b10111:
        casez_tmp_9 = stq_23_bits_uop_ctrl_op2_sel;
      5'b11000:
        casez_tmp_9 = stq_24_bits_uop_ctrl_op2_sel;
      5'b11001:
        casez_tmp_9 = stq_25_bits_uop_ctrl_op2_sel;
      5'b11010:
        casez_tmp_9 = stq_26_bits_uop_ctrl_op2_sel;
      5'b11011:
        casez_tmp_9 = stq_27_bits_uop_ctrl_op2_sel;
      5'b11100:
        casez_tmp_9 = stq_28_bits_uop_ctrl_op2_sel;
      5'b11101:
        casez_tmp_9 = stq_29_bits_uop_ctrl_op2_sel;
      5'b11110:
        casez_tmp_9 = stq_30_bits_uop_ctrl_op2_sel;
      default:
        casez_tmp_9 = stq_31_bits_uop_ctrl_op2_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_10;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_10 = stq_0_bits_uop_ctrl_imm_sel;
      5'b00001:
        casez_tmp_10 = stq_1_bits_uop_ctrl_imm_sel;
      5'b00010:
        casez_tmp_10 = stq_2_bits_uop_ctrl_imm_sel;
      5'b00011:
        casez_tmp_10 = stq_3_bits_uop_ctrl_imm_sel;
      5'b00100:
        casez_tmp_10 = stq_4_bits_uop_ctrl_imm_sel;
      5'b00101:
        casez_tmp_10 = stq_5_bits_uop_ctrl_imm_sel;
      5'b00110:
        casez_tmp_10 = stq_6_bits_uop_ctrl_imm_sel;
      5'b00111:
        casez_tmp_10 = stq_7_bits_uop_ctrl_imm_sel;
      5'b01000:
        casez_tmp_10 = stq_8_bits_uop_ctrl_imm_sel;
      5'b01001:
        casez_tmp_10 = stq_9_bits_uop_ctrl_imm_sel;
      5'b01010:
        casez_tmp_10 = stq_10_bits_uop_ctrl_imm_sel;
      5'b01011:
        casez_tmp_10 = stq_11_bits_uop_ctrl_imm_sel;
      5'b01100:
        casez_tmp_10 = stq_12_bits_uop_ctrl_imm_sel;
      5'b01101:
        casez_tmp_10 = stq_13_bits_uop_ctrl_imm_sel;
      5'b01110:
        casez_tmp_10 = stq_14_bits_uop_ctrl_imm_sel;
      5'b01111:
        casez_tmp_10 = stq_15_bits_uop_ctrl_imm_sel;
      5'b10000:
        casez_tmp_10 = stq_16_bits_uop_ctrl_imm_sel;
      5'b10001:
        casez_tmp_10 = stq_17_bits_uop_ctrl_imm_sel;
      5'b10010:
        casez_tmp_10 = stq_18_bits_uop_ctrl_imm_sel;
      5'b10011:
        casez_tmp_10 = stq_19_bits_uop_ctrl_imm_sel;
      5'b10100:
        casez_tmp_10 = stq_20_bits_uop_ctrl_imm_sel;
      5'b10101:
        casez_tmp_10 = stq_21_bits_uop_ctrl_imm_sel;
      5'b10110:
        casez_tmp_10 = stq_22_bits_uop_ctrl_imm_sel;
      5'b10111:
        casez_tmp_10 = stq_23_bits_uop_ctrl_imm_sel;
      5'b11000:
        casez_tmp_10 = stq_24_bits_uop_ctrl_imm_sel;
      5'b11001:
        casez_tmp_10 = stq_25_bits_uop_ctrl_imm_sel;
      5'b11010:
        casez_tmp_10 = stq_26_bits_uop_ctrl_imm_sel;
      5'b11011:
        casez_tmp_10 = stq_27_bits_uop_ctrl_imm_sel;
      5'b11100:
        casez_tmp_10 = stq_28_bits_uop_ctrl_imm_sel;
      5'b11101:
        casez_tmp_10 = stq_29_bits_uop_ctrl_imm_sel;
      5'b11110:
        casez_tmp_10 = stq_30_bits_uop_ctrl_imm_sel;
      default:
        casez_tmp_10 = stq_31_bits_uop_ctrl_imm_sel;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_11;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_11 = stq_0_bits_uop_ctrl_op_fcn;
      5'b00001:
        casez_tmp_11 = stq_1_bits_uop_ctrl_op_fcn;
      5'b00010:
        casez_tmp_11 = stq_2_bits_uop_ctrl_op_fcn;
      5'b00011:
        casez_tmp_11 = stq_3_bits_uop_ctrl_op_fcn;
      5'b00100:
        casez_tmp_11 = stq_4_bits_uop_ctrl_op_fcn;
      5'b00101:
        casez_tmp_11 = stq_5_bits_uop_ctrl_op_fcn;
      5'b00110:
        casez_tmp_11 = stq_6_bits_uop_ctrl_op_fcn;
      5'b00111:
        casez_tmp_11 = stq_7_bits_uop_ctrl_op_fcn;
      5'b01000:
        casez_tmp_11 = stq_8_bits_uop_ctrl_op_fcn;
      5'b01001:
        casez_tmp_11 = stq_9_bits_uop_ctrl_op_fcn;
      5'b01010:
        casez_tmp_11 = stq_10_bits_uop_ctrl_op_fcn;
      5'b01011:
        casez_tmp_11 = stq_11_bits_uop_ctrl_op_fcn;
      5'b01100:
        casez_tmp_11 = stq_12_bits_uop_ctrl_op_fcn;
      5'b01101:
        casez_tmp_11 = stq_13_bits_uop_ctrl_op_fcn;
      5'b01110:
        casez_tmp_11 = stq_14_bits_uop_ctrl_op_fcn;
      5'b01111:
        casez_tmp_11 = stq_15_bits_uop_ctrl_op_fcn;
      5'b10000:
        casez_tmp_11 = stq_16_bits_uop_ctrl_op_fcn;
      5'b10001:
        casez_tmp_11 = stq_17_bits_uop_ctrl_op_fcn;
      5'b10010:
        casez_tmp_11 = stq_18_bits_uop_ctrl_op_fcn;
      5'b10011:
        casez_tmp_11 = stq_19_bits_uop_ctrl_op_fcn;
      5'b10100:
        casez_tmp_11 = stq_20_bits_uop_ctrl_op_fcn;
      5'b10101:
        casez_tmp_11 = stq_21_bits_uop_ctrl_op_fcn;
      5'b10110:
        casez_tmp_11 = stq_22_bits_uop_ctrl_op_fcn;
      5'b10111:
        casez_tmp_11 = stq_23_bits_uop_ctrl_op_fcn;
      5'b11000:
        casez_tmp_11 = stq_24_bits_uop_ctrl_op_fcn;
      5'b11001:
        casez_tmp_11 = stq_25_bits_uop_ctrl_op_fcn;
      5'b11010:
        casez_tmp_11 = stq_26_bits_uop_ctrl_op_fcn;
      5'b11011:
        casez_tmp_11 = stq_27_bits_uop_ctrl_op_fcn;
      5'b11100:
        casez_tmp_11 = stq_28_bits_uop_ctrl_op_fcn;
      5'b11101:
        casez_tmp_11 = stq_29_bits_uop_ctrl_op_fcn;
      5'b11110:
        casez_tmp_11 = stq_30_bits_uop_ctrl_op_fcn;
      default:
        casez_tmp_11 = stq_31_bits_uop_ctrl_op_fcn;
    endcase
  end // always @(*)
  reg         casez_tmp_12;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_12 = stq_0_bits_uop_ctrl_fcn_dw;
      5'b00001:
        casez_tmp_12 = stq_1_bits_uop_ctrl_fcn_dw;
      5'b00010:
        casez_tmp_12 = stq_2_bits_uop_ctrl_fcn_dw;
      5'b00011:
        casez_tmp_12 = stq_3_bits_uop_ctrl_fcn_dw;
      5'b00100:
        casez_tmp_12 = stq_4_bits_uop_ctrl_fcn_dw;
      5'b00101:
        casez_tmp_12 = stq_5_bits_uop_ctrl_fcn_dw;
      5'b00110:
        casez_tmp_12 = stq_6_bits_uop_ctrl_fcn_dw;
      5'b00111:
        casez_tmp_12 = stq_7_bits_uop_ctrl_fcn_dw;
      5'b01000:
        casez_tmp_12 = stq_8_bits_uop_ctrl_fcn_dw;
      5'b01001:
        casez_tmp_12 = stq_9_bits_uop_ctrl_fcn_dw;
      5'b01010:
        casez_tmp_12 = stq_10_bits_uop_ctrl_fcn_dw;
      5'b01011:
        casez_tmp_12 = stq_11_bits_uop_ctrl_fcn_dw;
      5'b01100:
        casez_tmp_12 = stq_12_bits_uop_ctrl_fcn_dw;
      5'b01101:
        casez_tmp_12 = stq_13_bits_uop_ctrl_fcn_dw;
      5'b01110:
        casez_tmp_12 = stq_14_bits_uop_ctrl_fcn_dw;
      5'b01111:
        casez_tmp_12 = stq_15_bits_uop_ctrl_fcn_dw;
      5'b10000:
        casez_tmp_12 = stq_16_bits_uop_ctrl_fcn_dw;
      5'b10001:
        casez_tmp_12 = stq_17_bits_uop_ctrl_fcn_dw;
      5'b10010:
        casez_tmp_12 = stq_18_bits_uop_ctrl_fcn_dw;
      5'b10011:
        casez_tmp_12 = stq_19_bits_uop_ctrl_fcn_dw;
      5'b10100:
        casez_tmp_12 = stq_20_bits_uop_ctrl_fcn_dw;
      5'b10101:
        casez_tmp_12 = stq_21_bits_uop_ctrl_fcn_dw;
      5'b10110:
        casez_tmp_12 = stq_22_bits_uop_ctrl_fcn_dw;
      5'b10111:
        casez_tmp_12 = stq_23_bits_uop_ctrl_fcn_dw;
      5'b11000:
        casez_tmp_12 = stq_24_bits_uop_ctrl_fcn_dw;
      5'b11001:
        casez_tmp_12 = stq_25_bits_uop_ctrl_fcn_dw;
      5'b11010:
        casez_tmp_12 = stq_26_bits_uop_ctrl_fcn_dw;
      5'b11011:
        casez_tmp_12 = stq_27_bits_uop_ctrl_fcn_dw;
      5'b11100:
        casez_tmp_12 = stq_28_bits_uop_ctrl_fcn_dw;
      5'b11101:
        casez_tmp_12 = stq_29_bits_uop_ctrl_fcn_dw;
      5'b11110:
        casez_tmp_12 = stq_30_bits_uop_ctrl_fcn_dw;
      default:
        casez_tmp_12 = stq_31_bits_uop_ctrl_fcn_dw;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_13;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_13 = stq_0_bits_uop_ctrl_csr_cmd;
      5'b00001:
        casez_tmp_13 = stq_1_bits_uop_ctrl_csr_cmd;
      5'b00010:
        casez_tmp_13 = stq_2_bits_uop_ctrl_csr_cmd;
      5'b00011:
        casez_tmp_13 = stq_3_bits_uop_ctrl_csr_cmd;
      5'b00100:
        casez_tmp_13 = stq_4_bits_uop_ctrl_csr_cmd;
      5'b00101:
        casez_tmp_13 = stq_5_bits_uop_ctrl_csr_cmd;
      5'b00110:
        casez_tmp_13 = stq_6_bits_uop_ctrl_csr_cmd;
      5'b00111:
        casez_tmp_13 = stq_7_bits_uop_ctrl_csr_cmd;
      5'b01000:
        casez_tmp_13 = stq_8_bits_uop_ctrl_csr_cmd;
      5'b01001:
        casez_tmp_13 = stq_9_bits_uop_ctrl_csr_cmd;
      5'b01010:
        casez_tmp_13 = stq_10_bits_uop_ctrl_csr_cmd;
      5'b01011:
        casez_tmp_13 = stq_11_bits_uop_ctrl_csr_cmd;
      5'b01100:
        casez_tmp_13 = stq_12_bits_uop_ctrl_csr_cmd;
      5'b01101:
        casez_tmp_13 = stq_13_bits_uop_ctrl_csr_cmd;
      5'b01110:
        casez_tmp_13 = stq_14_bits_uop_ctrl_csr_cmd;
      5'b01111:
        casez_tmp_13 = stq_15_bits_uop_ctrl_csr_cmd;
      5'b10000:
        casez_tmp_13 = stq_16_bits_uop_ctrl_csr_cmd;
      5'b10001:
        casez_tmp_13 = stq_17_bits_uop_ctrl_csr_cmd;
      5'b10010:
        casez_tmp_13 = stq_18_bits_uop_ctrl_csr_cmd;
      5'b10011:
        casez_tmp_13 = stq_19_bits_uop_ctrl_csr_cmd;
      5'b10100:
        casez_tmp_13 = stq_20_bits_uop_ctrl_csr_cmd;
      5'b10101:
        casez_tmp_13 = stq_21_bits_uop_ctrl_csr_cmd;
      5'b10110:
        casez_tmp_13 = stq_22_bits_uop_ctrl_csr_cmd;
      5'b10111:
        casez_tmp_13 = stq_23_bits_uop_ctrl_csr_cmd;
      5'b11000:
        casez_tmp_13 = stq_24_bits_uop_ctrl_csr_cmd;
      5'b11001:
        casez_tmp_13 = stq_25_bits_uop_ctrl_csr_cmd;
      5'b11010:
        casez_tmp_13 = stq_26_bits_uop_ctrl_csr_cmd;
      5'b11011:
        casez_tmp_13 = stq_27_bits_uop_ctrl_csr_cmd;
      5'b11100:
        casez_tmp_13 = stq_28_bits_uop_ctrl_csr_cmd;
      5'b11101:
        casez_tmp_13 = stq_29_bits_uop_ctrl_csr_cmd;
      5'b11110:
        casez_tmp_13 = stq_30_bits_uop_ctrl_csr_cmd;
      default:
        casez_tmp_13 = stq_31_bits_uop_ctrl_csr_cmd;
    endcase
  end // always @(*)
  reg         casez_tmp_14;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_14 = stq_0_bits_uop_ctrl_is_load;
      5'b00001:
        casez_tmp_14 = stq_1_bits_uop_ctrl_is_load;
      5'b00010:
        casez_tmp_14 = stq_2_bits_uop_ctrl_is_load;
      5'b00011:
        casez_tmp_14 = stq_3_bits_uop_ctrl_is_load;
      5'b00100:
        casez_tmp_14 = stq_4_bits_uop_ctrl_is_load;
      5'b00101:
        casez_tmp_14 = stq_5_bits_uop_ctrl_is_load;
      5'b00110:
        casez_tmp_14 = stq_6_bits_uop_ctrl_is_load;
      5'b00111:
        casez_tmp_14 = stq_7_bits_uop_ctrl_is_load;
      5'b01000:
        casez_tmp_14 = stq_8_bits_uop_ctrl_is_load;
      5'b01001:
        casez_tmp_14 = stq_9_bits_uop_ctrl_is_load;
      5'b01010:
        casez_tmp_14 = stq_10_bits_uop_ctrl_is_load;
      5'b01011:
        casez_tmp_14 = stq_11_bits_uop_ctrl_is_load;
      5'b01100:
        casez_tmp_14 = stq_12_bits_uop_ctrl_is_load;
      5'b01101:
        casez_tmp_14 = stq_13_bits_uop_ctrl_is_load;
      5'b01110:
        casez_tmp_14 = stq_14_bits_uop_ctrl_is_load;
      5'b01111:
        casez_tmp_14 = stq_15_bits_uop_ctrl_is_load;
      5'b10000:
        casez_tmp_14 = stq_16_bits_uop_ctrl_is_load;
      5'b10001:
        casez_tmp_14 = stq_17_bits_uop_ctrl_is_load;
      5'b10010:
        casez_tmp_14 = stq_18_bits_uop_ctrl_is_load;
      5'b10011:
        casez_tmp_14 = stq_19_bits_uop_ctrl_is_load;
      5'b10100:
        casez_tmp_14 = stq_20_bits_uop_ctrl_is_load;
      5'b10101:
        casez_tmp_14 = stq_21_bits_uop_ctrl_is_load;
      5'b10110:
        casez_tmp_14 = stq_22_bits_uop_ctrl_is_load;
      5'b10111:
        casez_tmp_14 = stq_23_bits_uop_ctrl_is_load;
      5'b11000:
        casez_tmp_14 = stq_24_bits_uop_ctrl_is_load;
      5'b11001:
        casez_tmp_14 = stq_25_bits_uop_ctrl_is_load;
      5'b11010:
        casez_tmp_14 = stq_26_bits_uop_ctrl_is_load;
      5'b11011:
        casez_tmp_14 = stq_27_bits_uop_ctrl_is_load;
      5'b11100:
        casez_tmp_14 = stq_28_bits_uop_ctrl_is_load;
      5'b11101:
        casez_tmp_14 = stq_29_bits_uop_ctrl_is_load;
      5'b11110:
        casez_tmp_14 = stq_30_bits_uop_ctrl_is_load;
      default:
        casez_tmp_14 = stq_31_bits_uop_ctrl_is_load;
    endcase
  end // always @(*)
  reg         casez_tmp_15;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_15 = stq_0_bits_uop_ctrl_is_sta;
      5'b00001:
        casez_tmp_15 = stq_1_bits_uop_ctrl_is_sta;
      5'b00010:
        casez_tmp_15 = stq_2_bits_uop_ctrl_is_sta;
      5'b00011:
        casez_tmp_15 = stq_3_bits_uop_ctrl_is_sta;
      5'b00100:
        casez_tmp_15 = stq_4_bits_uop_ctrl_is_sta;
      5'b00101:
        casez_tmp_15 = stq_5_bits_uop_ctrl_is_sta;
      5'b00110:
        casez_tmp_15 = stq_6_bits_uop_ctrl_is_sta;
      5'b00111:
        casez_tmp_15 = stq_7_bits_uop_ctrl_is_sta;
      5'b01000:
        casez_tmp_15 = stq_8_bits_uop_ctrl_is_sta;
      5'b01001:
        casez_tmp_15 = stq_9_bits_uop_ctrl_is_sta;
      5'b01010:
        casez_tmp_15 = stq_10_bits_uop_ctrl_is_sta;
      5'b01011:
        casez_tmp_15 = stq_11_bits_uop_ctrl_is_sta;
      5'b01100:
        casez_tmp_15 = stq_12_bits_uop_ctrl_is_sta;
      5'b01101:
        casez_tmp_15 = stq_13_bits_uop_ctrl_is_sta;
      5'b01110:
        casez_tmp_15 = stq_14_bits_uop_ctrl_is_sta;
      5'b01111:
        casez_tmp_15 = stq_15_bits_uop_ctrl_is_sta;
      5'b10000:
        casez_tmp_15 = stq_16_bits_uop_ctrl_is_sta;
      5'b10001:
        casez_tmp_15 = stq_17_bits_uop_ctrl_is_sta;
      5'b10010:
        casez_tmp_15 = stq_18_bits_uop_ctrl_is_sta;
      5'b10011:
        casez_tmp_15 = stq_19_bits_uop_ctrl_is_sta;
      5'b10100:
        casez_tmp_15 = stq_20_bits_uop_ctrl_is_sta;
      5'b10101:
        casez_tmp_15 = stq_21_bits_uop_ctrl_is_sta;
      5'b10110:
        casez_tmp_15 = stq_22_bits_uop_ctrl_is_sta;
      5'b10111:
        casez_tmp_15 = stq_23_bits_uop_ctrl_is_sta;
      5'b11000:
        casez_tmp_15 = stq_24_bits_uop_ctrl_is_sta;
      5'b11001:
        casez_tmp_15 = stq_25_bits_uop_ctrl_is_sta;
      5'b11010:
        casez_tmp_15 = stq_26_bits_uop_ctrl_is_sta;
      5'b11011:
        casez_tmp_15 = stq_27_bits_uop_ctrl_is_sta;
      5'b11100:
        casez_tmp_15 = stq_28_bits_uop_ctrl_is_sta;
      5'b11101:
        casez_tmp_15 = stq_29_bits_uop_ctrl_is_sta;
      5'b11110:
        casez_tmp_15 = stq_30_bits_uop_ctrl_is_sta;
      default:
        casez_tmp_15 = stq_31_bits_uop_ctrl_is_sta;
    endcase
  end // always @(*)
  reg         casez_tmp_16;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_16 = stq_0_bits_uop_ctrl_is_std;
      5'b00001:
        casez_tmp_16 = stq_1_bits_uop_ctrl_is_std;
      5'b00010:
        casez_tmp_16 = stq_2_bits_uop_ctrl_is_std;
      5'b00011:
        casez_tmp_16 = stq_3_bits_uop_ctrl_is_std;
      5'b00100:
        casez_tmp_16 = stq_4_bits_uop_ctrl_is_std;
      5'b00101:
        casez_tmp_16 = stq_5_bits_uop_ctrl_is_std;
      5'b00110:
        casez_tmp_16 = stq_6_bits_uop_ctrl_is_std;
      5'b00111:
        casez_tmp_16 = stq_7_bits_uop_ctrl_is_std;
      5'b01000:
        casez_tmp_16 = stq_8_bits_uop_ctrl_is_std;
      5'b01001:
        casez_tmp_16 = stq_9_bits_uop_ctrl_is_std;
      5'b01010:
        casez_tmp_16 = stq_10_bits_uop_ctrl_is_std;
      5'b01011:
        casez_tmp_16 = stq_11_bits_uop_ctrl_is_std;
      5'b01100:
        casez_tmp_16 = stq_12_bits_uop_ctrl_is_std;
      5'b01101:
        casez_tmp_16 = stq_13_bits_uop_ctrl_is_std;
      5'b01110:
        casez_tmp_16 = stq_14_bits_uop_ctrl_is_std;
      5'b01111:
        casez_tmp_16 = stq_15_bits_uop_ctrl_is_std;
      5'b10000:
        casez_tmp_16 = stq_16_bits_uop_ctrl_is_std;
      5'b10001:
        casez_tmp_16 = stq_17_bits_uop_ctrl_is_std;
      5'b10010:
        casez_tmp_16 = stq_18_bits_uop_ctrl_is_std;
      5'b10011:
        casez_tmp_16 = stq_19_bits_uop_ctrl_is_std;
      5'b10100:
        casez_tmp_16 = stq_20_bits_uop_ctrl_is_std;
      5'b10101:
        casez_tmp_16 = stq_21_bits_uop_ctrl_is_std;
      5'b10110:
        casez_tmp_16 = stq_22_bits_uop_ctrl_is_std;
      5'b10111:
        casez_tmp_16 = stq_23_bits_uop_ctrl_is_std;
      5'b11000:
        casez_tmp_16 = stq_24_bits_uop_ctrl_is_std;
      5'b11001:
        casez_tmp_16 = stq_25_bits_uop_ctrl_is_std;
      5'b11010:
        casez_tmp_16 = stq_26_bits_uop_ctrl_is_std;
      5'b11011:
        casez_tmp_16 = stq_27_bits_uop_ctrl_is_std;
      5'b11100:
        casez_tmp_16 = stq_28_bits_uop_ctrl_is_std;
      5'b11101:
        casez_tmp_16 = stq_29_bits_uop_ctrl_is_std;
      5'b11110:
        casez_tmp_16 = stq_30_bits_uop_ctrl_is_std;
      default:
        casez_tmp_16 = stq_31_bits_uop_ctrl_is_std;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_17;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_17 = stq_0_bits_uop_iw_state;
      5'b00001:
        casez_tmp_17 = stq_1_bits_uop_iw_state;
      5'b00010:
        casez_tmp_17 = stq_2_bits_uop_iw_state;
      5'b00011:
        casez_tmp_17 = stq_3_bits_uop_iw_state;
      5'b00100:
        casez_tmp_17 = stq_4_bits_uop_iw_state;
      5'b00101:
        casez_tmp_17 = stq_5_bits_uop_iw_state;
      5'b00110:
        casez_tmp_17 = stq_6_bits_uop_iw_state;
      5'b00111:
        casez_tmp_17 = stq_7_bits_uop_iw_state;
      5'b01000:
        casez_tmp_17 = stq_8_bits_uop_iw_state;
      5'b01001:
        casez_tmp_17 = stq_9_bits_uop_iw_state;
      5'b01010:
        casez_tmp_17 = stq_10_bits_uop_iw_state;
      5'b01011:
        casez_tmp_17 = stq_11_bits_uop_iw_state;
      5'b01100:
        casez_tmp_17 = stq_12_bits_uop_iw_state;
      5'b01101:
        casez_tmp_17 = stq_13_bits_uop_iw_state;
      5'b01110:
        casez_tmp_17 = stq_14_bits_uop_iw_state;
      5'b01111:
        casez_tmp_17 = stq_15_bits_uop_iw_state;
      5'b10000:
        casez_tmp_17 = stq_16_bits_uop_iw_state;
      5'b10001:
        casez_tmp_17 = stq_17_bits_uop_iw_state;
      5'b10010:
        casez_tmp_17 = stq_18_bits_uop_iw_state;
      5'b10011:
        casez_tmp_17 = stq_19_bits_uop_iw_state;
      5'b10100:
        casez_tmp_17 = stq_20_bits_uop_iw_state;
      5'b10101:
        casez_tmp_17 = stq_21_bits_uop_iw_state;
      5'b10110:
        casez_tmp_17 = stq_22_bits_uop_iw_state;
      5'b10111:
        casez_tmp_17 = stq_23_bits_uop_iw_state;
      5'b11000:
        casez_tmp_17 = stq_24_bits_uop_iw_state;
      5'b11001:
        casez_tmp_17 = stq_25_bits_uop_iw_state;
      5'b11010:
        casez_tmp_17 = stq_26_bits_uop_iw_state;
      5'b11011:
        casez_tmp_17 = stq_27_bits_uop_iw_state;
      5'b11100:
        casez_tmp_17 = stq_28_bits_uop_iw_state;
      5'b11101:
        casez_tmp_17 = stq_29_bits_uop_iw_state;
      5'b11110:
        casez_tmp_17 = stq_30_bits_uop_iw_state;
      default:
        casez_tmp_17 = stq_31_bits_uop_iw_state;
    endcase
  end // always @(*)
  reg         casez_tmp_18;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_18 = stq_0_bits_uop_iw_p1_poisoned;
      5'b00001:
        casez_tmp_18 = stq_1_bits_uop_iw_p1_poisoned;
      5'b00010:
        casez_tmp_18 = stq_2_bits_uop_iw_p1_poisoned;
      5'b00011:
        casez_tmp_18 = stq_3_bits_uop_iw_p1_poisoned;
      5'b00100:
        casez_tmp_18 = stq_4_bits_uop_iw_p1_poisoned;
      5'b00101:
        casez_tmp_18 = stq_5_bits_uop_iw_p1_poisoned;
      5'b00110:
        casez_tmp_18 = stq_6_bits_uop_iw_p1_poisoned;
      5'b00111:
        casez_tmp_18 = stq_7_bits_uop_iw_p1_poisoned;
      5'b01000:
        casez_tmp_18 = stq_8_bits_uop_iw_p1_poisoned;
      5'b01001:
        casez_tmp_18 = stq_9_bits_uop_iw_p1_poisoned;
      5'b01010:
        casez_tmp_18 = stq_10_bits_uop_iw_p1_poisoned;
      5'b01011:
        casez_tmp_18 = stq_11_bits_uop_iw_p1_poisoned;
      5'b01100:
        casez_tmp_18 = stq_12_bits_uop_iw_p1_poisoned;
      5'b01101:
        casez_tmp_18 = stq_13_bits_uop_iw_p1_poisoned;
      5'b01110:
        casez_tmp_18 = stq_14_bits_uop_iw_p1_poisoned;
      5'b01111:
        casez_tmp_18 = stq_15_bits_uop_iw_p1_poisoned;
      5'b10000:
        casez_tmp_18 = stq_16_bits_uop_iw_p1_poisoned;
      5'b10001:
        casez_tmp_18 = stq_17_bits_uop_iw_p1_poisoned;
      5'b10010:
        casez_tmp_18 = stq_18_bits_uop_iw_p1_poisoned;
      5'b10011:
        casez_tmp_18 = stq_19_bits_uop_iw_p1_poisoned;
      5'b10100:
        casez_tmp_18 = stq_20_bits_uop_iw_p1_poisoned;
      5'b10101:
        casez_tmp_18 = stq_21_bits_uop_iw_p1_poisoned;
      5'b10110:
        casez_tmp_18 = stq_22_bits_uop_iw_p1_poisoned;
      5'b10111:
        casez_tmp_18 = stq_23_bits_uop_iw_p1_poisoned;
      5'b11000:
        casez_tmp_18 = stq_24_bits_uop_iw_p1_poisoned;
      5'b11001:
        casez_tmp_18 = stq_25_bits_uop_iw_p1_poisoned;
      5'b11010:
        casez_tmp_18 = stq_26_bits_uop_iw_p1_poisoned;
      5'b11011:
        casez_tmp_18 = stq_27_bits_uop_iw_p1_poisoned;
      5'b11100:
        casez_tmp_18 = stq_28_bits_uop_iw_p1_poisoned;
      5'b11101:
        casez_tmp_18 = stq_29_bits_uop_iw_p1_poisoned;
      5'b11110:
        casez_tmp_18 = stq_30_bits_uop_iw_p1_poisoned;
      default:
        casez_tmp_18 = stq_31_bits_uop_iw_p1_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_19;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_19 = stq_0_bits_uop_iw_p2_poisoned;
      5'b00001:
        casez_tmp_19 = stq_1_bits_uop_iw_p2_poisoned;
      5'b00010:
        casez_tmp_19 = stq_2_bits_uop_iw_p2_poisoned;
      5'b00011:
        casez_tmp_19 = stq_3_bits_uop_iw_p2_poisoned;
      5'b00100:
        casez_tmp_19 = stq_4_bits_uop_iw_p2_poisoned;
      5'b00101:
        casez_tmp_19 = stq_5_bits_uop_iw_p2_poisoned;
      5'b00110:
        casez_tmp_19 = stq_6_bits_uop_iw_p2_poisoned;
      5'b00111:
        casez_tmp_19 = stq_7_bits_uop_iw_p2_poisoned;
      5'b01000:
        casez_tmp_19 = stq_8_bits_uop_iw_p2_poisoned;
      5'b01001:
        casez_tmp_19 = stq_9_bits_uop_iw_p2_poisoned;
      5'b01010:
        casez_tmp_19 = stq_10_bits_uop_iw_p2_poisoned;
      5'b01011:
        casez_tmp_19 = stq_11_bits_uop_iw_p2_poisoned;
      5'b01100:
        casez_tmp_19 = stq_12_bits_uop_iw_p2_poisoned;
      5'b01101:
        casez_tmp_19 = stq_13_bits_uop_iw_p2_poisoned;
      5'b01110:
        casez_tmp_19 = stq_14_bits_uop_iw_p2_poisoned;
      5'b01111:
        casez_tmp_19 = stq_15_bits_uop_iw_p2_poisoned;
      5'b10000:
        casez_tmp_19 = stq_16_bits_uop_iw_p2_poisoned;
      5'b10001:
        casez_tmp_19 = stq_17_bits_uop_iw_p2_poisoned;
      5'b10010:
        casez_tmp_19 = stq_18_bits_uop_iw_p2_poisoned;
      5'b10011:
        casez_tmp_19 = stq_19_bits_uop_iw_p2_poisoned;
      5'b10100:
        casez_tmp_19 = stq_20_bits_uop_iw_p2_poisoned;
      5'b10101:
        casez_tmp_19 = stq_21_bits_uop_iw_p2_poisoned;
      5'b10110:
        casez_tmp_19 = stq_22_bits_uop_iw_p2_poisoned;
      5'b10111:
        casez_tmp_19 = stq_23_bits_uop_iw_p2_poisoned;
      5'b11000:
        casez_tmp_19 = stq_24_bits_uop_iw_p2_poisoned;
      5'b11001:
        casez_tmp_19 = stq_25_bits_uop_iw_p2_poisoned;
      5'b11010:
        casez_tmp_19 = stq_26_bits_uop_iw_p2_poisoned;
      5'b11011:
        casez_tmp_19 = stq_27_bits_uop_iw_p2_poisoned;
      5'b11100:
        casez_tmp_19 = stq_28_bits_uop_iw_p2_poisoned;
      5'b11101:
        casez_tmp_19 = stq_29_bits_uop_iw_p2_poisoned;
      5'b11110:
        casez_tmp_19 = stq_30_bits_uop_iw_p2_poisoned;
      default:
        casez_tmp_19 = stq_31_bits_uop_iw_p2_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_20;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_20 = stq_0_bits_uop_is_br;
      5'b00001:
        casez_tmp_20 = stq_1_bits_uop_is_br;
      5'b00010:
        casez_tmp_20 = stq_2_bits_uop_is_br;
      5'b00011:
        casez_tmp_20 = stq_3_bits_uop_is_br;
      5'b00100:
        casez_tmp_20 = stq_4_bits_uop_is_br;
      5'b00101:
        casez_tmp_20 = stq_5_bits_uop_is_br;
      5'b00110:
        casez_tmp_20 = stq_6_bits_uop_is_br;
      5'b00111:
        casez_tmp_20 = stq_7_bits_uop_is_br;
      5'b01000:
        casez_tmp_20 = stq_8_bits_uop_is_br;
      5'b01001:
        casez_tmp_20 = stq_9_bits_uop_is_br;
      5'b01010:
        casez_tmp_20 = stq_10_bits_uop_is_br;
      5'b01011:
        casez_tmp_20 = stq_11_bits_uop_is_br;
      5'b01100:
        casez_tmp_20 = stq_12_bits_uop_is_br;
      5'b01101:
        casez_tmp_20 = stq_13_bits_uop_is_br;
      5'b01110:
        casez_tmp_20 = stq_14_bits_uop_is_br;
      5'b01111:
        casez_tmp_20 = stq_15_bits_uop_is_br;
      5'b10000:
        casez_tmp_20 = stq_16_bits_uop_is_br;
      5'b10001:
        casez_tmp_20 = stq_17_bits_uop_is_br;
      5'b10010:
        casez_tmp_20 = stq_18_bits_uop_is_br;
      5'b10011:
        casez_tmp_20 = stq_19_bits_uop_is_br;
      5'b10100:
        casez_tmp_20 = stq_20_bits_uop_is_br;
      5'b10101:
        casez_tmp_20 = stq_21_bits_uop_is_br;
      5'b10110:
        casez_tmp_20 = stq_22_bits_uop_is_br;
      5'b10111:
        casez_tmp_20 = stq_23_bits_uop_is_br;
      5'b11000:
        casez_tmp_20 = stq_24_bits_uop_is_br;
      5'b11001:
        casez_tmp_20 = stq_25_bits_uop_is_br;
      5'b11010:
        casez_tmp_20 = stq_26_bits_uop_is_br;
      5'b11011:
        casez_tmp_20 = stq_27_bits_uop_is_br;
      5'b11100:
        casez_tmp_20 = stq_28_bits_uop_is_br;
      5'b11101:
        casez_tmp_20 = stq_29_bits_uop_is_br;
      5'b11110:
        casez_tmp_20 = stq_30_bits_uop_is_br;
      default:
        casez_tmp_20 = stq_31_bits_uop_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_21;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_21 = stq_0_bits_uop_is_jalr;
      5'b00001:
        casez_tmp_21 = stq_1_bits_uop_is_jalr;
      5'b00010:
        casez_tmp_21 = stq_2_bits_uop_is_jalr;
      5'b00011:
        casez_tmp_21 = stq_3_bits_uop_is_jalr;
      5'b00100:
        casez_tmp_21 = stq_4_bits_uop_is_jalr;
      5'b00101:
        casez_tmp_21 = stq_5_bits_uop_is_jalr;
      5'b00110:
        casez_tmp_21 = stq_6_bits_uop_is_jalr;
      5'b00111:
        casez_tmp_21 = stq_7_bits_uop_is_jalr;
      5'b01000:
        casez_tmp_21 = stq_8_bits_uop_is_jalr;
      5'b01001:
        casez_tmp_21 = stq_9_bits_uop_is_jalr;
      5'b01010:
        casez_tmp_21 = stq_10_bits_uop_is_jalr;
      5'b01011:
        casez_tmp_21 = stq_11_bits_uop_is_jalr;
      5'b01100:
        casez_tmp_21 = stq_12_bits_uop_is_jalr;
      5'b01101:
        casez_tmp_21 = stq_13_bits_uop_is_jalr;
      5'b01110:
        casez_tmp_21 = stq_14_bits_uop_is_jalr;
      5'b01111:
        casez_tmp_21 = stq_15_bits_uop_is_jalr;
      5'b10000:
        casez_tmp_21 = stq_16_bits_uop_is_jalr;
      5'b10001:
        casez_tmp_21 = stq_17_bits_uop_is_jalr;
      5'b10010:
        casez_tmp_21 = stq_18_bits_uop_is_jalr;
      5'b10011:
        casez_tmp_21 = stq_19_bits_uop_is_jalr;
      5'b10100:
        casez_tmp_21 = stq_20_bits_uop_is_jalr;
      5'b10101:
        casez_tmp_21 = stq_21_bits_uop_is_jalr;
      5'b10110:
        casez_tmp_21 = stq_22_bits_uop_is_jalr;
      5'b10111:
        casez_tmp_21 = stq_23_bits_uop_is_jalr;
      5'b11000:
        casez_tmp_21 = stq_24_bits_uop_is_jalr;
      5'b11001:
        casez_tmp_21 = stq_25_bits_uop_is_jalr;
      5'b11010:
        casez_tmp_21 = stq_26_bits_uop_is_jalr;
      5'b11011:
        casez_tmp_21 = stq_27_bits_uop_is_jalr;
      5'b11100:
        casez_tmp_21 = stq_28_bits_uop_is_jalr;
      5'b11101:
        casez_tmp_21 = stq_29_bits_uop_is_jalr;
      5'b11110:
        casez_tmp_21 = stq_30_bits_uop_is_jalr;
      default:
        casez_tmp_21 = stq_31_bits_uop_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_22;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_22 = stq_0_bits_uop_is_jal;
      5'b00001:
        casez_tmp_22 = stq_1_bits_uop_is_jal;
      5'b00010:
        casez_tmp_22 = stq_2_bits_uop_is_jal;
      5'b00011:
        casez_tmp_22 = stq_3_bits_uop_is_jal;
      5'b00100:
        casez_tmp_22 = stq_4_bits_uop_is_jal;
      5'b00101:
        casez_tmp_22 = stq_5_bits_uop_is_jal;
      5'b00110:
        casez_tmp_22 = stq_6_bits_uop_is_jal;
      5'b00111:
        casez_tmp_22 = stq_7_bits_uop_is_jal;
      5'b01000:
        casez_tmp_22 = stq_8_bits_uop_is_jal;
      5'b01001:
        casez_tmp_22 = stq_9_bits_uop_is_jal;
      5'b01010:
        casez_tmp_22 = stq_10_bits_uop_is_jal;
      5'b01011:
        casez_tmp_22 = stq_11_bits_uop_is_jal;
      5'b01100:
        casez_tmp_22 = stq_12_bits_uop_is_jal;
      5'b01101:
        casez_tmp_22 = stq_13_bits_uop_is_jal;
      5'b01110:
        casez_tmp_22 = stq_14_bits_uop_is_jal;
      5'b01111:
        casez_tmp_22 = stq_15_bits_uop_is_jal;
      5'b10000:
        casez_tmp_22 = stq_16_bits_uop_is_jal;
      5'b10001:
        casez_tmp_22 = stq_17_bits_uop_is_jal;
      5'b10010:
        casez_tmp_22 = stq_18_bits_uop_is_jal;
      5'b10011:
        casez_tmp_22 = stq_19_bits_uop_is_jal;
      5'b10100:
        casez_tmp_22 = stq_20_bits_uop_is_jal;
      5'b10101:
        casez_tmp_22 = stq_21_bits_uop_is_jal;
      5'b10110:
        casez_tmp_22 = stq_22_bits_uop_is_jal;
      5'b10111:
        casez_tmp_22 = stq_23_bits_uop_is_jal;
      5'b11000:
        casez_tmp_22 = stq_24_bits_uop_is_jal;
      5'b11001:
        casez_tmp_22 = stq_25_bits_uop_is_jal;
      5'b11010:
        casez_tmp_22 = stq_26_bits_uop_is_jal;
      5'b11011:
        casez_tmp_22 = stq_27_bits_uop_is_jal;
      5'b11100:
        casez_tmp_22 = stq_28_bits_uop_is_jal;
      5'b11101:
        casez_tmp_22 = stq_29_bits_uop_is_jal;
      5'b11110:
        casez_tmp_22 = stq_30_bits_uop_is_jal;
      default:
        casez_tmp_22 = stq_31_bits_uop_is_jal;
    endcase
  end // always @(*)
  reg         casez_tmp_23;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_23 = stq_0_bits_uop_is_sfb;
      5'b00001:
        casez_tmp_23 = stq_1_bits_uop_is_sfb;
      5'b00010:
        casez_tmp_23 = stq_2_bits_uop_is_sfb;
      5'b00011:
        casez_tmp_23 = stq_3_bits_uop_is_sfb;
      5'b00100:
        casez_tmp_23 = stq_4_bits_uop_is_sfb;
      5'b00101:
        casez_tmp_23 = stq_5_bits_uop_is_sfb;
      5'b00110:
        casez_tmp_23 = stq_6_bits_uop_is_sfb;
      5'b00111:
        casez_tmp_23 = stq_7_bits_uop_is_sfb;
      5'b01000:
        casez_tmp_23 = stq_8_bits_uop_is_sfb;
      5'b01001:
        casez_tmp_23 = stq_9_bits_uop_is_sfb;
      5'b01010:
        casez_tmp_23 = stq_10_bits_uop_is_sfb;
      5'b01011:
        casez_tmp_23 = stq_11_bits_uop_is_sfb;
      5'b01100:
        casez_tmp_23 = stq_12_bits_uop_is_sfb;
      5'b01101:
        casez_tmp_23 = stq_13_bits_uop_is_sfb;
      5'b01110:
        casez_tmp_23 = stq_14_bits_uop_is_sfb;
      5'b01111:
        casez_tmp_23 = stq_15_bits_uop_is_sfb;
      5'b10000:
        casez_tmp_23 = stq_16_bits_uop_is_sfb;
      5'b10001:
        casez_tmp_23 = stq_17_bits_uop_is_sfb;
      5'b10010:
        casez_tmp_23 = stq_18_bits_uop_is_sfb;
      5'b10011:
        casez_tmp_23 = stq_19_bits_uop_is_sfb;
      5'b10100:
        casez_tmp_23 = stq_20_bits_uop_is_sfb;
      5'b10101:
        casez_tmp_23 = stq_21_bits_uop_is_sfb;
      5'b10110:
        casez_tmp_23 = stq_22_bits_uop_is_sfb;
      5'b10111:
        casez_tmp_23 = stq_23_bits_uop_is_sfb;
      5'b11000:
        casez_tmp_23 = stq_24_bits_uop_is_sfb;
      5'b11001:
        casez_tmp_23 = stq_25_bits_uop_is_sfb;
      5'b11010:
        casez_tmp_23 = stq_26_bits_uop_is_sfb;
      5'b11011:
        casez_tmp_23 = stq_27_bits_uop_is_sfb;
      5'b11100:
        casez_tmp_23 = stq_28_bits_uop_is_sfb;
      5'b11101:
        casez_tmp_23 = stq_29_bits_uop_is_sfb;
      5'b11110:
        casez_tmp_23 = stq_30_bits_uop_is_sfb;
      default:
        casez_tmp_23 = stq_31_bits_uop_is_sfb;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_24;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_24 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_24 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_24 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_24 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_24 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_24 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_24 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_24 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_24 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_24 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_24 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_24 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_24 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_24 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_24 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_24 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_24 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_24 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_24 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_24 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_24 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_24 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_24 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_24 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_24 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_24 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_24 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_24 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_24 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_24 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_24 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_24 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_25;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_25 = stq_0_bits_uop_br_tag;
      5'b00001:
        casez_tmp_25 = stq_1_bits_uop_br_tag;
      5'b00010:
        casez_tmp_25 = stq_2_bits_uop_br_tag;
      5'b00011:
        casez_tmp_25 = stq_3_bits_uop_br_tag;
      5'b00100:
        casez_tmp_25 = stq_4_bits_uop_br_tag;
      5'b00101:
        casez_tmp_25 = stq_5_bits_uop_br_tag;
      5'b00110:
        casez_tmp_25 = stq_6_bits_uop_br_tag;
      5'b00111:
        casez_tmp_25 = stq_7_bits_uop_br_tag;
      5'b01000:
        casez_tmp_25 = stq_8_bits_uop_br_tag;
      5'b01001:
        casez_tmp_25 = stq_9_bits_uop_br_tag;
      5'b01010:
        casez_tmp_25 = stq_10_bits_uop_br_tag;
      5'b01011:
        casez_tmp_25 = stq_11_bits_uop_br_tag;
      5'b01100:
        casez_tmp_25 = stq_12_bits_uop_br_tag;
      5'b01101:
        casez_tmp_25 = stq_13_bits_uop_br_tag;
      5'b01110:
        casez_tmp_25 = stq_14_bits_uop_br_tag;
      5'b01111:
        casez_tmp_25 = stq_15_bits_uop_br_tag;
      5'b10000:
        casez_tmp_25 = stq_16_bits_uop_br_tag;
      5'b10001:
        casez_tmp_25 = stq_17_bits_uop_br_tag;
      5'b10010:
        casez_tmp_25 = stq_18_bits_uop_br_tag;
      5'b10011:
        casez_tmp_25 = stq_19_bits_uop_br_tag;
      5'b10100:
        casez_tmp_25 = stq_20_bits_uop_br_tag;
      5'b10101:
        casez_tmp_25 = stq_21_bits_uop_br_tag;
      5'b10110:
        casez_tmp_25 = stq_22_bits_uop_br_tag;
      5'b10111:
        casez_tmp_25 = stq_23_bits_uop_br_tag;
      5'b11000:
        casez_tmp_25 = stq_24_bits_uop_br_tag;
      5'b11001:
        casez_tmp_25 = stq_25_bits_uop_br_tag;
      5'b11010:
        casez_tmp_25 = stq_26_bits_uop_br_tag;
      5'b11011:
        casez_tmp_25 = stq_27_bits_uop_br_tag;
      5'b11100:
        casez_tmp_25 = stq_28_bits_uop_br_tag;
      5'b11101:
        casez_tmp_25 = stq_29_bits_uop_br_tag;
      5'b11110:
        casez_tmp_25 = stq_30_bits_uop_br_tag;
      default:
        casez_tmp_25 = stq_31_bits_uop_br_tag;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_26;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_26 = stq_0_bits_uop_ftq_idx;
      5'b00001:
        casez_tmp_26 = stq_1_bits_uop_ftq_idx;
      5'b00010:
        casez_tmp_26 = stq_2_bits_uop_ftq_idx;
      5'b00011:
        casez_tmp_26 = stq_3_bits_uop_ftq_idx;
      5'b00100:
        casez_tmp_26 = stq_4_bits_uop_ftq_idx;
      5'b00101:
        casez_tmp_26 = stq_5_bits_uop_ftq_idx;
      5'b00110:
        casez_tmp_26 = stq_6_bits_uop_ftq_idx;
      5'b00111:
        casez_tmp_26 = stq_7_bits_uop_ftq_idx;
      5'b01000:
        casez_tmp_26 = stq_8_bits_uop_ftq_idx;
      5'b01001:
        casez_tmp_26 = stq_9_bits_uop_ftq_idx;
      5'b01010:
        casez_tmp_26 = stq_10_bits_uop_ftq_idx;
      5'b01011:
        casez_tmp_26 = stq_11_bits_uop_ftq_idx;
      5'b01100:
        casez_tmp_26 = stq_12_bits_uop_ftq_idx;
      5'b01101:
        casez_tmp_26 = stq_13_bits_uop_ftq_idx;
      5'b01110:
        casez_tmp_26 = stq_14_bits_uop_ftq_idx;
      5'b01111:
        casez_tmp_26 = stq_15_bits_uop_ftq_idx;
      5'b10000:
        casez_tmp_26 = stq_16_bits_uop_ftq_idx;
      5'b10001:
        casez_tmp_26 = stq_17_bits_uop_ftq_idx;
      5'b10010:
        casez_tmp_26 = stq_18_bits_uop_ftq_idx;
      5'b10011:
        casez_tmp_26 = stq_19_bits_uop_ftq_idx;
      5'b10100:
        casez_tmp_26 = stq_20_bits_uop_ftq_idx;
      5'b10101:
        casez_tmp_26 = stq_21_bits_uop_ftq_idx;
      5'b10110:
        casez_tmp_26 = stq_22_bits_uop_ftq_idx;
      5'b10111:
        casez_tmp_26 = stq_23_bits_uop_ftq_idx;
      5'b11000:
        casez_tmp_26 = stq_24_bits_uop_ftq_idx;
      5'b11001:
        casez_tmp_26 = stq_25_bits_uop_ftq_idx;
      5'b11010:
        casez_tmp_26 = stq_26_bits_uop_ftq_idx;
      5'b11011:
        casez_tmp_26 = stq_27_bits_uop_ftq_idx;
      5'b11100:
        casez_tmp_26 = stq_28_bits_uop_ftq_idx;
      5'b11101:
        casez_tmp_26 = stq_29_bits_uop_ftq_idx;
      5'b11110:
        casez_tmp_26 = stq_30_bits_uop_ftq_idx;
      default:
        casez_tmp_26 = stq_31_bits_uop_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_27;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_27 = stq_0_bits_uop_edge_inst;
      5'b00001:
        casez_tmp_27 = stq_1_bits_uop_edge_inst;
      5'b00010:
        casez_tmp_27 = stq_2_bits_uop_edge_inst;
      5'b00011:
        casez_tmp_27 = stq_3_bits_uop_edge_inst;
      5'b00100:
        casez_tmp_27 = stq_4_bits_uop_edge_inst;
      5'b00101:
        casez_tmp_27 = stq_5_bits_uop_edge_inst;
      5'b00110:
        casez_tmp_27 = stq_6_bits_uop_edge_inst;
      5'b00111:
        casez_tmp_27 = stq_7_bits_uop_edge_inst;
      5'b01000:
        casez_tmp_27 = stq_8_bits_uop_edge_inst;
      5'b01001:
        casez_tmp_27 = stq_9_bits_uop_edge_inst;
      5'b01010:
        casez_tmp_27 = stq_10_bits_uop_edge_inst;
      5'b01011:
        casez_tmp_27 = stq_11_bits_uop_edge_inst;
      5'b01100:
        casez_tmp_27 = stq_12_bits_uop_edge_inst;
      5'b01101:
        casez_tmp_27 = stq_13_bits_uop_edge_inst;
      5'b01110:
        casez_tmp_27 = stq_14_bits_uop_edge_inst;
      5'b01111:
        casez_tmp_27 = stq_15_bits_uop_edge_inst;
      5'b10000:
        casez_tmp_27 = stq_16_bits_uop_edge_inst;
      5'b10001:
        casez_tmp_27 = stq_17_bits_uop_edge_inst;
      5'b10010:
        casez_tmp_27 = stq_18_bits_uop_edge_inst;
      5'b10011:
        casez_tmp_27 = stq_19_bits_uop_edge_inst;
      5'b10100:
        casez_tmp_27 = stq_20_bits_uop_edge_inst;
      5'b10101:
        casez_tmp_27 = stq_21_bits_uop_edge_inst;
      5'b10110:
        casez_tmp_27 = stq_22_bits_uop_edge_inst;
      5'b10111:
        casez_tmp_27 = stq_23_bits_uop_edge_inst;
      5'b11000:
        casez_tmp_27 = stq_24_bits_uop_edge_inst;
      5'b11001:
        casez_tmp_27 = stq_25_bits_uop_edge_inst;
      5'b11010:
        casez_tmp_27 = stq_26_bits_uop_edge_inst;
      5'b11011:
        casez_tmp_27 = stq_27_bits_uop_edge_inst;
      5'b11100:
        casez_tmp_27 = stq_28_bits_uop_edge_inst;
      5'b11101:
        casez_tmp_27 = stq_29_bits_uop_edge_inst;
      5'b11110:
        casez_tmp_27 = stq_30_bits_uop_edge_inst;
      default:
        casez_tmp_27 = stq_31_bits_uop_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_28;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_28 = stq_0_bits_uop_pc_lob;
      5'b00001:
        casez_tmp_28 = stq_1_bits_uop_pc_lob;
      5'b00010:
        casez_tmp_28 = stq_2_bits_uop_pc_lob;
      5'b00011:
        casez_tmp_28 = stq_3_bits_uop_pc_lob;
      5'b00100:
        casez_tmp_28 = stq_4_bits_uop_pc_lob;
      5'b00101:
        casez_tmp_28 = stq_5_bits_uop_pc_lob;
      5'b00110:
        casez_tmp_28 = stq_6_bits_uop_pc_lob;
      5'b00111:
        casez_tmp_28 = stq_7_bits_uop_pc_lob;
      5'b01000:
        casez_tmp_28 = stq_8_bits_uop_pc_lob;
      5'b01001:
        casez_tmp_28 = stq_9_bits_uop_pc_lob;
      5'b01010:
        casez_tmp_28 = stq_10_bits_uop_pc_lob;
      5'b01011:
        casez_tmp_28 = stq_11_bits_uop_pc_lob;
      5'b01100:
        casez_tmp_28 = stq_12_bits_uop_pc_lob;
      5'b01101:
        casez_tmp_28 = stq_13_bits_uop_pc_lob;
      5'b01110:
        casez_tmp_28 = stq_14_bits_uop_pc_lob;
      5'b01111:
        casez_tmp_28 = stq_15_bits_uop_pc_lob;
      5'b10000:
        casez_tmp_28 = stq_16_bits_uop_pc_lob;
      5'b10001:
        casez_tmp_28 = stq_17_bits_uop_pc_lob;
      5'b10010:
        casez_tmp_28 = stq_18_bits_uop_pc_lob;
      5'b10011:
        casez_tmp_28 = stq_19_bits_uop_pc_lob;
      5'b10100:
        casez_tmp_28 = stq_20_bits_uop_pc_lob;
      5'b10101:
        casez_tmp_28 = stq_21_bits_uop_pc_lob;
      5'b10110:
        casez_tmp_28 = stq_22_bits_uop_pc_lob;
      5'b10111:
        casez_tmp_28 = stq_23_bits_uop_pc_lob;
      5'b11000:
        casez_tmp_28 = stq_24_bits_uop_pc_lob;
      5'b11001:
        casez_tmp_28 = stq_25_bits_uop_pc_lob;
      5'b11010:
        casez_tmp_28 = stq_26_bits_uop_pc_lob;
      5'b11011:
        casez_tmp_28 = stq_27_bits_uop_pc_lob;
      5'b11100:
        casez_tmp_28 = stq_28_bits_uop_pc_lob;
      5'b11101:
        casez_tmp_28 = stq_29_bits_uop_pc_lob;
      5'b11110:
        casez_tmp_28 = stq_30_bits_uop_pc_lob;
      default:
        casez_tmp_28 = stq_31_bits_uop_pc_lob;
    endcase
  end // always @(*)
  reg         casez_tmp_29;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_29 = stq_0_bits_uop_taken;
      5'b00001:
        casez_tmp_29 = stq_1_bits_uop_taken;
      5'b00010:
        casez_tmp_29 = stq_2_bits_uop_taken;
      5'b00011:
        casez_tmp_29 = stq_3_bits_uop_taken;
      5'b00100:
        casez_tmp_29 = stq_4_bits_uop_taken;
      5'b00101:
        casez_tmp_29 = stq_5_bits_uop_taken;
      5'b00110:
        casez_tmp_29 = stq_6_bits_uop_taken;
      5'b00111:
        casez_tmp_29 = stq_7_bits_uop_taken;
      5'b01000:
        casez_tmp_29 = stq_8_bits_uop_taken;
      5'b01001:
        casez_tmp_29 = stq_9_bits_uop_taken;
      5'b01010:
        casez_tmp_29 = stq_10_bits_uop_taken;
      5'b01011:
        casez_tmp_29 = stq_11_bits_uop_taken;
      5'b01100:
        casez_tmp_29 = stq_12_bits_uop_taken;
      5'b01101:
        casez_tmp_29 = stq_13_bits_uop_taken;
      5'b01110:
        casez_tmp_29 = stq_14_bits_uop_taken;
      5'b01111:
        casez_tmp_29 = stq_15_bits_uop_taken;
      5'b10000:
        casez_tmp_29 = stq_16_bits_uop_taken;
      5'b10001:
        casez_tmp_29 = stq_17_bits_uop_taken;
      5'b10010:
        casez_tmp_29 = stq_18_bits_uop_taken;
      5'b10011:
        casez_tmp_29 = stq_19_bits_uop_taken;
      5'b10100:
        casez_tmp_29 = stq_20_bits_uop_taken;
      5'b10101:
        casez_tmp_29 = stq_21_bits_uop_taken;
      5'b10110:
        casez_tmp_29 = stq_22_bits_uop_taken;
      5'b10111:
        casez_tmp_29 = stq_23_bits_uop_taken;
      5'b11000:
        casez_tmp_29 = stq_24_bits_uop_taken;
      5'b11001:
        casez_tmp_29 = stq_25_bits_uop_taken;
      5'b11010:
        casez_tmp_29 = stq_26_bits_uop_taken;
      5'b11011:
        casez_tmp_29 = stq_27_bits_uop_taken;
      5'b11100:
        casez_tmp_29 = stq_28_bits_uop_taken;
      5'b11101:
        casez_tmp_29 = stq_29_bits_uop_taken;
      5'b11110:
        casez_tmp_29 = stq_30_bits_uop_taken;
      default:
        casez_tmp_29 = stq_31_bits_uop_taken;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_30;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_30 = stq_0_bits_uop_imm_packed;
      5'b00001:
        casez_tmp_30 = stq_1_bits_uop_imm_packed;
      5'b00010:
        casez_tmp_30 = stq_2_bits_uop_imm_packed;
      5'b00011:
        casez_tmp_30 = stq_3_bits_uop_imm_packed;
      5'b00100:
        casez_tmp_30 = stq_4_bits_uop_imm_packed;
      5'b00101:
        casez_tmp_30 = stq_5_bits_uop_imm_packed;
      5'b00110:
        casez_tmp_30 = stq_6_bits_uop_imm_packed;
      5'b00111:
        casez_tmp_30 = stq_7_bits_uop_imm_packed;
      5'b01000:
        casez_tmp_30 = stq_8_bits_uop_imm_packed;
      5'b01001:
        casez_tmp_30 = stq_9_bits_uop_imm_packed;
      5'b01010:
        casez_tmp_30 = stq_10_bits_uop_imm_packed;
      5'b01011:
        casez_tmp_30 = stq_11_bits_uop_imm_packed;
      5'b01100:
        casez_tmp_30 = stq_12_bits_uop_imm_packed;
      5'b01101:
        casez_tmp_30 = stq_13_bits_uop_imm_packed;
      5'b01110:
        casez_tmp_30 = stq_14_bits_uop_imm_packed;
      5'b01111:
        casez_tmp_30 = stq_15_bits_uop_imm_packed;
      5'b10000:
        casez_tmp_30 = stq_16_bits_uop_imm_packed;
      5'b10001:
        casez_tmp_30 = stq_17_bits_uop_imm_packed;
      5'b10010:
        casez_tmp_30 = stq_18_bits_uop_imm_packed;
      5'b10011:
        casez_tmp_30 = stq_19_bits_uop_imm_packed;
      5'b10100:
        casez_tmp_30 = stq_20_bits_uop_imm_packed;
      5'b10101:
        casez_tmp_30 = stq_21_bits_uop_imm_packed;
      5'b10110:
        casez_tmp_30 = stq_22_bits_uop_imm_packed;
      5'b10111:
        casez_tmp_30 = stq_23_bits_uop_imm_packed;
      5'b11000:
        casez_tmp_30 = stq_24_bits_uop_imm_packed;
      5'b11001:
        casez_tmp_30 = stq_25_bits_uop_imm_packed;
      5'b11010:
        casez_tmp_30 = stq_26_bits_uop_imm_packed;
      5'b11011:
        casez_tmp_30 = stq_27_bits_uop_imm_packed;
      5'b11100:
        casez_tmp_30 = stq_28_bits_uop_imm_packed;
      5'b11101:
        casez_tmp_30 = stq_29_bits_uop_imm_packed;
      5'b11110:
        casez_tmp_30 = stq_30_bits_uop_imm_packed;
      default:
        casez_tmp_30 = stq_31_bits_uop_imm_packed;
    endcase
  end // always @(*)
  reg  [11:0] casez_tmp_31;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_31 = stq_0_bits_uop_csr_addr;
      5'b00001:
        casez_tmp_31 = stq_1_bits_uop_csr_addr;
      5'b00010:
        casez_tmp_31 = stq_2_bits_uop_csr_addr;
      5'b00011:
        casez_tmp_31 = stq_3_bits_uop_csr_addr;
      5'b00100:
        casez_tmp_31 = stq_4_bits_uop_csr_addr;
      5'b00101:
        casez_tmp_31 = stq_5_bits_uop_csr_addr;
      5'b00110:
        casez_tmp_31 = stq_6_bits_uop_csr_addr;
      5'b00111:
        casez_tmp_31 = stq_7_bits_uop_csr_addr;
      5'b01000:
        casez_tmp_31 = stq_8_bits_uop_csr_addr;
      5'b01001:
        casez_tmp_31 = stq_9_bits_uop_csr_addr;
      5'b01010:
        casez_tmp_31 = stq_10_bits_uop_csr_addr;
      5'b01011:
        casez_tmp_31 = stq_11_bits_uop_csr_addr;
      5'b01100:
        casez_tmp_31 = stq_12_bits_uop_csr_addr;
      5'b01101:
        casez_tmp_31 = stq_13_bits_uop_csr_addr;
      5'b01110:
        casez_tmp_31 = stq_14_bits_uop_csr_addr;
      5'b01111:
        casez_tmp_31 = stq_15_bits_uop_csr_addr;
      5'b10000:
        casez_tmp_31 = stq_16_bits_uop_csr_addr;
      5'b10001:
        casez_tmp_31 = stq_17_bits_uop_csr_addr;
      5'b10010:
        casez_tmp_31 = stq_18_bits_uop_csr_addr;
      5'b10011:
        casez_tmp_31 = stq_19_bits_uop_csr_addr;
      5'b10100:
        casez_tmp_31 = stq_20_bits_uop_csr_addr;
      5'b10101:
        casez_tmp_31 = stq_21_bits_uop_csr_addr;
      5'b10110:
        casez_tmp_31 = stq_22_bits_uop_csr_addr;
      5'b10111:
        casez_tmp_31 = stq_23_bits_uop_csr_addr;
      5'b11000:
        casez_tmp_31 = stq_24_bits_uop_csr_addr;
      5'b11001:
        casez_tmp_31 = stq_25_bits_uop_csr_addr;
      5'b11010:
        casez_tmp_31 = stq_26_bits_uop_csr_addr;
      5'b11011:
        casez_tmp_31 = stq_27_bits_uop_csr_addr;
      5'b11100:
        casez_tmp_31 = stq_28_bits_uop_csr_addr;
      5'b11101:
        casez_tmp_31 = stq_29_bits_uop_csr_addr;
      5'b11110:
        casez_tmp_31 = stq_30_bits_uop_csr_addr;
      default:
        casez_tmp_31 = stq_31_bits_uop_csr_addr;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_32;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_32 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_32 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_32 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_32 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_32 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_32 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_32 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_32 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_32 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_32 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_32 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_32 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_32 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_32 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_32 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_32 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_32 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_32 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_32 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_32 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_32 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_32 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_32 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_32 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_32 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_32 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_32 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_32 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_32 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_32 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_32 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_32 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_33;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_33 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_33 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_33 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_33 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_33 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_33 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_33 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_33 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_33 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_33 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_33 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_33 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_33 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_33 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_33 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_33 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_33 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_33 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_33 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_33 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_33 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_33 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_33 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_33 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_33 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_33 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_33 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_33 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_33 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_33 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_33 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_33 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_34;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_34 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_34 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_34 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_34 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_34 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_34 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_34 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_34 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_34 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_34 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_34 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_34 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_34 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_34 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_34 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_34 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_34 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_34 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_34 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_34 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_34 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_34 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_34 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_34 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_34 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_34 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_34 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_34 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_34 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_34 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_34 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_34 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_35;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_35 = stq_0_bits_uop_rxq_idx;
      5'b00001:
        casez_tmp_35 = stq_1_bits_uop_rxq_idx;
      5'b00010:
        casez_tmp_35 = stq_2_bits_uop_rxq_idx;
      5'b00011:
        casez_tmp_35 = stq_3_bits_uop_rxq_idx;
      5'b00100:
        casez_tmp_35 = stq_4_bits_uop_rxq_idx;
      5'b00101:
        casez_tmp_35 = stq_5_bits_uop_rxq_idx;
      5'b00110:
        casez_tmp_35 = stq_6_bits_uop_rxq_idx;
      5'b00111:
        casez_tmp_35 = stq_7_bits_uop_rxq_idx;
      5'b01000:
        casez_tmp_35 = stq_8_bits_uop_rxq_idx;
      5'b01001:
        casez_tmp_35 = stq_9_bits_uop_rxq_idx;
      5'b01010:
        casez_tmp_35 = stq_10_bits_uop_rxq_idx;
      5'b01011:
        casez_tmp_35 = stq_11_bits_uop_rxq_idx;
      5'b01100:
        casez_tmp_35 = stq_12_bits_uop_rxq_idx;
      5'b01101:
        casez_tmp_35 = stq_13_bits_uop_rxq_idx;
      5'b01110:
        casez_tmp_35 = stq_14_bits_uop_rxq_idx;
      5'b01111:
        casez_tmp_35 = stq_15_bits_uop_rxq_idx;
      5'b10000:
        casez_tmp_35 = stq_16_bits_uop_rxq_idx;
      5'b10001:
        casez_tmp_35 = stq_17_bits_uop_rxq_idx;
      5'b10010:
        casez_tmp_35 = stq_18_bits_uop_rxq_idx;
      5'b10011:
        casez_tmp_35 = stq_19_bits_uop_rxq_idx;
      5'b10100:
        casez_tmp_35 = stq_20_bits_uop_rxq_idx;
      5'b10101:
        casez_tmp_35 = stq_21_bits_uop_rxq_idx;
      5'b10110:
        casez_tmp_35 = stq_22_bits_uop_rxq_idx;
      5'b10111:
        casez_tmp_35 = stq_23_bits_uop_rxq_idx;
      5'b11000:
        casez_tmp_35 = stq_24_bits_uop_rxq_idx;
      5'b11001:
        casez_tmp_35 = stq_25_bits_uop_rxq_idx;
      5'b11010:
        casez_tmp_35 = stq_26_bits_uop_rxq_idx;
      5'b11011:
        casez_tmp_35 = stq_27_bits_uop_rxq_idx;
      5'b11100:
        casez_tmp_35 = stq_28_bits_uop_rxq_idx;
      5'b11101:
        casez_tmp_35 = stq_29_bits_uop_rxq_idx;
      5'b11110:
        casez_tmp_35 = stq_30_bits_uop_rxq_idx;
      default:
        casez_tmp_35 = stq_31_bits_uop_rxq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_36;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_36 = stq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_36 = stq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_36 = stq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_36 = stq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_36 = stq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_36 = stq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_36 = stq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_36 = stq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_36 = stq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_36 = stq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_36 = stq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_36 = stq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_36 = stq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_36 = stq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_36 = stq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_36 = stq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_36 = stq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_36 = stq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_36 = stq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_36 = stq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_36 = stq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_36 = stq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_36 = stq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_36 = stq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_36 = stq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_36 = stq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_36 = stq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_36 = stq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_36 = stq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_36 = stq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_36 = stq_30_bits_uop_pdst;
      default:
        casez_tmp_36 = stq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_37;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_37 = stq_0_bits_uop_prs1;
      5'b00001:
        casez_tmp_37 = stq_1_bits_uop_prs1;
      5'b00010:
        casez_tmp_37 = stq_2_bits_uop_prs1;
      5'b00011:
        casez_tmp_37 = stq_3_bits_uop_prs1;
      5'b00100:
        casez_tmp_37 = stq_4_bits_uop_prs1;
      5'b00101:
        casez_tmp_37 = stq_5_bits_uop_prs1;
      5'b00110:
        casez_tmp_37 = stq_6_bits_uop_prs1;
      5'b00111:
        casez_tmp_37 = stq_7_bits_uop_prs1;
      5'b01000:
        casez_tmp_37 = stq_8_bits_uop_prs1;
      5'b01001:
        casez_tmp_37 = stq_9_bits_uop_prs1;
      5'b01010:
        casez_tmp_37 = stq_10_bits_uop_prs1;
      5'b01011:
        casez_tmp_37 = stq_11_bits_uop_prs1;
      5'b01100:
        casez_tmp_37 = stq_12_bits_uop_prs1;
      5'b01101:
        casez_tmp_37 = stq_13_bits_uop_prs1;
      5'b01110:
        casez_tmp_37 = stq_14_bits_uop_prs1;
      5'b01111:
        casez_tmp_37 = stq_15_bits_uop_prs1;
      5'b10000:
        casez_tmp_37 = stq_16_bits_uop_prs1;
      5'b10001:
        casez_tmp_37 = stq_17_bits_uop_prs1;
      5'b10010:
        casez_tmp_37 = stq_18_bits_uop_prs1;
      5'b10011:
        casez_tmp_37 = stq_19_bits_uop_prs1;
      5'b10100:
        casez_tmp_37 = stq_20_bits_uop_prs1;
      5'b10101:
        casez_tmp_37 = stq_21_bits_uop_prs1;
      5'b10110:
        casez_tmp_37 = stq_22_bits_uop_prs1;
      5'b10111:
        casez_tmp_37 = stq_23_bits_uop_prs1;
      5'b11000:
        casez_tmp_37 = stq_24_bits_uop_prs1;
      5'b11001:
        casez_tmp_37 = stq_25_bits_uop_prs1;
      5'b11010:
        casez_tmp_37 = stq_26_bits_uop_prs1;
      5'b11011:
        casez_tmp_37 = stq_27_bits_uop_prs1;
      5'b11100:
        casez_tmp_37 = stq_28_bits_uop_prs1;
      5'b11101:
        casez_tmp_37 = stq_29_bits_uop_prs1;
      5'b11110:
        casez_tmp_37 = stq_30_bits_uop_prs1;
      default:
        casez_tmp_37 = stq_31_bits_uop_prs1;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_38;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_38 = stq_0_bits_uop_prs2;
      5'b00001:
        casez_tmp_38 = stq_1_bits_uop_prs2;
      5'b00010:
        casez_tmp_38 = stq_2_bits_uop_prs2;
      5'b00011:
        casez_tmp_38 = stq_3_bits_uop_prs2;
      5'b00100:
        casez_tmp_38 = stq_4_bits_uop_prs2;
      5'b00101:
        casez_tmp_38 = stq_5_bits_uop_prs2;
      5'b00110:
        casez_tmp_38 = stq_6_bits_uop_prs2;
      5'b00111:
        casez_tmp_38 = stq_7_bits_uop_prs2;
      5'b01000:
        casez_tmp_38 = stq_8_bits_uop_prs2;
      5'b01001:
        casez_tmp_38 = stq_9_bits_uop_prs2;
      5'b01010:
        casez_tmp_38 = stq_10_bits_uop_prs2;
      5'b01011:
        casez_tmp_38 = stq_11_bits_uop_prs2;
      5'b01100:
        casez_tmp_38 = stq_12_bits_uop_prs2;
      5'b01101:
        casez_tmp_38 = stq_13_bits_uop_prs2;
      5'b01110:
        casez_tmp_38 = stq_14_bits_uop_prs2;
      5'b01111:
        casez_tmp_38 = stq_15_bits_uop_prs2;
      5'b10000:
        casez_tmp_38 = stq_16_bits_uop_prs2;
      5'b10001:
        casez_tmp_38 = stq_17_bits_uop_prs2;
      5'b10010:
        casez_tmp_38 = stq_18_bits_uop_prs2;
      5'b10011:
        casez_tmp_38 = stq_19_bits_uop_prs2;
      5'b10100:
        casez_tmp_38 = stq_20_bits_uop_prs2;
      5'b10101:
        casez_tmp_38 = stq_21_bits_uop_prs2;
      5'b10110:
        casez_tmp_38 = stq_22_bits_uop_prs2;
      5'b10111:
        casez_tmp_38 = stq_23_bits_uop_prs2;
      5'b11000:
        casez_tmp_38 = stq_24_bits_uop_prs2;
      5'b11001:
        casez_tmp_38 = stq_25_bits_uop_prs2;
      5'b11010:
        casez_tmp_38 = stq_26_bits_uop_prs2;
      5'b11011:
        casez_tmp_38 = stq_27_bits_uop_prs2;
      5'b11100:
        casez_tmp_38 = stq_28_bits_uop_prs2;
      5'b11101:
        casez_tmp_38 = stq_29_bits_uop_prs2;
      5'b11110:
        casez_tmp_38 = stq_30_bits_uop_prs2;
      default:
        casez_tmp_38 = stq_31_bits_uop_prs2;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_39;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_39 = stq_0_bits_uop_prs3;
      5'b00001:
        casez_tmp_39 = stq_1_bits_uop_prs3;
      5'b00010:
        casez_tmp_39 = stq_2_bits_uop_prs3;
      5'b00011:
        casez_tmp_39 = stq_3_bits_uop_prs3;
      5'b00100:
        casez_tmp_39 = stq_4_bits_uop_prs3;
      5'b00101:
        casez_tmp_39 = stq_5_bits_uop_prs3;
      5'b00110:
        casez_tmp_39 = stq_6_bits_uop_prs3;
      5'b00111:
        casez_tmp_39 = stq_7_bits_uop_prs3;
      5'b01000:
        casez_tmp_39 = stq_8_bits_uop_prs3;
      5'b01001:
        casez_tmp_39 = stq_9_bits_uop_prs3;
      5'b01010:
        casez_tmp_39 = stq_10_bits_uop_prs3;
      5'b01011:
        casez_tmp_39 = stq_11_bits_uop_prs3;
      5'b01100:
        casez_tmp_39 = stq_12_bits_uop_prs3;
      5'b01101:
        casez_tmp_39 = stq_13_bits_uop_prs3;
      5'b01110:
        casez_tmp_39 = stq_14_bits_uop_prs3;
      5'b01111:
        casez_tmp_39 = stq_15_bits_uop_prs3;
      5'b10000:
        casez_tmp_39 = stq_16_bits_uop_prs3;
      5'b10001:
        casez_tmp_39 = stq_17_bits_uop_prs3;
      5'b10010:
        casez_tmp_39 = stq_18_bits_uop_prs3;
      5'b10011:
        casez_tmp_39 = stq_19_bits_uop_prs3;
      5'b10100:
        casez_tmp_39 = stq_20_bits_uop_prs3;
      5'b10101:
        casez_tmp_39 = stq_21_bits_uop_prs3;
      5'b10110:
        casez_tmp_39 = stq_22_bits_uop_prs3;
      5'b10111:
        casez_tmp_39 = stq_23_bits_uop_prs3;
      5'b11000:
        casez_tmp_39 = stq_24_bits_uop_prs3;
      5'b11001:
        casez_tmp_39 = stq_25_bits_uop_prs3;
      5'b11010:
        casez_tmp_39 = stq_26_bits_uop_prs3;
      5'b11011:
        casez_tmp_39 = stq_27_bits_uop_prs3;
      5'b11100:
        casez_tmp_39 = stq_28_bits_uop_prs3;
      5'b11101:
        casez_tmp_39 = stq_29_bits_uop_prs3;
      5'b11110:
        casez_tmp_39 = stq_30_bits_uop_prs3;
      default:
        casez_tmp_39 = stq_31_bits_uop_prs3;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_40;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_40 = stq_0_bits_uop_ppred;
      5'b00001:
        casez_tmp_40 = stq_1_bits_uop_ppred;
      5'b00010:
        casez_tmp_40 = stq_2_bits_uop_ppred;
      5'b00011:
        casez_tmp_40 = stq_3_bits_uop_ppred;
      5'b00100:
        casez_tmp_40 = stq_4_bits_uop_ppred;
      5'b00101:
        casez_tmp_40 = stq_5_bits_uop_ppred;
      5'b00110:
        casez_tmp_40 = stq_6_bits_uop_ppred;
      5'b00111:
        casez_tmp_40 = stq_7_bits_uop_ppred;
      5'b01000:
        casez_tmp_40 = stq_8_bits_uop_ppred;
      5'b01001:
        casez_tmp_40 = stq_9_bits_uop_ppred;
      5'b01010:
        casez_tmp_40 = stq_10_bits_uop_ppred;
      5'b01011:
        casez_tmp_40 = stq_11_bits_uop_ppred;
      5'b01100:
        casez_tmp_40 = stq_12_bits_uop_ppred;
      5'b01101:
        casez_tmp_40 = stq_13_bits_uop_ppred;
      5'b01110:
        casez_tmp_40 = stq_14_bits_uop_ppred;
      5'b01111:
        casez_tmp_40 = stq_15_bits_uop_ppred;
      5'b10000:
        casez_tmp_40 = stq_16_bits_uop_ppred;
      5'b10001:
        casez_tmp_40 = stq_17_bits_uop_ppred;
      5'b10010:
        casez_tmp_40 = stq_18_bits_uop_ppred;
      5'b10011:
        casez_tmp_40 = stq_19_bits_uop_ppred;
      5'b10100:
        casez_tmp_40 = stq_20_bits_uop_ppred;
      5'b10101:
        casez_tmp_40 = stq_21_bits_uop_ppred;
      5'b10110:
        casez_tmp_40 = stq_22_bits_uop_ppred;
      5'b10111:
        casez_tmp_40 = stq_23_bits_uop_ppred;
      5'b11000:
        casez_tmp_40 = stq_24_bits_uop_ppred;
      5'b11001:
        casez_tmp_40 = stq_25_bits_uop_ppred;
      5'b11010:
        casez_tmp_40 = stq_26_bits_uop_ppred;
      5'b11011:
        casez_tmp_40 = stq_27_bits_uop_ppred;
      5'b11100:
        casez_tmp_40 = stq_28_bits_uop_ppred;
      5'b11101:
        casez_tmp_40 = stq_29_bits_uop_ppred;
      5'b11110:
        casez_tmp_40 = stq_30_bits_uop_ppred;
      default:
        casez_tmp_40 = stq_31_bits_uop_ppred;
    endcase
  end // always @(*)
  reg         casez_tmp_41;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_41 = stq_0_bits_uop_prs1_busy;
      5'b00001:
        casez_tmp_41 = stq_1_bits_uop_prs1_busy;
      5'b00010:
        casez_tmp_41 = stq_2_bits_uop_prs1_busy;
      5'b00011:
        casez_tmp_41 = stq_3_bits_uop_prs1_busy;
      5'b00100:
        casez_tmp_41 = stq_4_bits_uop_prs1_busy;
      5'b00101:
        casez_tmp_41 = stq_5_bits_uop_prs1_busy;
      5'b00110:
        casez_tmp_41 = stq_6_bits_uop_prs1_busy;
      5'b00111:
        casez_tmp_41 = stq_7_bits_uop_prs1_busy;
      5'b01000:
        casez_tmp_41 = stq_8_bits_uop_prs1_busy;
      5'b01001:
        casez_tmp_41 = stq_9_bits_uop_prs1_busy;
      5'b01010:
        casez_tmp_41 = stq_10_bits_uop_prs1_busy;
      5'b01011:
        casez_tmp_41 = stq_11_bits_uop_prs1_busy;
      5'b01100:
        casez_tmp_41 = stq_12_bits_uop_prs1_busy;
      5'b01101:
        casez_tmp_41 = stq_13_bits_uop_prs1_busy;
      5'b01110:
        casez_tmp_41 = stq_14_bits_uop_prs1_busy;
      5'b01111:
        casez_tmp_41 = stq_15_bits_uop_prs1_busy;
      5'b10000:
        casez_tmp_41 = stq_16_bits_uop_prs1_busy;
      5'b10001:
        casez_tmp_41 = stq_17_bits_uop_prs1_busy;
      5'b10010:
        casez_tmp_41 = stq_18_bits_uop_prs1_busy;
      5'b10011:
        casez_tmp_41 = stq_19_bits_uop_prs1_busy;
      5'b10100:
        casez_tmp_41 = stq_20_bits_uop_prs1_busy;
      5'b10101:
        casez_tmp_41 = stq_21_bits_uop_prs1_busy;
      5'b10110:
        casez_tmp_41 = stq_22_bits_uop_prs1_busy;
      5'b10111:
        casez_tmp_41 = stq_23_bits_uop_prs1_busy;
      5'b11000:
        casez_tmp_41 = stq_24_bits_uop_prs1_busy;
      5'b11001:
        casez_tmp_41 = stq_25_bits_uop_prs1_busy;
      5'b11010:
        casez_tmp_41 = stq_26_bits_uop_prs1_busy;
      5'b11011:
        casez_tmp_41 = stq_27_bits_uop_prs1_busy;
      5'b11100:
        casez_tmp_41 = stq_28_bits_uop_prs1_busy;
      5'b11101:
        casez_tmp_41 = stq_29_bits_uop_prs1_busy;
      5'b11110:
        casez_tmp_41 = stq_30_bits_uop_prs1_busy;
      default:
        casez_tmp_41 = stq_31_bits_uop_prs1_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_42;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_42 = stq_0_bits_uop_prs2_busy;
      5'b00001:
        casez_tmp_42 = stq_1_bits_uop_prs2_busy;
      5'b00010:
        casez_tmp_42 = stq_2_bits_uop_prs2_busy;
      5'b00011:
        casez_tmp_42 = stq_3_bits_uop_prs2_busy;
      5'b00100:
        casez_tmp_42 = stq_4_bits_uop_prs2_busy;
      5'b00101:
        casez_tmp_42 = stq_5_bits_uop_prs2_busy;
      5'b00110:
        casez_tmp_42 = stq_6_bits_uop_prs2_busy;
      5'b00111:
        casez_tmp_42 = stq_7_bits_uop_prs2_busy;
      5'b01000:
        casez_tmp_42 = stq_8_bits_uop_prs2_busy;
      5'b01001:
        casez_tmp_42 = stq_9_bits_uop_prs2_busy;
      5'b01010:
        casez_tmp_42 = stq_10_bits_uop_prs2_busy;
      5'b01011:
        casez_tmp_42 = stq_11_bits_uop_prs2_busy;
      5'b01100:
        casez_tmp_42 = stq_12_bits_uop_prs2_busy;
      5'b01101:
        casez_tmp_42 = stq_13_bits_uop_prs2_busy;
      5'b01110:
        casez_tmp_42 = stq_14_bits_uop_prs2_busy;
      5'b01111:
        casez_tmp_42 = stq_15_bits_uop_prs2_busy;
      5'b10000:
        casez_tmp_42 = stq_16_bits_uop_prs2_busy;
      5'b10001:
        casez_tmp_42 = stq_17_bits_uop_prs2_busy;
      5'b10010:
        casez_tmp_42 = stq_18_bits_uop_prs2_busy;
      5'b10011:
        casez_tmp_42 = stq_19_bits_uop_prs2_busy;
      5'b10100:
        casez_tmp_42 = stq_20_bits_uop_prs2_busy;
      5'b10101:
        casez_tmp_42 = stq_21_bits_uop_prs2_busy;
      5'b10110:
        casez_tmp_42 = stq_22_bits_uop_prs2_busy;
      5'b10111:
        casez_tmp_42 = stq_23_bits_uop_prs2_busy;
      5'b11000:
        casez_tmp_42 = stq_24_bits_uop_prs2_busy;
      5'b11001:
        casez_tmp_42 = stq_25_bits_uop_prs2_busy;
      5'b11010:
        casez_tmp_42 = stq_26_bits_uop_prs2_busy;
      5'b11011:
        casez_tmp_42 = stq_27_bits_uop_prs2_busy;
      5'b11100:
        casez_tmp_42 = stq_28_bits_uop_prs2_busy;
      5'b11101:
        casez_tmp_42 = stq_29_bits_uop_prs2_busy;
      5'b11110:
        casez_tmp_42 = stq_30_bits_uop_prs2_busy;
      default:
        casez_tmp_42 = stq_31_bits_uop_prs2_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_43;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_43 = stq_0_bits_uop_prs3_busy;
      5'b00001:
        casez_tmp_43 = stq_1_bits_uop_prs3_busy;
      5'b00010:
        casez_tmp_43 = stq_2_bits_uop_prs3_busy;
      5'b00011:
        casez_tmp_43 = stq_3_bits_uop_prs3_busy;
      5'b00100:
        casez_tmp_43 = stq_4_bits_uop_prs3_busy;
      5'b00101:
        casez_tmp_43 = stq_5_bits_uop_prs3_busy;
      5'b00110:
        casez_tmp_43 = stq_6_bits_uop_prs3_busy;
      5'b00111:
        casez_tmp_43 = stq_7_bits_uop_prs3_busy;
      5'b01000:
        casez_tmp_43 = stq_8_bits_uop_prs3_busy;
      5'b01001:
        casez_tmp_43 = stq_9_bits_uop_prs3_busy;
      5'b01010:
        casez_tmp_43 = stq_10_bits_uop_prs3_busy;
      5'b01011:
        casez_tmp_43 = stq_11_bits_uop_prs3_busy;
      5'b01100:
        casez_tmp_43 = stq_12_bits_uop_prs3_busy;
      5'b01101:
        casez_tmp_43 = stq_13_bits_uop_prs3_busy;
      5'b01110:
        casez_tmp_43 = stq_14_bits_uop_prs3_busy;
      5'b01111:
        casez_tmp_43 = stq_15_bits_uop_prs3_busy;
      5'b10000:
        casez_tmp_43 = stq_16_bits_uop_prs3_busy;
      5'b10001:
        casez_tmp_43 = stq_17_bits_uop_prs3_busy;
      5'b10010:
        casez_tmp_43 = stq_18_bits_uop_prs3_busy;
      5'b10011:
        casez_tmp_43 = stq_19_bits_uop_prs3_busy;
      5'b10100:
        casez_tmp_43 = stq_20_bits_uop_prs3_busy;
      5'b10101:
        casez_tmp_43 = stq_21_bits_uop_prs3_busy;
      5'b10110:
        casez_tmp_43 = stq_22_bits_uop_prs3_busy;
      5'b10111:
        casez_tmp_43 = stq_23_bits_uop_prs3_busy;
      5'b11000:
        casez_tmp_43 = stq_24_bits_uop_prs3_busy;
      5'b11001:
        casez_tmp_43 = stq_25_bits_uop_prs3_busy;
      5'b11010:
        casez_tmp_43 = stq_26_bits_uop_prs3_busy;
      5'b11011:
        casez_tmp_43 = stq_27_bits_uop_prs3_busy;
      5'b11100:
        casez_tmp_43 = stq_28_bits_uop_prs3_busy;
      5'b11101:
        casez_tmp_43 = stq_29_bits_uop_prs3_busy;
      5'b11110:
        casez_tmp_43 = stq_30_bits_uop_prs3_busy;
      default:
        casez_tmp_43 = stq_31_bits_uop_prs3_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_44;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_44 = stq_0_bits_uop_ppred_busy;
      5'b00001:
        casez_tmp_44 = stq_1_bits_uop_ppred_busy;
      5'b00010:
        casez_tmp_44 = stq_2_bits_uop_ppred_busy;
      5'b00011:
        casez_tmp_44 = stq_3_bits_uop_ppred_busy;
      5'b00100:
        casez_tmp_44 = stq_4_bits_uop_ppred_busy;
      5'b00101:
        casez_tmp_44 = stq_5_bits_uop_ppred_busy;
      5'b00110:
        casez_tmp_44 = stq_6_bits_uop_ppred_busy;
      5'b00111:
        casez_tmp_44 = stq_7_bits_uop_ppred_busy;
      5'b01000:
        casez_tmp_44 = stq_8_bits_uop_ppred_busy;
      5'b01001:
        casez_tmp_44 = stq_9_bits_uop_ppred_busy;
      5'b01010:
        casez_tmp_44 = stq_10_bits_uop_ppred_busy;
      5'b01011:
        casez_tmp_44 = stq_11_bits_uop_ppred_busy;
      5'b01100:
        casez_tmp_44 = stq_12_bits_uop_ppred_busy;
      5'b01101:
        casez_tmp_44 = stq_13_bits_uop_ppred_busy;
      5'b01110:
        casez_tmp_44 = stq_14_bits_uop_ppred_busy;
      5'b01111:
        casez_tmp_44 = stq_15_bits_uop_ppred_busy;
      5'b10000:
        casez_tmp_44 = stq_16_bits_uop_ppred_busy;
      5'b10001:
        casez_tmp_44 = stq_17_bits_uop_ppred_busy;
      5'b10010:
        casez_tmp_44 = stq_18_bits_uop_ppred_busy;
      5'b10011:
        casez_tmp_44 = stq_19_bits_uop_ppred_busy;
      5'b10100:
        casez_tmp_44 = stq_20_bits_uop_ppred_busy;
      5'b10101:
        casez_tmp_44 = stq_21_bits_uop_ppred_busy;
      5'b10110:
        casez_tmp_44 = stq_22_bits_uop_ppred_busy;
      5'b10111:
        casez_tmp_44 = stq_23_bits_uop_ppred_busy;
      5'b11000:
        casez_tmp_44 = stq_24_bits_uop_ppred_busy;
      5'b11001:
        casez_tmp_44 = stq_25_bits_uop_ppred_busy;
      5'b11010:
        casez_tmp_44 = stq_26_bits_uop_ppred_busy;
      5'b11011:
        casez_tmp_44 = stq_27_bits_uop_ppred_busy;
      5'b11100:
        casez_tmp_44 = stq_28_bits_uop_ppred_busy;
      5'b11101:
        casez_tmp_44 = stq_29_bits_uop_ppred_busy;
      5'b11110:
        casez_tmp_44 = stq_30_bits_uop_ppred_busy;
      default:
        casez_tmp_44 = stq_31_bits_uop_ppred_busy;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_45;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_45 = stq_0_bits_uop_stale_pdst;
      5'b00001:
        casez_tmp_45 = stq_1_bits_uop_stale_pdst;
      5'b00010:
        casez_tmp_45 = stq_2_bits_uop_stale_pdst;
      5'b00011:
        casez_tmp_45 = stq_3_bits_uop_stale_pdst;
      5'b00100:
        casez_tmp_45 = stq_4_bits_uop_stale_pdst;
      5'b00101:
        casez_tmp_45 = stq_5_bits_uop_stale_pdst;
      5'b00110:
        casez_tmp_45 = stq_6_bits_uop_stale_pdst;
      5'b00111:
        casez_tmp_45 = stq_7_bits_uop_stale_pdst;
      5'b01000:
        casez_tmp_45 = stq_8_bits_uop_stale_pdst;
      5'b01001:
        casez_tmp_45 = stq_9_bits_uop_stale_pdst;
      5'b01010:
        casez_tmp_45 = stq_10_bits_uop_stale_pdst;
      5'b01011:
        casez_tmp_45 = stq_11_bits_uop_stale_pdst;
      5'b01100:
        casez_tmp_45 = stq_12_bits_uop_stale_pdst;
      5'b01101:
        casez_tmp_45 = stq_13_bits_uop_stale_pdst;
      5'b01110:
        casez_tmp_45 = stq_14_bits_uop_stale_pdst;
      5'b01111:
        casez_tmp_45 = stq_15_bits_uop_stale_pdst;
      5'b10000:
        casez_tmp_45 = stq_16_bits_uop_stale_pdst;
      5'b10001:
        casez_tmp_45 = stq_17_bits_uop_stale_pdst;
      5'b10010:
        casez_tmp_45 = stq_18_bits_uop_stale_pdst;
      5'b10011:
        casez_tmp_45 = stq_19_bits_uop_stale_pdst;
      5'b10100:
        casez_tmp_45 = stq_20_bits_uop_stale_pdst;
      5'b10101:
        casez_tmp_45 = stq_21_bits_uop_stale_pdst;
      5'b10110:
        casez_tmp_45 = stq_22_bits_uop_stale_pdst;
      5'b10111:
        casez_tmp_45 = stq_23_bits_uop_stale_pdst;
      5'b11000:
        casez_tmp_45 = stq_24_bits_uop_stale_pdst;
      5'b11001:
        casez_tmp_45 = stq_25_bits_uop_stale_pdst;
      5'b11010:
        casez_tmp_45 = stq_26_bits_uop_stale_pdst;
      5'b11011:
        casez_tmp_45 = stq_27_bits_uop_stale_pdst;
      5'b11100:
        casez_tmp_45 = stq_28_bits_uop_stale_pdst;
      5'b11101:
        casez_tmp_45 = stq_29_bits_uop_stale_pdst;
      5'b11110:
        casez_tmp_45 = stq_30_bits_uop_stale_pdst;
      default:
        casez_tmp_45 = stq_31_bits_uop_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_46;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_46 = stq_0_bits_uop_exception;
      5'b00001:
        casez_tmp_46 = stq_1_bits_uop_exception;
      5'b00010:
        casez_tmp_46 = stq_2_bits_uop_exception;
      5'b00011:
        casez_tmp_46 = stq_3_bits_uop_exception;
      5'b00100:
        casez_tmp_46 = stq_4_bits_uop_exception;
      5'b00101:
        casez_tmp_46 = stq_5_bits_uop_exception;
      5'b00110:
        casez_tmp_46 = stq_6_bits_uop_exception;
      5'b00111:
        casez_tmp_46 = stq_7_bits_uop_exception;
      5'b01000:
        casez_tmp_46 = stq_8_bits_uop_exception;
      5'b01001:
        casez_tmp_46 = stq_9_bits_uop_exception;
      5'b01010:
        casez_tmp_46 = stq_10_bits_uop_exception;
      5'b01011:
        casez_tmp_46 = stq_11_bits_uop_exception;
      5'b01100:
        casez_tmp_46 = stq_12_bits_uop_exception;
      5'b01101:
        casez_tmp_46 = stq_13_bits_uop_exception;
      5'b01110:
        casez_tmp_46 = stq_14_bits_uop_exception;
      5'b01111:
        casez_tmp_46 = stq_15_bits_uop_exception;
      5'b10000:
        casez_tmp_46 = stq_16_bits_uop_exception;
      5'b10001:
        casez_tmp_46 = stq_17_bits_uop_exception;
      5'b10010:
        casez_tmp_46 = stq_18_bits_uop_exception;
      5'b10011:
        casez_tmp_46 = stq_19_bits_uop_exception;
      5'b10100:
        casez_tmp_46 = stq_20_bits_uop_exception;
      5'b10101:
        casez_tmp_46 = stq_21_bits_uop_exception;
      5'b10110:
        casez_tmp_46 = stq_22_bits_uop_exception;
      5'b10111:
        casez_tmp_46 = stq_23_bits_uop_exception;
      5'b11000:
        casez_tmp_46 = stq_24_bits_uop_exception;
      5'b11001:
        casez_tmp_46 = stq_25_bits_uop_exception;
      5'b11010:
        casez_tmp_46 = stq_26_bits_uop_exception;
      5'b11011:
        casez_tmp_46 = stq_27_bits_uop_exception;
      5'b11100:
        casez_tmp_46 = stq_28_bits_uop_exception;
      5'b11101:
        casez_tmp_46 = stq_29_bits_uop_exception;
      5'b11110:
        casez_tmp_46 = stq_30_bits_uop_exception;
      default:
        casez_tmp_46 = stq_31_bits_uop_exception;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_47;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_47 = stq_0_bits_uop_exc_cause;
      5'b00001:
        casez_tmp_47 = stq_1_bits_uop_exc_cause;
      5'b00010:
        casez_tmp_47 = stq_2_bits_uop_exc_cause;
      5'b00011:
        casez_tmp_47 = stq_3_bits_uop_exc_cause;
      5'b00100:
        casez_tmp_47 = stq_4_bits_uop_exc_cause;
      5'b00101:
        casez_tmp_47 = stq_5_bits_uop_exc_cause;
      5'b00110:
        casez_tmp_47 = stq_6_bits_uop_exc_cause;
      5'b00111:
        casez_tmp_47 = stq_7_bits_uop_exc_cause;
      5'b01000:
        casez_tmp_47 = stq_8_bits_uop_exc_cause;
      5'b01001:
        casez_tmp_47 = stq_9_bits_uop_exc_cause;
      5'b01010:
        casez_tmp_47 = stq_10_bits_uop_exc_cause;
      5'b01011:
        casez_tmp_47 = stq_11_bits_uop_exc_cause;
      5'b01100:
        casez_tmp_47 = stq_12_bits_uop_exc_cause;
      5'b01101:
        casez_tmp_47 = stq_13_bits_uop_exc_cause;
      5'b01110:
        casez_tmp_47 = stq_14_bits_uop_exc_cause;
      5'b01111:
        casez_tmp_47 = stq_15_bits_uop_exc_cause;
      5'b10000:
        casez_tmp_47 = stq_16_bits_uop_exc_cause;
      5'b10001:
        casez_tmp_47 = stq_17_bits_uop_exc_cause;
      5'b10010:
        casez_tmp_47 = stq_18_bits_uop_exc_cause;
      5'b10011:
        casez_tmp_47 = stq_19_bits_uop_exc_cause;
      5'b10100:
        casez_tmp_47 = stq_20_bits_uop_exc_cause;
      5'b10101:
        casez_tmp_47 = stq_21_bits_uop_exc_cause;
      5'b10110:
        casez_tmp_47 = stq_22_bits_uop_exc_cause;
      5'b10111:
        casez_tmp_47 = stq_23_bits_uop_exc_cause;
      5'b11000:
        casez_tmp_47 = stq_24_bits_uop_exc_cause;
      5'b11001:
        casez_tmp_47 = stq_25_bits_uop_exc_cause;
      5'b11010:
        casez_tmp_47 = stq_26_bits_uop_exc_cause;
      5'b11011:
        casez_tmp_47 = stq_27_bits_uop_exc_cause;
      5'b11100:
        casez_tmp_47 = stq_28_bits_uop_exc_cause;
      5'b11101:
        casez_tmp_47 = stq_29_bits_uop_exc_cause;
      5'b11110:
        casez_tmp_47 = stq_30_bits_uop_exc_cause;
      default:
        casez_tmp_47 = stq_31_bits_uop_exc_cause;
    endcase
  end // always @(*)
  reg         casez_tmp_48;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_48 = stq_0_bits_uop_bypassable;
      5'b00001:
        casez_tmp_48 = stq_1_bits_uop_bypassable;
      5'b00010:
        casez_tmp_48 = stq_2_bits_uop_bypassable;
      5'b00011:
        casez_tmp_48 = stq_3_bits_uop_bypassable;
      5'b00100:
        casez_tmp_48 = stq_4_bits_uop_bypassable;
      5'b00101:
        casez_tmp_48 = stq_5_bits_uop_bypassable;
      5'b00110:
        casez_tmp_48 = stq_6_bits_uop_bypassable;
      5'b00111:
        casez_tmp_48 = stq_7_bits_uop_bypassable;
      5'b01000:
        casez_tmp_48 = stq_8_bits_uop_bypassable;
      5'b01001:
        casez_tmp_48 = stq_9_bits_uop_bypassable;
      5'b01010:
        casez_tmp_48 = stq_10_bits_uop_bypassable;
      5'b01011:
        casez_tmp_48 = stq_11_bits_uop_bypassable;
      5'b01100:
        casez_tmp_48 = stq_12_bits_uop_bypassable;
      5'b01101:
        casez_tmp_48 = stq_13_bits_uop_bypassable;
      5'b01110:
        casez_tmp_48 = stq_14_bits_uop_bypassable;
      5'b01111:
        casez_tmp_48 = stq_15_bits_uop_bypassable;
      5'b10000:
        casez_tmp_48 = stq_16_bits_uop_bypassable;
      5'b10001:
        casez_tmp_48 = stq_17_bits_uop_bypassable;
      5'b10010:
        casez_tmp_48 = stq_18_bits_uop_bypassable;
      5'b10011:
        casez_tmp_48 = stq_19_bits_uop_bypassable;
      5'b10100:
        casez_tmp_48 = stq_20_bits_uop_bypassable;
      5'b10101:
        casez_tmp_48 = stq_21_bits_uop_bypassable;
      5'b10110:
        casez_tmp_48 = stq_22_bits_uop_bypassable;
      5'b10111:
        casez_tmp_48 = stq_23_bits_uop_bypassable;
      5'b11000:
        casez_tmp_48 = stq_24_bits_uop_bypassable;
      5'b11001:
        casez_tmp_48 = stq_25_bits_uop_bypassable;
      5'b11010:
        casez_tmp_48 = stq_26_bits_uop_bypassable;
      5'b11011:
        casez_tmp_48 = stq_27_bits_uop_bypassable;
      5'b11100:
        casez_tmp_48 = stq_28_bits_uop_bypassable;
      5'b11101:
        casez_tmp_48 = stq_29_bits_uop_bypassable;
      5'b11110:
        casez_tmp_48 = stq_30_bits_uop_bypassable;
      default:
        casez_tmp_48 = stq_31_bits_uop_bypassable;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_49;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_49 = stq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_49 = stq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_49 = stq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_49 = stq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_49 = stq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_49 = stq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_49 = stq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_49 = stq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_49 = stq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_49 = stq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_49 = stq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_49 = stq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_49 = stq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_49 = stq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_49 = stq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_49 = stq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_49 = stq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_49 = stq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_49 = stq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_49 = stq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_49 = stq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_49 = stq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_49 = stq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_49 = stq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_49 = stq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_49 = stq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_49 = stq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_49 = stq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_49 = stq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_49 = stq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_49 = stq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_49 = stq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_50;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_50 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_50 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_50 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_50 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_50 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_50 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_50 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_50 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_50 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_50 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_50 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_50 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_50 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_50 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_50 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_50 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_50 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_50 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_50 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_50 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_50 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_50 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_50 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_50 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_50 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_50 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_50 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_50 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_50 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_50 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_50 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_50 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_51;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_51 = stq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_51 = stq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_51 = stq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_51 = stq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_51 = stq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_51 = stq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_51 = stq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_51 = stq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_51 = stq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_51 = stq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_51 = stq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_51 = stq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_51 = stq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_51 = stq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_51 = stq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_51 = stq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_51 = stq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_51 = stq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_51 = stq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_51 = stq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_51 = stq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_51 = stq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_51 = stq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_51 = stq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_51 = stq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_51 = stq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_51 = stq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_51 = stq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_51 = stq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_51 = stq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_51 = stq_30_bits_uop_mem_signed;
      default:
        casez_tmp_51 = stq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  reg         casez_tmp_52;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_52 = stq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_52 = stq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_52 = stq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_52 = stq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_52 = stq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_52 = stq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_52 = stq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_52 = stq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_52 = stq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_52 = stq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_52 = stq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_52 = stq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_52 = stq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_52 = stq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_52 = stq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_52 = stq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_52 = stq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_52 = stq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_52 = stq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_52 = stq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_52 = stq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_52 = stq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_52 = stq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_52 = stq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_52 = stq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_52 = stq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_52 = stq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_52 = stq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_52 = stq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_52 = stq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_52 = stq_30_bits_uop_is_fence;
      default:
        casez_tmp_52 = stq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  reg         casez_tmp_53;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_53 = stq_0_bits_uop_is_fencei;
      5'b00001:
        casez_tmp_53 = stq_1_bits_uop_is_fencei;
      5'b00010:
        casez_tmp_53 = stq_2_bits_uop_is_fencei;
      5'b00011:
        casez_tmp_53 = stq_3_bits_uop_is_fencei;
      5'b00100:
        casez_tmp_53 = stq_4_bits_uop_is_fencei;
      5'b00101:
        casez_tmp_53 = stq_5_bits_uop_is_fencei;
      5'b00110:
        casez_tmp_53 = stq_6_bits_uop_is_fencei;
      5'b00111:
        casez_tmp_53 = stq_7_bits_uop_is_fencei;
      5'b01000:
        casez_tmp_53 = stq_8_bits_uop_is_fencei;
      5'b01001:
        casez_tmp_53 = stq_9_bits_uop_is_fencei;
      5'b01010:
        casez_tmp_53 = stq_10_bits_uop_is_fencei;
      5'b01011:
        casez_tmp_53 = stq_11_bits_uop_is_fencei;
      5'b01100:
        casez_tmp_53 = stq_12_bits_uop_is_fencei;
      5'b01101:
        casez_tmp_53 = stq_13_bits_uop_is_fencei;
      5'b01110:
        casez_tmp_53 = stq_14_bits_uop_is_fencei;
      5'b01111:
        casez_tmp_53 = stq_15_bits_uop_is_fencei;
      5'b10000:
        casez_tmp_53 = stq_16_bits_uop_is_fencei;
      5'b10001:
        casez_tmp_53 = stq_17_bits_uop_is_fencei;
      5'b10010:
        casez_tmp_53 = stq_18_bits_uop_is_fencei;
      5'b10011:
        casez_tmp_53 = stq_19_bits_uop_is_fencei;
      5'b10100:
        casez_tmp_53 = stq_20_bits_uop_is_fencei;
      5'b10101:
        casez_tmp_53 = stq_21_bits_uop_is_fencei;
      5'b10110:
        casez_tmp_53 = stq_22_bits_uop_is_fencei;
      5'b10111:
        casez_tmp_53 = stq_23_bits_uop_is_fencei;
      5'b11000:
        casez_tmp_53 = stq_24_bits_uop_is_fencei;
      5'b11001:
        casez_tmp_53 = stq_25_bits_uop_is_fencei;
      5'b11010:
        casez_tmp_53 = stq_26_bits_uop_is_fencei;
      5'b11011:
        casez_tmp_53 = stq_27_bits_uop_is_fencei;
      5'b11100:
        casez_tmp_53 = stq_28_bits_uop_is_fencei;
      5'b11101:
        casez_tmp_53 = stq_29_bits_uop_is_fencei;
      5'b11110:
        casez_tmp_53 = stq_30_bits_uop_is_fencei;
      default:
        casez_tmp_53 = stq_31_bits_uop_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_54;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_54 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_54 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_54 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_54 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_54 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_54 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_54 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_54 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_54 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_54 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_54 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_54 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_54 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_54 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_54 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_54 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_54 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_54 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_54 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_54 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_54 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_54 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_54 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_54 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_54 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_54 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_54 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_54 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_54 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_54 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_54 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_54 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_55;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_55 = stq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_55 = stq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_55 = stq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_55 = stq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_55 = stq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_55 = stq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_55 = stq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_55 = stq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_55 = stq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_55 = stq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_55 = stq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_55 = stq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_55 = stq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_55 = stq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_55 = stq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_55 = stq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_55 = stq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_55 = stq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_55 = stq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_55 = stq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_55 = stq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_55 = stq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_55 = stq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_55 = stq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_55 = stq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_55 = stq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_55 = stq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_55 = stq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_55 = stq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_55 = stq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_55 = stq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_55 = stq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_56;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_56 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_56 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_56 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_56 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_56 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_56 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_56 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_56 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_56 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_56 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_56 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_56 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_56 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_56 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_56 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_56 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_56 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_56 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_56 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_56 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_56 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_56 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_56 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_56 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_56 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_56 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_56 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_56 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_56 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_56 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_56 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_56 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_57;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_57 = stq_0_bits_uop_is_sys_pc2epc;
      5'b00001:
        casez_tmp_57 = stq_1_bits_uop_is_sys_pc2epc;
      5'b00010:
        casez_tmp_57 = stq_2_bits_uop_is_sys_pc2epc;
      5'b00011:
        casez_tmp_57 = stq_3_bits_uop_is_sys_pc2epc;
      5'b00100:
        casez_tmp_57 = stq_4_bits_uop_is_sys_pc2epc;
      5'b00101:
        casez_tmp_57 = stq_5_bits_uop_is_sys_pc2epc;
      5'b00110:
        casez_tmp_57 = stq_6_bits_uop_is_sys_pc2epc;
      5'b00111:
        casez_tmp_57 = stq_7_bits_uop_is_sys_pc2epc;
      5'b01000:
        casez_tmp_57 = stq_8_bits_uop_is_sys_pc2epc;
      5'b01001:
        casez_tmp_57 = stq_9_bits_uop_is_sys_pc2epc;
      5'b01010:
        casez_tmp_57 = stq_10_bits_uop_is_sys_pc2epc;
      5'b01011:
        casez_tmp_57 = stq_11_bits_uop_is_sys_pc2epc;
      5'b01100:
        casez_tmp_57 = stq_12_bits_uop_is_sys_pc2epc;
      5'b01101:
        casez_tmp_57 = stq_13_bits_uop_is_sys_pc2epc;
      5'b01110:
        casez_tmp_57 = stq_14_bits_uop_is_sys_pc2epc;
      5'b01111:
        casez_tmp_57 = stq_15_bits_uop_is_sys_pc2epc;
      5'b10000:
        casez_tmp_57 = stq_16_bits_uop_is_sys_pc2epc;
      5'b10001:
        casez_tmp_57 = stq_17_bits_uop_is_sys_pc2epc;
      5'b10010:
        casez_tmp_57 = stq_18_bits_uop_is_sys_pc2epc;
      5'b10011:
        casez_tmp_57 = stq_19_bits_uop_is_sys_pc2epc;
      5'b10100:
        casez_tmp_57 = stq_20_bits_uop_is_sys_pc2epc;
      5'b10101:
        casez_tmp_57 = stq_21_bits_uop_is_sys_pc2epc;
      5'b10110:
        casez_tmp_57 = stq_22_bits_uop_is_sys_pc2epc;
      5'b10111:
        casez_tmp_57 = stq_23_bits_uop_is_sys_pc2epc;
      5'b11000:
        casez_tmp_57 = stq_24_bits_uop_is_sys_pc2epc;
      5'b11001:
        casez_tmp_57 = stq_25_bits_uop_is_sys_pc2epc;
      5'b11010:
        casez_tmp_57 = stq_26_bits_uop_is_sys_pc2epc;
      5'b11011:
        casez_tmp_57 = stq_27_bits_uop_is_sys_pc2epc;
      5'b11100:
        casez_tmp_57 = stq_28_bits_uop_is_sys_pc2epc;
      5'b11101:
        casez_tmp_57 = stq_29_bits_uop_is_sys_pc2epc;
      5'b11110:
        casez_tmp_57 = stq_30_bits_uop_is_sys_pc2epc;
      default:
        casez_tmp_57 = stq_31_bits_uop_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_58;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_58 = stq_0_bits_uop_is_unique;
      5'b00001:
        casez_tmp_58 = stq_1_bits_uop_is_unique;
      5'b00010:
        casez_tmp_58 = stq_2_bits_uop_is_unique;
      5'b00011:
        casez_tmp_58 = stq_3_bits_uop_is_unique;
      5'b00100:
        casez_tmp_58 = stq_4_bits_uop_is_unique;
      5'b00101:
        casez_tmp_58 = stq_5_bits_uop_is_unique;
      5'b00110:
        casez_tmp_58 = stq_6_bits_uop_is_unique;
      5'b00111:
        casez_tmp_58 = stq_7_bits_uop_is_unique;
      5'b01000:
        casez_tmp_58 = stq_8_bits_uop_is_unique;
      5'b01001:
        casez_tmp_58 = stq_9_bits_uop_is_unique;
      5'b01010:
        casez_tmp_58 = stq_10_bits_uop_is_unique;
      5'b01011:
        casez_tmp_58 = stq_11_bits_uop_is_unique;
      5'b01100:
        casez_tmp_58 = stq_12_bits_uop_is_unique;
      5'b01101:
        casez_tmp_58 = stq_13_bits_uop_is_unique;
      5'b01110:
        casez_tmp_58 = stq_14_bits_uop_is_unique;
      5'b01111:
        casez_tmp_58 = stq_15_bits_uop_is_unique;
      5'b10000:
        casez_tmp_58 = stq_16_bits_uop_is_unique;
      5'b10001:
        casez_tmp_58 = stq_17_bits_uop_is_unique;
      5'b10010:
        casez_tmp_58 = stq_18_bits_uop_is_unique;
      5'b10011:
        casez_tmp_58 = stq_19_bits_uop_is_unique;
      5'b10100:
        casez_tmp_58 = stq_20_bits_uop_is_unique;
      5'b10101:
        casez_tmp_58 = stq_21_bits_uop_is_unique;
      5'b10110:
        casez_tmp_58 = stq_22_bits_uop_is_unique;
      5'b10111:
        casez_tmp_58 = stq_23_bits_uop_is_unique;
      5'b11000:
        casez_tmp_58 = stq_24_bits_uop_is_unique;
      5'b11001:
        casez_tmp_58 = stq_25_bits_uop_is_unique;
      5'b11010:
        casez_tmp_58 = stq_26_bits_uop_is_unique;
      5'b11011:
        casez_tmp_58 = stq_27_bits_uop_is_unique;
      5'b11100:
        casez_tmp_58 = stq_28_bits_uop_is_unique;
      5'b11101:
        casez_tmp_58 = stq_29_bits_uop_is_unique;
      5'b11110:
        casez_tmp_58 = stq_30_bits_uop_is_unique;
      default:
        casez_tmp_58 = stq_31_bits_uop_is_unique;
    endcase
  end // always @(*)
  reg         casez_tmp_59;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_59 = stq_0_bits_uop_flush_on_commit;
      5'b00001:
        casez_tmp_59 = stq_1_bits_uop_flush_on_commit;
      5'b00010:
        casez_tmp_59 = stq_2_bits_uop_flush_on_commit;
      5'b00011:
        casez_tmp_59 = stq_3_bits_uop_flush_on_commit;
      5'b00100:
        casez_tmp_59 = stq_4_bits_uop_flush_on_commit;
      5'b00101:
        casez_tmp_59 = stq_5_bits_uop_flush_on_commit;
      5'b00110:
        casez_tmp_59 = stq_6_bits_uop_flush_on_commit;
      5'b00111:
        casez_tmp_59 = stq_7_bits_uop_flush_on_commit;
      5'b01000:
        casez_tmp_59 = stq_8_bits_uop_flush_on_commit;
      5'b01001:
        casez_tmp_59 = stq_9_bits_uop_flush_on_commit;
      5'b01010:
        casez_tmp_59 = stq_10_bits_uop_flush_on_commit;
      5'b01011:
        casez_tmp_59 = stq_11_bits_uop_flush_on_commit;
      5'b01100:
        casez_tmp_59 = stq_12_bits_uop_flush_on_commit;
      5'b01101:
        casez_tmp_59 = stq_13_bits_uop_flush_on_commit;
      5'b01110:
        casez_tmp_59 = stq_14_bits_uop_flush_on_commit;
      5'b01111:
        casez_tmp_59 = stq_15_bits_uop_flush_on_commit;
      5'b10000:
        casez_tmp_59 = stq_16_bits_uop_flush_on_commit;
      5'b10001:
        casez_tmp_59 = stq_17_bits_uop_flush_on_commit;
      5'b10010:
        casez_tmp_59 = stq_18_bits_uop_flush_on_commit;
      5'b10011:
        casez_tmp_59 = stq_19_bits_uop_flush_on_commit;
      5'b10100:
        casez_tmp_59 = stq_20_bits_uop_flush_on_commit;
      5'b10101:
        casez_tmp_59 = stq_21_bits_uop_flush_on_commit;
      5'b10110:
        casez_tmp_59 = stq_22_bits_uop_flush_on_commit;
      5'b10111:
        casez_tmp_59 = stq_23_bits_uop_flush_on_commit;
      5'b11000:
        casez_tmp_59 = stq_24_bits_uop_flush_on_commit;
      5'b11001:
        casez_tmp_59 = stq_25_bits_uop_flush_on_commit;
      5'b11010:
        casez_tmp_59 = stq_26_bits_uop_flush_on_commit;
      5'b11011:
        casez_tmp_59 = stq_27_bits_uop_flush_on_commit;
      5'b11100:
        casez_tmp_59 = stq_28_bits_uop_flush_on_commit;
      5'b11101:
        casez_tmp_59 = stq_29_bits_uop_flush_on_commit;
      5'b11110:
        casez_tmp_59 = stq_30_bits_uop_flush_on_commit;
      default:
        casez_tmp_59 = stq_31_bits_uop_flush_on_commit;
    endcase
  end // always @(*)
  reg         casez_tmp_60;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_60 = stq_0_bits_uop_ldst_is_rs1;
      5'b00001:
        casez_tmp_60 = stq_1_bits_uop_ldst_is_rs1;
      5'b00010:
        casez_tmp_60 = stq_2_bits_uop_ldst_is_rs1;
      5'b00011:
        casez_tmp_60 = stq_3_bits_uop_ldst_is_rs1;
      5'b00100:
        casez_tmp_60 = stq_4_bits_uop_ldst_is_rs1;
      5'b00101:
        casez_tmp_60 = stq_5_bits_uop_ldst_is_rs1;
      5'b00110:
        casez_tmp_60 = stq_6_bits_uop_ldst_is_rs1;
      5'b00111:
        casez_tmp_60 = stq_7_bits_uop_ldst_is_rs1;
      5'b01000:
        casez_tmp_60 = stq_8_bits_uop_ldst_is_rs1;
      5'b01001:
        casez_tmp_60 = stq_9_bits_uop_ldst_is_rs1;
      5'b01010:
        casez_tmp_60 = stq_10_bits_uop_ldst_is_rs1;
      5'b01011:
        casez_tmp_60 = stq_11_bits_uop_ldst_is_rs1;
      5'b01100:
        casez_tmp_60 = stq_12_bits_uop_ldst_is_rs1;
      5'b01101:
        casez_tmp_60 = stq_13_bits_uop_ldst_is_rs1;
      5'b01110:
        casez_tmp_60 = stq_14_bits_uop_ldst_is_rs1;
      5'b01111:
        casez_tmp_60 = stq_15_bits_uop_ldst_is_rs1;
      5'b10000:
        casez_tmp_60 = stq_16_bits_uop_ldst_is_rs1;
      5'b10001:
        casez_tmp_60 = stq_17_bits_uop_ldst_is_rs1;
      5'b10010:
        casez_tmp_60 = stq_18_bits_uop_ldst_is_rs1;
      5'b10011:
        casez_tmp_60 = stq_19_bits_uop_ldst_is_rs1;
      5'b10100:
        casez_tmp_60 = stq_20_bits_uop_ldst_is_rs1;
      5'b10101:
        casez_tmp_60 = stq_21_bits_uop_ldst_is_rs1;
      5'b10110:
        casez_tmp_60 = stq_22_bits_uop_ldst_is_rs1;
      5'b10111:
        casez_tmp_60 = stq_23_bits_uop_ldst_is_rs1;
      5'b11000:
        casez_tmp_60 = stq_24_bits_uop_ldst_is_rs1;
      5'b11001:
        casez_tmp_60 = stq_25_bits_uop_ldst_is_rs1;
      5'b11010:
        casez_tmp_60 = stq_26_bits_uop_ldst_is_rs1;
      5'b11011:
        casez_tmp_60 = stq_27_bits_uop_ldst_is_rs1;
      5'b11100:
        casez_tmp_60 = stq_28_bits_uop_ldst_is_rs1;
      5'b11101:
        casez_tmp_60 = stq_29_bits_uop_ldst_is_rs1;
      5'b11110:
        casez_tmp_60 = stq_30_bits_uop_ldst_is_rs1;
      default:
        casez_tmp_60 = stq_31_bits_uop_ldst_is_rs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_61;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_61 = stq_0_bits_uop_ldst;
      5'b00001:
        casez_tmp_61 = stq_1_bits_uop_ldst;
      5'b00010:
        casez_tmp_61 = stq_2_bits_uop_ldst;
      5'b00011:
        casez_tmp_61 = stq_3_bits_uop_ldst;
      5'b00100:
        casez_tmp_61 = stq_4_bits_uop_ldst;
      5'b00101:
        casez_tmp_61 = stq_5_bits_uop_ldst;
      5'b00110:
        casez_tmp_61 = stq_6_bits_uop_ldst;
      5'b00111:
        casez_tmp_61 = stq_7_bits_uop_ldst;
      5'b01000:
        casez_tmp_61 = stq_8_bits_uop_ldst;
      5'b01001:
        casez_tmp_61 = stq_9_bits_uop_ldst;
      5'b01010:
        casez_tmp_61 = stq_10_bits_uop_ldst;
      5'b01011:
        casez_tmp_61 = stq_11_bits_uop_ldst;
      5'b01100:
        casez_tmp_61 = stq_12_bits_uop_ldst;
      5'b01101:
        casez_tmp_61 = stq_13_bits_uop_ldst;
      5'b01110:
        casez_tmp_61 = stq_14_bits_uop_ldst;
      5'b01111:
        casez_tmp_61 = stq_15_bits_uop_ldst;
      5'b10000:
        casez_tmp_61 = stq_16_bits_uop_ldst;
      5'b10001:
        casez_tmp_61 = stq_17_bits_uop_ldst;
      5'b10010:
        casez_tmp_61 = stq_18_bits_uop_ldst;
      5'b10011:
        casez_tmp_61 = stq_19_bits_uop_ldst;
      5'b10100:
        casez_tmp_61 = stq_20_bits_uop_ldst;
      5'b10101:
        casez_tmp_61 = stq_21_bits_uop_ldst;
      5'b10110:
        casez_tmp_61 = stq_22_bits_uop_ldst;
      5'b10111:
        casez_tmp_61 = stq_23_bits_uop_ldst;
      5'b11000:
        casez_tmp_61 = stq_24_bits_uop_ldst;
      5'b11001:
        casez_tmp_61 = stq_25_bits_uop_ldst;
      5'b11010:
        casez_tmp_61 = stq_26_bits_uop_ldst;
      5'b11011:
        casez_tmp_61 = stq_27_bits_uop_ldst;
      5'b11100:
        casez_tmp_61 = stq_28_bits_uop_ldst;
      5'b11101:
        casez_tmp_61 = stq_29_bits_uop_ldst;
      5'b11110:
        casez_tmp_61 = stq_30_bits_uop_ldst;
      default:
        casez_tmp_61 = stq_31_bits_uop_ldst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_62;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_62 = stq_0_bits_uop_lrs1;
      5'b00001:
        casez_tmp_62 = stq_1_bits_uop_lrs1;
      5'b00010:
        casez_tmp_62 = stq_2_bits_uop_lrs1;
      5'b00011:
        casez_tmp_62 = stq_3_bits_uop_lrs1;
      5'b00100:
        casez_tmp_62 = stq_4_bits_uop_lrs1;
      5'b00101:
        casez_tmp_62 = stq_5_bits_uop_lrs1;
      5'b00110:
        casez_tmp_62 = stq_6_bits_uop_lrs1;
      5'b00111:
        casez_tmp_62 = stq_7_bits_uop_lrs1;
      5'b01000:
        casez_tmp_62 = stq_8_bits_uop_lrs1;
      5'b01001:
        casez_tmp_62 = stq_9_bits_uop_lrs1;
      5'b01010:
        casez_tmp_62 = stq_10_bits_uop_lrs1;
      5'b01011:
        casez_tmp_62 = stq_11_bits_uop_lrs1;
      5'b01100:
        casez_tmp_62 = stq_12_bits_uop_lrs1;
      5'b01101:
        casez_tmp_62 = stq_13_bits_uop_lrs1;
      5'b01110:
        casez_tmp_62 = stq_14_bits_uop_lrs1;
      5'b01111:
        casez_tmp_62 = stq_15_bits_uop_lrs1;
      5'b10000:
        casez_tmp_62 = stq_16_bits_uop_lrs1;
      5'b10001:
        casez_tmp_62 = stq_17_bits_uop_lrs1;
      5'b10010:
        casez_tmp_62 = stq_18_bits_uop_lrs1;
      5'b10011:
        casez_tmp_62 = stq_19_bits_uop_lrs1;
      5'b10100:
        casez_tmp_62 = stq_20_bits_uop_lrs1;
      5'b10101:
        casez_tmp_62 = stq_21_bits_uop_lrs1;
      5'b10110:
        casez_tmp_62 = stq_22_bits_uop_lrs1;
      5'b10111:
        casez_tmp_62 = stq_23_bits_uop_lrs1;
      5'b11000:
        casez_tmp_62 = stq_24_bits_uop_lrs1;
      5'b11001:
        casez_tmp_62 = stq_25_bits_uop_lrs1;
      5'b11010:
        casez_tmp_62 = stq_26_bits_uop_lrs1;
      5'b11011:
        casez_tmp_62 = stq_27_bits_uop_lrs1;
      5'b11100:
        casez_tmp_62 = stq_28_bits_uop_lrs1;
      5'b11101:
        casez_tmp_62 = stq_29_bits_uop_lrs1;
      5'b11110:
        casez_tmp_62 = stq_30_bits_uop_lrs1;
      default:
        casez_tmp_62 = stq_31_bits_uop_lrs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_63;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_63 = stq_0_bits_uop_lrs2;
      5'b00001:
        casez_tmp_63 = stq_1_bits_uop_lrs2;
      5'b00010:
        casez_tmp_63 = stq_2_bits_uop_lrs2;
      5'b00011:
        casez_tmp_63 = stq_3_bits_uop_lrs2;
      5'b00100:
        casez_tmp_63 = stq_4_bits_uop_lrs2;
      5'b00101:
        casez_tmp_63 = stq_5_bits_uop_lrs2;
      5'b00110:
        casez_tmp_63 = stq_6_bits_uop_lrs2;
      5'b00111:
        casez_tmp_63 = stq_7_bits_uop_lrs2;
      5'b01000:
        casez_tmp_63 = stq_8_bits_uop_lrs2;
      5'b01001:
        casez_tmp_63 = stq_9_bits_uop_lrs2;
      5'b01010:
        casez_tmp_63 = stq_10_bits_uop_lrs2;
      5'b01011:
        casez_tmp_63 = stq_11_bits_uop_lrs2;
      5'b01100:
        casez_tmp_63 = stq_12_bits_uop_lrs2;
      5'b01101:
        casez_tmp_63 = stq_13_bits_uop_lrs2;
      5'b01110:
        casez_tmp_63 = stq_14_bits_uop_lrs2;
      5'b01111:
        casez_tmp_63 = stq_15_bits_uop_lrs2;
      5'b10000:
        casez_tmp_63 = stq_16_bits_uop_lrs2;
      5'b10001:
        casez_tmp_63 = stq_17_bits_uop_lrs2;
      5'b10010:
        casez_tmp_63 = stq_18_bits_uop_lrs2;
      5'b10011:
        casez_tmp_63 = stq_19_bits_uop_lrs2;
      5'b10100:
        casez_tmp_63 = stq_20_bits_uop_lrs2;
      5'b10101:
        casez_tmp_63 = stq_21_bits_uop_lrs2;
      5'b10110:
        casez_tmp_63 = stq_22_bits_uop_lrs2;
      5'b10111:
        casez_tmp_63 = stq_23_bits_uop_lrs2;
      5'b11000:
        casez_tmp_63 = stq_24_bits_uop_lrs2;
      5'b11001:
        casez_tmp_63 = stq_25_bits_uop_lrs2;
      5'b11010:
        casez_tmp_63 = stq_26_bits_uop_lrs2;
      5'b11011:
        casez_tmp_63 = stq_27_bits_uop_lrs2;
      5'b11100:
        casez_tmp_63 = stq_28_bits_uop_lrs2;
      5'b11101:
        casez_tmp_63 = stq_29_bits_uop_lrs2;
      5'b11110:
        casez_tmp_63 = stq_30_bits_uop_lrs2;
      default:
        casez_tmp_63 = stq_31_bits_uop_lrs2;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_64;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_64 = stq_0_bits_uop_lrs3;
      5'b00001:
        casez_tmp_64 = stq_1_bits_uop_lrs3;
      5'b00010:
        casez_tmp_64 = stq_2_bits_uop_lrs3;
      5'b00011:
        casez_tmp_64 = stq_3_bits_uop_lrs3;
      5'b00100:
        casez_tmp_64 = stq_4_bits_uop_lrs3;
      5'b00101:
        casez_tmp_64 = stq_5_bits_uop_lrs3;
      5'b00110:
        casez_tmp_64 = stq_6_bits_uop_lrs3;
      5'b00111:
        casez_tmp_64 = stq_7_bits_uop_lrs3;
      5'b01000:
        casez_tmp_64 = stq_8_bits_uop_lrs3;
      5'b01001:
        casez_tmp_64 = stq_9_bits_uop_lrs3;
      5'b01010:
        casez_tmp_64 = stq_10_bits_uop_lrs3;
      5'b01011:
        casez_tmp_64 = stq_11_bits_uop_lrs3;
      5'b01100:
        casez_tmp_64 = stq_12_bits_uop_lrs3;
      5'b01101:
        casez_tmp_64 = stq_13_bits_uop_lrs3;
      5'b01110:
        casez_tmp_64 = stq_14_bits_uop_lrs3;
      5'b01111:
        casez_tmp_64 = stq_15_bits_uop_lrs3;
      5'b10000:
        casez_tmp_64 = stq_16_bits_uop_lrs3;
      5'b10001:
        casez_tmp_64 = stq_17_bits_uop_lrs3;
      5'b10010:
        casez_tmp_64 = stq_18_bits_uop_lrs3;
      5'b10011:
        casez_tmp_64 = stq_19_bits_uop_lrs3;
      5'b10100:
        casez_tmp_64 = stq_20_bits_uop_lrs3;
      5'b10101:
        casez_tmp_64 = stq_21_bits_uop_lrs3;
      5'b10110:
        casez_tmp_64 = stq_22_bits_uop_lrs3;
      5'b10111:
        casez_tmp_64 = stq_23_bits_uop_lrs3;
      5'b11000:
        casez_tmp_64 = stq_24_bits_uop_lrs3;
      5'b11001:
        casez_tmp_64 = stq_25_bits_uop_lrs3;
      5'b11010:
        casez_tmp_64 = stq_26_bits_uop_lrs3;
      5'b11011:
        casez_tmp_64 = stq_27_bits_uop_lrs3;
      5'b11100:
        casez_tmp_64 = stq_28_bits_uop_lrs3;
      5'b11101:
        casez_tmp_64 = stq_29_bits_uop_lrs3;
      5'b11110:
        casez_tmp_64 = stq_30_bits_uop_lrs3;
      default:
        casez_tmp_64 = stq_31_bits_uop_lrs3;
    endcase
  end // always @(*)
  reg         casez_tmp_65;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_65 = stq_0_bits_uop_ldst_val;
      5'b00001:
        casez_tmp_65 = stq_1_bits_uop_ldst_val;
      5'b00010:
        casez_tmp_65 = stq_2_bits_uop_ldst_val;
      5'b00011:
        casez_tmp_65 = stq_3_bits_uop_ldst_val;
      5'b00100:
        casez_tmp_65 = stq_4_bits_uop_ldst_val;
      5'b00101:
        casez_tmp_65 = stq_5_bits_uop_ldst_val;
      5'b00110:
        casez_tmp_65 = stq_6_bits_uop_ldst_val;
      5'b00111:
        casez_tmp_65 = stq_7_bits_uop_ldst_val;
      5'b01000:
        casez_tmp_65 = stq_8_bits_uop_ldst_val;
      5'b01001:
        casez_tmp_65 = stq_9_bits_uop_ldst_val;
      5'b01010:
        casez_tmp_65 = stq_10_bits_uop_ldst_val;
      5'b01011:
        casez_tmp_65 = stq_11_bits_uop_ldst_val;
      5'b01100:
        casez_tmp_65 = stq_12_bits_uop_ldst_val;
      5'b01101:
        casez_tmp_65 = stq_13_bits_uop_ldst_val;
      5'b01110:
        casez_tmp_65 = stq_14_bits_uop_ldst_val;
      5'b01111:
        casez_tmp_65 = stq_15_bits_uop_ldst_val;
      5'b10000:
        casez_tmp_65 = stq_16_bits_uop_ldst_val;
      5'b10001:
        casez_tmp_65 = stq_17_bits_uop_ldst_val;
      5'b10010:
        casez_tmp_65 = stq_18_bits_uop_ldst_val;
      5'b10011:
        casez_tmp_65 = stq_19_bits_uop_ldst_val;
      5'b10100:
        casez_tmp_65 = stq_20_bits_uop_ldst_val;
      5'b10101:
        casez_tmp_65 = stq_21_bits_uop_ldst_val;
      5'b10110:
        casez_tmp_65 = stq_22_bits_uop_ldst_val;
      5'b10111:
        casez_tmp_65 = stq_23_bits_uop_ldst_val;
      5'b11000:
        casez_tmp_65 = stq_24_bits_uop_ldst_val;
      5'b11001:
        casez_tmp_65 = stq_25_bits_uop_ldst_val;
      5'b11010:
        casez_tmp_65 = stq_26_bits_uop_ldst_val;
      5'b11011:
        casez_tmp_65 = stq_27_bits_uop_ldst_val;
      5'b11100:
        casez_tmp_65 = stq_28_bits_uop_ldst_val;
      5'b11101:
        casez_tmp_65 = stq_29_bits_uop_ldst_val;
      5'b11110:
        casez_tmp_65 = stq_30_bits_uop_ldst_val;
      default:
        casez_tmp_65 = stq_31_bits_uop_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_66;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_66 = stq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_66 = stq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_66 = stq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_66 = stq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_66 = stq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_66 = stq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_66 = stq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_66 = stq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_66 = stq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_66 = stq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_66 = stq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_66 = stq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_66 = stq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_66 = stq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_66 = stq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_66 = stq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_66 = stq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_66 = stq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_66 = stq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_66 = stq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_66 = stq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_66 = stq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_66 = stq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_66 = stq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_66 = stq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_66 = stq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_66 = stq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_66 = stq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_66 = stq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_66 = stq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_66 = stq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_66 = stq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_67;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_67 = stq_0_bits_uop_lrs1_rtype;
      5'b00001:
        casez_tmp_67 = stq_1_bits_uop_lrs1_rtype;
      5'b00010:
        casez_tmp_67 = stq_2_bits_uop_lrs1_rtype;
      5'b00011:
        casez_tmp_67 = stq_3_bits_uop_lrs1_rtype;
      5'b00100:
        casez_tmp_67 = stq_4_bits_uop_lrs1_rtype;
      5'b00101:
        casez_tmp_67 = stq_5_bits_uop_lrs1_rtype;
      5'b00110:
        casez_tmp_67 = stq_6_bits_uop_lrs1_rtype;
      5'b00111:
        casez_tmp_67 = stq_7_bits_uop_lrs1_rtype;
      5'b01000:
        casez_tmp_67 = stq_8_bits_uop_lrs1_rtype;
      5'b01001:
        casez_tmp_67 = stq_9_bits_uop_lrs1_rtype;
      5'b01010:
        casez_tmp_67 = stq_10_bits_uop_lrs1_rtype;
      5'b01011:
        casez_tmp_67 = stq_11_bits_uop_lrs1_rtype;
      5'b01100:
        casez_tmp_67 = stq_12_bits_uop_lrs1_rtype;
      5'b01101:
        casez_tmp_67 = stq_13_bits_uop_lrs1_rtype;
      5'b01110:
        casez_tmp_67 = stq_14_bits_uop_lrs1_rtype;
      5'b01111:
        casez_tmp_67 = stq_15_bits_uop_lrs1_rtype;
      5'b10000:
        casez_tmp_67 = stq_16_bits_uop_lrs1_rtype;
      5'b10001:
        casez_tmp_67 = stq_17_bits_uop_lrs1_rtype;
      5'b10010:
        casez_tmp_67 = stq_18_bits_uop_lrs1_rtype;
      5'b10011:
        casez_tmp_67 = stq_19_bits_uop_lrs1_rtype;
      5'b10100:
        casez_tmp_67 = stq_20_bits_uop_lrs1_rtype;
      5'b10101:
        casez_tmp_67 = stq_21_bits_uop_lrs1_rtype;
      5'b10110:
        casez_tmp_67 = stq_22_bits_uop_lrs1_rtype;
      5'b10111:
        casez_tmp_67 = stq_23_bits_uop_lrs1_rtype;
      5'b11000:
        casez_tmp_67 = stq_24_bits_uop_lrs1_rtype;
      5'b11001:
        casez_tmp_67 = stq_25_bits_uop_lrs1_rtype;
      5'b11010:
        casez_tmp_67 = stq_26_bits_uop_lrs1_rtype;
      5'b11011:
        casez_tmp_67 = stq_27_bits_uop_lrs1_rtype;
      5'b11100:
        casez_tmp_67 = stq_28_bits_uop_lrs1_rtype;
      5'b11101:
        casez_tmp_67 = stq_29_bits_uop_lrs1_rtype;
      5'b11110:
        casez_tmp_67 = stq_30_bits_uop_lrs1_rtype;
      default:
        casez_tmp_67 = stq_31_bits_uop_lrs1_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_68;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_68 = stq_0_bits_uop_lrs2_rtype;
      5'b00001:
        casez_tmp_68 = stq_1_bits_uop_lrs2_rtype;
      5'b00010:
        casez_tmp_68 = stq_2_bits_uop_lrs2_rtype;
      5'b00011:
        casez_tmp_68 = stq_3_bits_uop_lrs2_rtype;
      5'b00100:
        casez_tmp_68 = stq_4_bits_uop_lrs2_rtype;
      5'b00101:
        casez_tmp_68 = stq_5_bits_uop_lrs2_rtype;
      5'b00110:
        casez_tmp_68 = stq_6_bits_uop_lrs2_rtype;
      5'b00111:
        casez_tmp_68 = stq_7_bits_uop_lrs2_rtype;
      5'b01000:
        casez_tmp_68 = stq_8_bits_uop_lrs2_rtype;
      5'b01001:
        casez_tmp_68 = stq_9_bits_uop_lrs2_rtype;
      5'b01010:
        casez_tmp_68 = stq_10_bits_uop_lrs2_rtype;
      5'b01011:
        casez_tmp_68 = stq_11_bits_uop_lrs2_rtype;
      5'b01100:
        casez_tmp_68 = stq_12_bits_uop_lrs2_rtype;
      5'b01101:
        casez_tmp_68 = stq_13_bits_uop_lrs2_rtype;
      5'b01110:
        casez_tmp_68 = stq_14_bits_uop_lrs2_rtype;
      5'b01111:
        casez_tmp_68 = stq_15_bits_uop_lrs2_rtype;
      5'b10000:
        casez_tmp_68 = stq_16_bits_uop_lrs2_rtype;
      5'b10001:
        casez_tmp_68 = stq_17_bits_uop_lrs2_rtype;
      5'b10010:
        casez_tmp_68 = stq_18_bits_uop_lrs2_rtype;
      5'b10011:
        casez_tmp_68 = stq_19_bits_uop_lrs2_rtype;
      5'b10100:
        casez_tmp_68 = stq_20_bits_uop_lrs2_rtype;
      5'b10101:
        casez_tmp_68 = stq_21_bits_uop_lrs2_rtype;
      5'b10110:
        casez_tmp_68 = stq_22_bits_uop_lrs2_rtype;
      5'b10111:
        casez_tmp_68 = stq_23_bits_uop_lrs2_rtype;
      5'b11000:
        casez_tmp_68 = stq_24_bits_uop_lrs2_rtype;
      5'b11001:
        casez_tmp_68 = stq_25_bits_uop_lrs2_rtype;
      5'b11010:
        casez_tmp_68 = stq_26_bits_uop_lrs2_rtype;
      5'b11011:
        casez_tmp_68 = stq_27_bits_uop_lrs2_rtype;
      5'b11100:
        casez_tmp_68 = stq_28_bits_uop_lrs2_rtype;
      5'b11101:
        casez_tmp_68 = stq_29_bits_uop_lrs2_rtype;
      5'b11110:
        casez_tmp_68 = stq_30_bits_uop_lrs2_rtype;
      default:
        casez_tmp_68 = stq_31_bits_uop_lrs2_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_69;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_69 = stq_0_bits_uop_frs3_en;
      5'b00001:
        casez_tmp_69 = stq_1_bits_uop_frs3_en;
      5'b00010:
        casez_tmp_69 = stq_2_bits_uop_frs3_en;
      5'b00011:
        casez_tmp_69 = stq_3_bits_uop_frs3_en;
      5'b00100:
        casez_tmp_69 = stq_4_bits_uop_frs3_en;
      5'b00101:
        casez_tmp_69 = stq_5_bits_uop_frs3_en;
      5'b00110:
        casez_tmp_69 = stq_6_bits_uop_frs3_en;
      5'b00111:
        casez_tmp_69 = stq_7_bits_uop_frs3_en;
      5'b01000:
        casez_tmp_69 = stq_8_bits_uop_frs3_en;
      5'b01001:
        casez_tmp_69 = stq_9_bits_uop_frs3_en;
      5'b01010:
        casez_tmp_69 = stq_10_bits_uop_frs3_en;
      5'b01011:
        casez_tmp_69 = stq_11_bits_uop_frs3_en;
      5'b01100:
        casez_tmp_69 = stq_12_bits_uop_frs3_en;
      5'b01101:
        casez_tmp_69 = stq_13_bits_uop_frs3_en;
      5'b01110:
        casez_tmp_69 = stq_14_bits_uop_frs3_en;
      5'b01111:
        casez_tmp_69 = stq_15_bits_uop_frs3_en;
      5'b10000:
        casez_tmp_69 = stq_16_bits_uop_frs3_en;
      5'b10001:
        casez_tmp_69 = stq_17_bits_uop_frs3_en;
      5'b10010:
        casez_tmp_69 = stq_18_bits_uop_frs3_en;
      5'b10011:
        casez_tmp_69 = stq_19_bits_uop_frs3_en;
      5'b10100:
        casez_tmp_69 = stq_20_bits_uop_frs3_en;
      5'b10101:
        casez_tmp_69 = stq_21_bits_uop_frs3_en;
      5'b10110:
        casez_tmp_69 = stq_22_bits_uop_frs3_en;
      5'b10111:
        casez_tmp_69 = stq_23_bits_uop_frs3_en;
      5'b11000:
        casez_tmp_69 = stq_24_bits_uop_frs3_en;
      5'b11001:
        casez_tmp_69 = stq_25_bits_uop_frs3_en;
      5'b11010:
        casez_tmp_69 = stq_26_bits_uop_frs3_en;
      5'b11011:
        casez_tmp_69 = stq_27_bits_uop_frs3_en;
      5'b11100:
        casez_tmp_69 = stq_28_bits_uop_frs3_en;
      5'b11101:
        casez_tmp_69 = stq_29_bits_uop_frs3_en;
      5'b11110:
        casez_tmp_69 = stq_30_bits_uop_frs3_en;
      default:
        casez_tmp_69 = stq_31_bits_uop_frs3_en;
    endcase
  end // always @(*)
  reg         casez_tmp_70;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_70 = stq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_70 = stq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_70 = stq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_70 = stq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_70 = stq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_70 = stq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_70 = stq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_70 = stq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_70 = stq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_70 = stq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_70 = stq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_70 = stq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_70 = stq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_70 = stq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_70 = stq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_70 = stq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_70 = stq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_70 = stq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_70 = stq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_70 = stq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_70 = stq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_70 = stq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_70 = stq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_70 = stq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_70 = stq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_70 = stq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_70 = stq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_70 = stq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_70 = stq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_70 = stq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_70 = stq_30_bits_uop_fp_val;
      default:
        casez_tmp_70 = stq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  reg         casez_tmp_71;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_71 = stq_0_bits_uop_fp_single;
      5'b00001:
        casez_tmp_71 = stq_1_bits_uop_fp_single;
      5'b00010:
        casez_tmp_71 = stq_2_bits_uop_fp_single;
      5'b00011:
        casez_tmp_71 = stq_3_bits_uop_fp_single;
      5'b00100:
        casez_tmp_71 = stq_4_bits_uop_fp_single;
      5'b00101:
        casez_tmp_71 = stq_5_bits_uop_fp_single;
      5'b00110:
        casez_tmp_71 = stq_6_bits_uop_fp_single;
      5'b00111:
        casez_tmp_71 = stq_7_bits_uop_fp_single;
      5'b01000:
        casez_tmp_71 = stq_8_bits_uop_fp_single;
      5'b01001:
        casez_tmp_71 = stq_9_bits_uop_fp_single;
      5'b01010:
        casez_tmp_71 = stq_10_bits_uop_fp_single;
      5'b01011:
        casez_tmp_71 = stq_11_bits_uop_fp_single;
      5'b01100:
        casez_tmp_71 = stq_12_bits_uop_fp_single;
      5'b01101:
        casez_tmp_71 = stq_13_bits_uop_fp_single;
      5'b01110:
        casez_tmp_71 = stq_14_bits_uop_fp_single;
      5'b01111:
        casez_tmp_71 = stq_15_bits_uop_fp_single;
      5'b10000:
        casez_tmp_71 = stq_16_bits_uop_fp_single;
      5'b10001:
        casez_tmp_71 = stq_17_bits_uop_fp_single;
      5'b10010:
        casez_tmp_71 = stq_18_bits_uop_fp_single;
      5'b10011:
        casez_tmp_71 = stq_19_bits_uop_fp_single;
      5'b10100:
        casez_tmp_71 = stq_20_bits_uop_fp_single;
      5'b10101:
        casez_tmp_71 = stq_21_bits_uop_fp_single;
      5'b10110:
        casez_tmp_71 = stq_22_bits_uop_fp_single;
      5'b10111:
        casez_tmp_71 = stq_23_bits_uop_fp_single;
      5'b11000:
        casez_tmp_71 = stq_24_bits_uop_fp_single;
      5'b11001:
        casez_tmp_71 = stq_25_bits_uop_fp_single;
      5'b11010:
        casez_tmp_71 = stq_26_bits_uop_fp_single;
      5'b11011:
        casez_tmp_71 = stq_27_bits_uop_fp_single;
      5'b11100:
        casez_tmp_71 = stq_28_bits_uop_fp_single;
      5'b11101:
        casez_tmp_71 = stq_29_bits_uop_fp_single;
      5'b11110:
        casez_tmp_71 = stq_30_bits_uop_fp_single;
      default:
        casez_tmp_71 = stq_31_bits_uop_fp_single;
    endcase
  end // always @(*)
  reg         casez_tmp_72;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_72 = stq_0_bits_uop_xcpt_pf_if;
      5'b00001:
        casez_tmp_72 = stq_1_bits_uop_xcpt_pf_if;
      5'b00010:
        casez_tmp_72 = stq_2_bits_uop_xcpt_pf_if;
      5'b00011:
        casez_tmp_72 = stq_3_bits_uop_xcpt_pf_if;
      5'b00100:
        casez_tmp_72 = stq_4_bits_uop_xcpt_pf_if;
      5'b00101:
        casez_tmp_72 = stq_5_bits_uop_xcpt_pf_if;
      5'b00110:
        casez_tmp_72 = stq_6_bits_uop_xcpt_pf_if;
      5'b00111:
        casez_tmp_72 = stq_7_bits_uop_xcpt_pf_if;
      5'b01000:
        casez_tmp_72 = stq_8_bits_uop_xcpt_pf_if;
      5'b01001:
        casez_tmp_72 = stq_9_bits_uop_xcpt_pf_if;
      5'b01010:
        casez_tmp_72 = stq_10_bits_uop_xcpt_pf_if;
      5'b01011:
        casez_tmp_72 = stq_11_bits_uop_xcpt_pf_if;
      5'b01100:
        casez_tmp_72 = stq_12_bits_uop_xcpt_pf_if;
      5'b01101:
        casez_tmp_72 = stq_13_bits_uop_xcpt_pf_if;
      5'b01110:
        casez_tmp_72 = stq_14_bits_uop_xcpt_pf_if;
      5'b01111:
        casez_tmp_72 = stq_15_bits_uop_xcpt_pf_if;
      5'b10000:
        casez_tmp_72 = stq_16_bits_uop_xcpt_pf_if;
      5'b10001:
        casez_tmp_72 = stq_17_bits_uop_xcpt_pf_if;
      5'b10010:
        casez_tmp_72 = stq_18_bits_uop_xcpt_pf_if;
      5'b10011:
        casez_tmp_72 = stq_19_bits_uop_xcpt_pf_if;
      5'b10100:
        casez_tmp_72 = stq_20_bits_uop_xcpt_pf_if;
      5'b10101:
        casez_tmp_72 = stq_21_bits_uop_xcpt_pf_if;
      5'b10110:
        casez_tmp_72 = stq_22_bits_uop_xcpt_pf_if;
      5'b10111:
        casez_tmp_72 = stq_23_bits_uop_xcpt_pf_if;
      5'b11000:
        casez_tmp_72 = stq_24_bits_uop_xcpt_pf_if;
      5'b11001:
        casez_tmp_72 = stq_25_bits_uop_xcpt_pf_if;
      5'b11010:
        casez_tmp_72 = stq_26_bits_uop_xcpt_pf_if;
      5'b11011:
        casez_tmp_72 = stq_27_bits_uop_xcpt_pf_if;
      5'b11100:
        casez_tmp_72 = stq_28_bits_uop_xcpt_pf_if;
      5'b11101:
        casez_tmp_72 = stq_29_bits_uop_xcpt_pf_if;
      5'b11110:
        casez_tmp_72 = stq_30_bits_uop_xcpt_pf_if;
      default:
        casez_tmp_72 = stq_31_bits_uop_xcpt_pf_if;
    endcase
  end // always @(*)
  reg         casez_tmp_73;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_73 = stq_0_bits_uop_xcpt_ae_if;
      5'b00001:
        casez_tmp_73 = stq_1_bits_uop_xcpt_ae_if;
      5'b00010:
        casez_tmp_73 = stq_2_bits_uop_xcpt_ae_if;
      5'b00011:
        casez_tmp_73 = stq_3_bits_uop_xcpt_ae_if;
      5'b00100:
        casez_tmp_73 = stq_4_bits_uop_xcpt_ae_if;
      5'b00101:
        casez_tmp_73 = stq_5_bits_uop_xcpt_ae_if;
      5'b00110:
        casez_tmp_73 = stq_6_bits_uop_xcpt_ae_if;
      5'b00111:
        casez_tmp_73 = stq_7_bits_uop_xcpt_ae_if;
      5'b01000:
        casez_tmp_73 = stq_8_bits_uop_xcpt_ae_if;
      5'b01001:
        casez_tmp_73 = stq_9_bits_uop_xcpt_ae_if;
      5'b01010:
        casez_tmp_73 = stq_10_bits_uop_xcpt_ae_if;
      5'b01011:
        casez_tmp_73 = stq_11_bits_uop_xcpt_ae_if;
      5'b01100:
        casez_tmp_73 = stq_12_bits_uop_xcpt_ae_if;
      5'b01101:
        casez_tmp_73 = stq_13_bits_uop_xcpt_ae_if;
      5'b01110:
        casez_tmp_73 = stq_14_bits_uop_xcpt_ae_if;
      5'b01111:
        casez_tmp_73 = stq_15_bits_uop_xcpt_ae_if;
      5'b10000:
        casez_tmp_73 = stq_16_bits_uop_xcpt_ae_if;
      5'b10001:
        casez_tmp_73 = stq_17_bits_uop_xcpt_ae_if;
      5'b10010:
        casez_tmp_73 = stq_18_bits_uop_xcpt_ae_if;
      5'b10011:
        casez_tmp_73 = stq_19_bits_uop_xcpt_ae_if;
      5'b10100:
        casez_tmp_73 = stq_20_bits_uop_xcpt_ae_if;
      5'b10101:
        casez_tmp_73 = stq_21_bits_uop_xcpt_ae_if;
      5'b10110:
        casez_tmp_73 = stq_22_bits_uop_xcpt_ae_if;
      5'b10111:
        casez_tmp_73 = stq_23_bits_uop_xcpt_ae_if;
      5'b11000:
        casez_tmp_73 = stq_24_bits_uop_xcpt_ae_if;
      5'b11001:
        casez_tmp_73 = stq_25_bits_uop_xcpt_ae_if;
      5'b11010:
        casez_tmp_73 = stq_26_bits_uop_xcpt_ae_if;
      5'b11011:
        casez_tmp_73 = stq_27_bits_uop_xcpt_ae_if;
      5'b11100:
        casez_tmp_73 = stq_28_bits_uop_xcpt_ae_if;
      5'b11101:
        casez_tmp_73 = stq_29_bits_uop_xcpt_ae_if;
      5'b11110:
        casez_tmp_73 = stq_30_bits_uop_xcpt_ae_if;
      default:
        casez_tmp_73 = stq_31_bits_uop_xcpt_ae_if;
    endcase
  end // always @(*)
  reg         casez_tmp_74;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_74 = stq_0_bits_uop_xcpt_ma_if;
      5'b00001:
        casez_tmp_74 = stq_1_bits_uop_xcpt_ma_if;
      5'b00010:
        casez_tmp_74 = stq_2_bits_uop_xcpt_ma_if;
      5'b00011:
        casez_tmp_74 = stq_3_bits_uop_xcpt_ma_if;
      5'b00100:
        casez_tmp_74 = stq_4_bits_uop_xcpt_ma_if;
      5'b00101:
        casez_tmp_74 = stq_5_bits_uop_xcpt_ma_if;
      5'b00110:
        casez_tmp_74 = stq_6_bits_uop_xcpt_ma_if;
      5'b00111:
        casez_tmp_74 = stq_7_bits_uop_xcpt_ma_if;
      5'b01000:
        casez_tmp_74 = stq_8_bits_uop_xcpt_ma_if;
      5'b01001:
        casez_tmp_74 = stq_9_bits_uop_xcpt_ma_if;
      5'b01010:
        casez_tmp_74 = stq_10_bits_uop_xcpt_ma_if;
      5'b01011:
        casez_tmp_74 = stq_11_bits_uop_xcpt_ma_if;
      5'b01100:
        casez_tmp_74 = stq_12_bits_uop_xcpt_ma_if;
      5'b01101:
        casez_tmp_74 = stq_13_bits_uop_xcpt_ma_if;
      5'b01110:
        casez_tmp_74 = stq_14_bits_uop_xcpt_ma_if;
      5'b01111:
        casez_tmp_74 = stq_15_bits_uop_xcpt_ma_if;
      5'b10000:
        casez_tmp_74 = stq_16_bits_uop_xcpt_ma_if;
      5'b10001:
        casez_tmp_74 = stq_17_bits_uop_xcpt_ma_if;
      5'b10010:
        casez_tmp_74 = stq_18_bits_uop_xcpt_ma_if;
      5'b10011:
        casez_tmp_74 = stq_19_bits_uop_xcpt_ma_if;
      5'b10100:
        casez_tmp_74 = stq_20_bits_uop_xcpt_ma_if;
      5'b10101:
        casez_tmp_74 = stq_21_bits_uop_xcpt_ma_if;
      5'b10110:
        casez_tmp_74 = stq_22_bits_uop_xcpt_ma_if;
      5'b10111:
        casez_tmp_74 = stq_23_bits_uop_xcpt_ma_if;
      5'b11000:
        casez_tmp_74 = stq_24_bits_uop_xcpt_ma_if;
      5'b11001:
        casez_tmp_74 = stq_25_bits_uop_xcpt_ma_if;
      5'b11010:
        casez_tmp_74 = stq_26_bits_uop_xcpt_ma_if;
      5'b11011:
        casez_tmp_74 = stq_27_bits_uop_xcpt_ma_if;
      5'b11100:
        casez_tmp_74 = stq_28_bits_uop_xcpt_ma_if;
      5'b11101:
        casez_tmp_74 = stq_29_bits_uop_xcpt_ma_if;
      5'b11110:
        casez_tmp_74 = stq_30_bits_uop_xcpt_ma_if;
      default:
        casez_tmp_74 = stq_31_bits_uop_xcpt_ma_if;
    endcase
  end // always @(*)
  reg         casez_tmp_75;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_75 = stq_0_bits_uop_bp_debug_if;
      5'b00001:
        casez_tmp_75 = stq_1_bits_uop_bp_debug_if;
      5'b00010:
        casez_tmp_75 = stq_2_bits_uop_bp_debug_if;
      5'b00011:
        casez_tmp_75 = stq_3_bits_uop_bp_debug_if;
      5'b00100:
        casez_tmp_75 = stq_4_bits_uop_bp_debug_if;
      5'b00101:
        casez_tmp_75 = stq_5_bits_uop_bp_debug_if;
      5'b00110:
        casez_tmp_75 = stq_6_bits_uop_bp_debug_if;
      5'b00111:
        casez_tmp_75 = stq_7_bits_uop_bp_debug_if;
      5'b01000:
        casez_tmp_75 = stq_8_bits_uop_bp_debug_if;
      5'b01001:
        casez_tmp_75 = stq_9_bits_uop_bp_debug_if;
      5'b01010:
        casez_tmp_75 = stq_10_bits_uop_bp_debug_if;
      5'b01011:
        casez_tmp_75 = stq_11_bits_uop_bp_debug_if;
      5'b01100:
        casez_tmp_75 = stq_12_bits_uop_bp_debug_if;
      5'b01101:
        casez_tmp_75 = stq_13_bits_uop_bp_debug_if;
      5'b01110:
        casez_tmp_75 = stq_14_bits_uop_bp_debug_if;
      5'b01111:
        casez_tmp_75 = stq_15_bits_uop_bp_debug_if;
      5'b10000:
        casez_tmp_75 = stq_16_bits_uop_bp_debug_if;
      5'b10001:
        casez_tmp_75 = stq_17_bits_uop_bp_debug_if;
      5'b10010:
        casez_tmp_75 = stq_18_bits_uop_bp_debug_if;
      5'b10011:
        casez_tmp_75 = stq_19_bits_uop_bp_debug_if;
      5'b10100:
        casez_tmp_75 = stq_20_bits_uop_bp_debug_if;
      5'b10101:
        casez_tmp_75 = stq_21_bits_uop_bp_debug_if;
      5'b10110:
        casez_tmp_75 = stq_22_bits_uop_bp_debug_if;
      5'b10111:
        casez_tmp_75 = stq_23_bits_uop_bp_debug_if;
      5'b11000:
        casez_tmp_75 = stq_24_bits_uop_bp_debug_if;
      5'b11001:
        casez_tmp_75 = stq_25_bits_uop_bp_debug_if;
      5'b11010:
        casez_tmp_75 = stq_26_bits_uop_bp_debug_if;
      5'b11011:
        casez_tmp_75 = stq_27_bits_uop_bp_debug_if;
      5'b11100:
        casez_tmp_75 = stq_28_bits_uop_bp_debug_if;
      5'b11101:
        casez_tmp_75 = stq_29_bits_uop_bp_debug_if;
      5'b11110:
        casez_tmp_75 = stq_30_bits_uop_bp_debug_if;
      default:
        casez_tmp_75 = stq_31_bits_uop_bp_debug_if;
    endcase
  end // always @(*)
  reg         casez_tmp_76;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_76 = stq_0_bits_uop_bp_xcpt_if;
      5'b00001:
        casez_tmp_76 = stq_1_bits_uop_bp_xcpt_if;
      5'b00010:
        casez_tmp_76 = stq_2_bits_uop_bp_xcpt_if;
      5'b00011:
        casez_tmp_76 = stq_3_bits_uop_bp_xcpt_if;
      5'b00100:
        casez_tmp_76 = stq_4_bits_uop_bp_xcpt_if;
      5'b00101:
        casez_tmp_76 = stq_5_bits_uop_bp_xcpt_if;
      5'b00110:
        casez_tmp_76 = stq_6_bits_uop_bp_xcpt_if;
      5'b00111:
        casez_tmp_76 = stq_7_bits_uop_bp_xcpt_if;
      5'b01000:
        casez_tmp_76 = stq_8_bits_uop_bp_xcpt_if;
      5'b01001:
        casez_tmp_76 = stq_9_bits_uop_bp_xcpt_if;
      5'b01010:
        casez_tmp_76 = stq_10_bits_uop_bp_xcpt_if;
      5'b01011:
        casez_tmp_76 = stq_11_bits_uop_bp_xcpt_if;
      5'b01100:
        casez_tmp_76 = stq_12_bits_uop_bp_xcpt_if;
      5'b01101:
        casez_tmp_76 = stq_13_bits_uop_bp_xcpt_if;
      5'b01110:
        casez_tmp_76 = stq_14_bits_uop_bp_xcpt_if;
      5'b01111:
        casez_tmp_76 = stq_15_bits_uop_bp_xcpt_if;
      5'b10000:
        casez_tmp_76 = stq_16_bits_uop_bp_xcpt_if;
      5'b10001:
        casez_tmp_76 = stq_17_bits_uop_bp_xcpt_if;
      5'b10010:
        casez_tmp_76 = stq_18_bits_uop_bp_xcpt_if;
      5'b10011:
        casez_tmp_76 = stq_19_bits_uop_bp_xcpt_if;
      5'b10100:
        casez_tmp_76 = stq_20_bits_uop_bp_xcpt_if;
      5'b10101:
        casez_tmp_76 = stq_21_bits_uop_bp_xcpt_if;
      5'b10110:
        casez_tmp_76 = stq_22_bits_uop_bp_xcpt_if;
      5'b10111:
        casez_tmp_76 = stq_23_bits_uop_bp_xcpt_if;
      5'b11000:
        casez_tmp_76 = stq_24_bits_uop_bp_xcpt_if;
      5'b11001:
        casez_tmp_76 = stq_25_bits_uop_bp_xcpt_if;
      5'b11010:
        casez_tmp_76 = stq_26_bits_uop_bp_xcpt_if;
      5'b11011:
        casez_tmp_76 = stq_27_bits_uop_bp_xcpt_if;
      5'b11100:
        casez_tmp_76 = stq_28_bits_uop_bp_xcpt_if;
      5'b11101:
        casez_tmp_76 = stq_29_bits_uop_bp_xcpt_if;
      5'b11110:
        casez_tmp_76 = stq_30_bits_uop_bp_xcpt_if;
      default:
        casez_tmp_76 = stq_31_bits_uop_bp_xcpt_if;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_77;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_77 = stq_0_bits_uop_debug_fsrc;
      5'b00001:
        casez_tmp_77 = stq_1_bits_uop_debug_fsrc;
      5'b00010:
        casez_tmp_77 = stq_2_bits_uop_debug_fsrc;
      5'b00011:
        casez_tmp_77 = stq_3_bits_uop_debug_fsrc;
      5'b00100:
        casez_tmp_77 = stq_4_bits_uop_debug_fsrc;
      5'b00101:
        casez_tmp_77 = stq_5_bits_uop_debug_fsrc;
      5'b00110:
        casez_tmp_77 = stq_6_bits_uop_debug_fsrc;
      5'b00111:
        casez_tmp_77 = stq_7_bits_uop_debug_fsrc;
      5'b01000:
        casez_tmp_77 = stq_8_bits_uop_debug_fsrc;
      5'b01001:
        casez_tmp_77 = stq_9_bits_uop_debug_fsrc;
      5'b01010:
        casez_tmp_77 = stq_10_bits_uop_debug_fsrc;
      5'b01011:
        casez_tmp_77 = stq_11_bits_uop_debug_fsrc;
      5'b01100:
        casez_tmp_77 = stq_12_bits_uop_debug_fsrc;
      5'b01101:
        casez_tmp_77 = stq_13_bits_uop_debug_fsrc;
      5'b01110:
        casez_tmp_77 = stq_14_bits_uop_debug_fsrc;
      5'b01111:
        casez_tmp_77 = stq_15_bits_uop_debug_fsrc;
      5'b10000:
        casez_tmp_77 = stq_16_bits_uop_debug_fsrc;
      5'b10001:
        casez_tmp_77 = stq_17_bits_uop_debug_fsrc;
      5'b10010:
        casez_tmp_77 = stq_18_bits_uop_debug_fsrc;
      5'b10011:
        casez_tmp_77 = stq_19_bits_uop_debug_fsrc;
      5'b10100:
        casez_tmp_77 = stq_20_bits_uop_debug_fsrc;
      5'b10101:
        casez_tmp_77 = stq_21_bits_uop_debug_fsrc;
      5'b10110:
        casez_tmp_77 = stq_22_bits_uop_debug_fsrc;
      5'b10111:
        casez_tmp_77 = stq_23_bits_uop_debug_fsrc;
      5'b11000:
        casez_tmp_77 = stq_24_bits_uop_debug_fsrc;
      5'b11001:
        casez_tmp_77 = stq_25_bits_uop_debug_fsrc;
      5'b11010:
        casez_tmp_77 = stq_26_bits_uop_debug_fsrc;
      5'b11011:
        casez_tmp_77 = stq_27_bits_uop_debug_fsrc;
      5'b11100:
        casez_tmp_77 = stq_28_bits_uop_debug_fsrc;
      5'b11101:
        casez_tmp_77 = stq_29_bits_uop_debug_fsrc;
      5'b11110:
        casez_tmp_77 = stq_30_bits_uop_debug_fsrc;
      default:
        casez_tmp_77 = stq_31_bits_uop_debug_fsrc;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_78;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_78 = stq_0_bits_uop_debug_tsrc;
      5'b00001:
        casez_tmp_78 = stq_1_bits_uop_debug_tsrc;
      5'b00010:
        casez_tmp_78 = stq_2_bits_uop_debug_tsrc;
      5'b00011:
        casez_tmp_78 = stq_3_bits_uop_debug_tsrc;
      5'b00100:
        casez_tmp_78 = stq_4_bits_uop_debug_tsrc;
      5'b00101:
        casez_tmp_78 = stq_5_bits_uop_debug_tsrc;
      5'b00110:
        casez_tmp_78 = stq_6_bits_uop_debug_tsrc;
      5'b00111:
        casez_tmp_78 = stq_7_bits_uop_debug_tsrc;
      5'b01000:
        casez_tmp_78 = stq_8_bits_uop_debug_tsrc;
      5'b01001:
        casez_tmp_78 = stq_9_bits_uop_debug_tsrc;
      5'b01010:
        casez_tmp_78 = stq_10_bits_uop_debug_tsrc;
      5'b01011:
        casez_tmp_78 = stq_11_bits_uop_debug_tsrc;
      5'b01100:
        casez_tmp_78 = stq_12_bits_uop_debug_tsrc;
      5'b01101:
        casez_tmp_78 = stq_13_bits_uop_debug_tsrc;
      5'b01110:
        casez_tmp_78 = stq_14_bits_uop_debug_tsrc;
      5'b01111:
        casez_tmp_78 = stq_15_bits_uop_debug_tsrc;
      5'b10000:
        casez_tmp_78 = stq_16_bits_uop_debug_tsrc;
      5'b10001:
        casez_tmp_78 = stq_17_bits_uop_debug_tsrc;
      5'b10010:
        casez_tmp_78 = stq_18_bits_uop_debug_tsrc;
      5'b10011:
        casez_tmp_78 = stq_19_bits_uop_debug_tsrc;
      5'b10100:
        casez_tmp_78 = stq_20_bits_uop_debug_tsrc;
      5'b10101:
        casez_tmp_78 = stq_21_bits_uop_debug_tsrc;
      5'b10110:
        casez_tmp_78 = stq_22_bits_uop_debug_tsrc;
      5'b10111:
        casez_tmp_78 = stq_23_bits_uop_debug_tsrc;
      5'b11000:
        casez_tmp_78 = stq_24_bits_uop_debug_tsrc;
      5'b11001:
        casez_tmp_78 = stq_25_bits_uop_debug_tsrc;
      5'b11010:
        casez_tmp_78 = stq_26_bits_uop_debug_tsrc;
      5'b11011:
        casez_tmp_78 = stq_27_bits_uop_debug_tsrc;
      5'b11100:
        casez_tmp_78 = stq_28_bits_uop_debug_tsrc;
      5'b11101:
        casez_tmp_78 = stq_29_bits_uop_debug_tsrc;
      5'b11110:
        casez_tmp_78 = stq_30_bits_uop_debug_tsrc;
      default:
        casez_tmp_78 = stq_31_bits_uop_debug_tsrc;
    endcase
  end // always @(*)
  reg         casez_tmp_79;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_79 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_79 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_79 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_79 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_79 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_79 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_79 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_79 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_79 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_79 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_79 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_79 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_79 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_79 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_79 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_79 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_79 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_79 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_79 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_79 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_79 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_79 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_79 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_79 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_79 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_79 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_79 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_79 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_79 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_79 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_79 = stq_30_bits_addr_valid;
      default:
        casez_tmp_79 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_80;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_80 = stq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_80 = stq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_80 = stq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_80 = stq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_80 = stq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_80 = stq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_80 = stq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_80 = stq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_80 = stq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_80 = stq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_80 = stq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_80 = stq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_80 = stq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_80 = stq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_80 = stq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_80 = stq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_80 = stq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_80 = stq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_80 = stq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_80 = stq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_80 = stq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_80 = stq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_80 = stq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_80 = stq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_80 = stq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_80 = stq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_80 = stq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_80 = stq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_80 = stq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_80 = stq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_80 = stq_30_bits_addr_bits;
      default:
        casez_tmp_80 = stq_31_bits_addr_bits;
    endcase
  end // always @(*)
  reg         casez_tmp_81;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_81 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_81 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_81 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_81 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_81 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_81 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_81 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_81 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_81 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_81 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_81 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_81 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_81 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_81 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_81 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_81 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_81 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_81 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_81 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_81 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_81 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_81 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_81 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_81 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_81 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_81 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_81 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_81 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_81 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_81 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_81 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_81 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         casez_tmp_82;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_82 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_82 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_82 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_82 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_82 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_82 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_82 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_82 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_82 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_82 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_82 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_82 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_82 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_82 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_82 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_82 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_82 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_82 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_82 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_82 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_82 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_82 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_82 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_82 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_82 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_82 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_82 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_82 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_82 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_82 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_82 = stq_30_bits_data_valid;
      default:
        casez_tmp_82 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_83;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_83 = stq_0_bits_data_bits;
      5'b00001:
        casez_tmp_83 = stq_1_bits_data_bits;
      5'b00010:
        casez_tmp_83 = stq_2_bits_data_bits;
      5'b00011:
        casez_tmp_83 = stq_3_bits_data_bits;
      5'b00100:
        casez_tmp_83 = stq_4_bits_data_bits;
      5'b00101:
        casez_tmp_83 = stq_5_bits_data_bits;
      5'b00110:
        casez_tmp_83 = stq_6_bits_data_bits;
      5'b00111:
        casez_tmp_83 = stq_7_bits_data_bits;
      5'b01000:
        casez_tmp_83 = stq_8_bits_data_bits;
      5'b01001:
        casez_tmp_83 = stq_9_bits_data_bits;
      5'b01010:
        casez_tmp_83 = stq_10_bits_data_bits;
      5'b01011:
        casez_tmp_83 = stq_11_bits_data_bits;
      5'b01100:
        casez_tmp_83 = stq_12_bits_data_bits;
      5'b01101:
        casez_tmp_83 = stq_13_bits_data_bits;
      5'b01110:
        casez_tmp_83 = stq_14_bits_data_bits;
      5'b01111:
        casez_tmp_83 = stq_15_bits_data_bits;
      5'b10000:
        casez_tmp_83 = stq_16_bits_data_bits;
      5'b10001:
        casez_tmp_83 = stq_17_bits_data_bits;
      5'b10010:
        casez_tmp_83 = stq_18_bits_data_bits;
      5'b10011:
        casez_tmp_83 = stq_19_bits_data_bits;
      5'b10100:
        casez_tmp_83 = stq_20_bits_data_bits;
      5'b10101:
        casez_tmp_83 = stq_21_bits_data_bits;
      5'b10110:
        casez_tmp_83 = stq_22_bits_data_bits;
      5'b10111:
        casez_tmp_83 = stq_23_bits_data_bits;
      5'b11000:
        casez_tmp_83 = stq_24_bits_data_bits;
      5'b11001:
        casez_tmp_83 = stq_25_bits_data_bits;
      5'b11010:
        casez_tmp_83 = stq_26_bits_data_bits;
      5'b11011:
        casez_tmp_83 = stq_27_bits_data_bits;
      5'b11100:
        casez_tmp_83 = stq_28_bits_data_bits;
      5'b11101:
        casez_tmp_83 = stq_29_bits_data_bits;
      5'b11110:
        casez_tmp_83 = stq_30_bits_data_bits;
      default:
        casez_tmp_83 = stq_31_bits_data_bits;
    endcase
  end // always @(*)
  reg         casez_tmp_84;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_84 = stq_0_bits_committed;
      5'b00001:
        casez_tmp_84 = stq_1_bits_committed;
      5'b00010:
        casez_tmp_84 = stq_2_bits_committed;
      5'b00011:
        casez_tmp_84 = stq_3_bits_committed;
      5'b00100:
        casez_tmp_84 = stq_4_bits_committed;
      5'b00101:
        casez_tmp_84 = stq_5_bits_committed;
      5'b00110:
        casez_tmp_84 = stq_6_bits_committed;
      5'b00111:
        casez_tmp_84 = stq_7_bits_committed;
      5'b01000:
        casez_tmp_84 = stq_8_bits_committed;
      5'b01001:
        casez_tmp_84 = stq_9_bits_committed;
      5'b01010:
        casez_tmp_84 = stq_10_bits_committed;
      5'b01011:
        casez_tmp_84 = stq_11_bits_committed;
      5'b01100:
        casez_tmp_84 = stq_12_bits_committed;
      5'b01101:
        casez_tmp_84 = stq_13_bits_committed;
      5'b01110:
        casez_tmp_84 = stq_14_bits_committed;
      5'b01111:
        casez_tmp_84 = stq_15_bits_committed;
      5'b10000:
        casez_tmp_84 = stq_16_bits_committed;
      5'b10001:
        casez_tmp_84 = stq_17_bits_committed;
      5'b10010:
        casez_tmp_84 = stq_18_bits_committed;
      5'b10011:
        casez_tmp_84 = stq_19_bits_committed;
      5'b10100:
        casez_tmp_84 = stq_20_bits_committed;
      5'b10101:
        casez_tmp_84 = stq_21_bits_committed;
      5'b10110:
        casez_tmp_84 = stq_22_bits_committed;
      5'b10111:
        casez_tmp_84 = stq_23_bits_committed;
      5'b11000:
        casez_tmp_84 = stq_24_bits_committed;
      5'b11001:
        casez_tmp_84 = stq_25_bits_committed;
      5'b11010:
        casez_tmp_84 = stq_26_bits_committed;
      5'b11011:
        casez_tmp_84 = stq_27_bits_committed;
      5'b11100:
        casez_tmp_84 = stq_28_bits_committed;
      5'b11101:
        casez_tmp_84 = stq_29_bits_committed;
      5'b11110:
        casez_tmp_84 = stq_30_bits_committed;
      default:
        casez_tmp_84 = stq_31_bits_committed;
    endcase
  end // always @(*)
  reg  [2:0]  hella_state;
  reg  [39:0] hella_req_addr;
  reg  [63:0] hella_data_data;
  reg  [32:0] hella_paddr;
  reg         hella_xcpt_ma_ld;
  reg         hella_xcpt_ma_st;
  reg         hella_xcpt_pf_ld;
  reg         hella_xcpt_pf_st;
  reg         hella_xcpt_gf_ld;
  reg         hella_xcpt_gf_st;
  reg         hella_xcpt_ae_ld;
  reg         hella_xcpt_ae_st;
  reg  [31:0] live_store_mask;
  wire [4:0]  _GEN_3 = ldq_tail + 5'h1;
  wire [4:0]  _GEN_4 = stq_tail + 5'h1;
  wire        dis_ld_val = io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_ldq & ~io_core_dis_uops_0_bits_exception;
  wire        dis_st_val = io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_stq & ~io_core_dis_uops_0_bits_exception;
  reg         casez_tmp_85;
  always @(*) begin
    casez (ldq_tail)
      5'b00000:
        casez_tmp_85 = ldq_0_valid;
      5'b00001:
        casez_tmp_85 = ldq_1_valid;
      5'b00010:
        casez_tmp_85 = ldq_2_valid;
      5'b00011:
        casez_tmp_85 = ldq_3_valid;
      5'b00100:
        casez_tmp_85 = ldq_4_valid;
      5'b00101:
        casez_tmp_85 = ldq_5_valid;
      5'b00110:
        casez_tmp_85 = ldq_6_valid;
      5'b00111:
        casez_tmp_85 = ldq_7_valid;
      5'b01000:
        casez_tmp_85 = ldq_8_valid;
      5'b01001:
        casez_tmp_85 = ldq_9_valid;
      5'b01010:
        casez_tmp_85 = ldq_10_valid;
      5'b01011:
        casez_tmp_85 = ldq_11_valid;
      5'b01100:
        casez_tmp_85 = ldq_12_valid;
      5'b01101:
        casez_tmp_85 = ldq_13_valid;
      5'b01110:
        casez_tmp_85 = ldq_14_valid;
      5'b01111:
        casez_tmp_85 = ldq_15_valid;
      5'b10000:
        casez_tmp_85 = ldq_16_valid;
      5'b10001:
        casez_tmp_85 = ldq_17_valid;
      5'b10010:
        casez_tmp_85 = ldq_18_valid;
      5'b10011:
        casez_tmp_85 = ldq_19_valid;
      5'b10100:
        casez_tmp_85 = ldq_20_valid;
      5'b10101:
        casez_tmp_85 = ldq_21_valid;
      5'b10110:
        casez_tmp_85 = ldq_22_valid;
      5'b10111:
        casez_tmp_85 = ldq_23_valid;
      5'b11000:
        casez_tmp_85 = ldq_24_valid;
      5'b11001:
        casez_tmp_85 = ldq_25_valid;
      5'b11010:
        casez_tmp_85 = ldq_26_valid;
      5'b11011:
        casez_tmp_85 = ldq_27_valid;
      5'b11100:
        casez_tmp_85 = ldq_28_valid;
      5'b11101:
        casez_tmp_85 = ldq_29_valid;
      5'b11110:
        casez_tmp_85 = ldq_30_valid;
      default:
        casez_tmp_85 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_86;
  always @(*) begin
    casez (stq_tail)
      5'b00000:
        casez_tmp_86 = stq_0_valid;
      5'b00001:
        casez_tmp_86 = stq_1_valid;
      5'b00010:
        casez_tmp_86 = stq_2_valid;
      5'b00011:
        casez_tmp_86 = stq_3_valid;
      5'b00100:
        casez_tmp_86 = stq_4_valid;
      5'b00101:
        casez_tmp_86 = stq_5_valid;
      5'b00110:
        casez_tmp_86 = stq_6_valid;
      5'b00111:
        casez_tmp_86 = stq_7_valid;
      5'b01000:
        casez_tmp_86 = stq_8_valid;
      5'b01001:
        casez_tmp_86 = stq_9_valid;
      5'b01010:
        casez_tmp_86 = stq_10_valid;
      5'b01011:
        casez_tmp_86 = stq_11_valid;
      5'b01100:
        casez_tmp_86 = stq_12_valid;
      5'b01101:
        casez_tmp_86 = stq_13_valid;
      5'b01110:
        casez_tmp_86 = stq_14_valid;
      5'b01111:
        casez_tmp_86 = stq_15_valid;
      5'b10000:
        casez_tmp_86 = stq_16_valid;
      5'b10001:
        casez_tmp_86 = stq_17_valid;
      5'b10010:
        casez_tmp_86 = stq_18_valid;
      5'b10011:
        casez_tmp_86 = stq_19_valid;
      5'b10100:
        casez_tmp_86 = stq_20_valid;
      5'b10101:
        casez_tmp_86 = stq_21_valid;
      5'b10110:
        casez_tmp_86 = stq_22_valid;
      5'b10111:
        casez_tmp_86 = stq_23_valid;
      5'b11000:
        casez_tmp_86 = stq_24_valid;
      5'b11001:
        casez_tmp_86 = stq_25_valid;
      5'b11010:
        casez_tmp_86 = stq_26_valid;
      5'b11011:
        casez_tmp_86 = stq_27_valid;
      5'b11100:
        casez_tmp_86 = stq_28_valid;
      5'b11101:
        casez_tmp_86 = stq_29_valid;
      5'b11110:
        casez_tmp_86 = stq_30_valid;
      default:
        casez_tmp_86 = stq_31_valid;
    endcase
  end // always @(*)
  wire [4:0]  _GEN_5 = dis_ld_val ? _GEN_3 : ldq_tail;
  wire [4:0]  _GEN_6 = dis_st_val ? _GEN_4 : stq_tail;
  wire [4:0]  _GEN_7 = _GEN_5 + 5'h1;
  wire [4:0]  _GEN_8 = _GEN_6 + 5'h1;
  wire        dis_ld_val_1 = io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_ldq & ~io_core_dis_uops_1_bits_exception;
  wire        dis_st_val_1 = io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_stq & ~io_core_dis_uops_1_bits_exception;
  reg         casez_tmp_87;
  always @(*) begin
    casez (_GEN_5)
      5'b00000:
        casez_tmp_87 = ldq_0_valid;
      5'b00001:
        casez_tmp_87 = ldq_1_valid;
      5'b00010:
        casez_tmp_87 = ldq_2_valid;
      5'b00011:
        casez_tmp_87 = ldq_3_valid;
      5'b00100:
        casez_tmp_87 = ldq_4_valid;
      5'b00101:
        casez_tmp_87 = ldq_5_valid;
      5'b00110:
        casez_tmp_87 = ldq_6_valid;
      5'b00111:
        casez_tmp_87 = ldq_7_valid;
      5'b01000:
        casez_tmp_87 = ldq_8_valid;
      5'b01001:
        casez_tmp_87 = ldq_9_valid;
      5'b01010:
        casez_tmp_87 = ldq_10_valid;
      5'b01011:
        casez_tmp_87 = ldq_11_valid;
      5'b01100:
        casez_tmp_87 = ldq_12_valid;
      5'b01101:
        casez_tmp_87 = ldq_13_valid;
      5'b01110:
        casez_tmp_87 = ldq_14_valid;
      5'b01111:
        casez_tmp_87 = ldq_15_valid;
      5'b10000:
        casez_tmp_87 = ldq_16_valid;
      5'b10001:
        casez_tmp_87 = ldq_17_valid;
      5'b10010:
        casez_tmp_87 = ldq_18_valid;
      5'b10011:
        casez_tmp_87 = ldq_19_valid;
      5'b10100:
        casez_tmp_87 = ldq_20_valid;
      5'b10101:
        casez_tmp_87 = ldq_21_valid;
      5'b10110:
        casez_tmp_87 = ldq_22_valid;
      5'b10111:
        casez_tmp_87 = ldq_23_valid;
      5'b11000:
        casez_tmp_87 = ldq_24_valid;
      5'b11001:
        casez_tmp_87 = ldq_25_valid;
      5'b11010:
        casez_tmp_87 = ldq_26_valid;
      5'b11011:
        casez_tmp_87 = ldq_27_valid;
      5'b11100:
        casez_tmp_87 = ldq_28_valid;
      5'b11101:
        casez_tmp_87 = ldq_29_valid;
      5'b11110:
        casez_tmp_87 = ldq_30_valid;
      default:
        casez_tmp_87 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_88;
  always @(*) begin
    casez (_GEN_6)
      5'b00000:
        casez_tmp_88 = stq_0_valid;
      5'b00001:
        casez_tmp_88 = stq_1_valid;
      5'b00010:
        casez_tmp_88 = stq_2_valid;
      5'b00011:
        casez_tmp_88 = stq_3_valid;
      5'b00100:
        casez_tmp_88 = stq_4_valid;
      5'b00101:
        casez_tmp_88 = stq_5_valid;
      5'b00110:
        casez_tmp_88 = stq_6_valid;
      5'b00111:
        casez_tmp_88 = stq_7_valid;
      5'b01000:
        casez_tmp_88 = stq_8_valid;
      5'b01001:
        casez_tmp_88 = stq_9_valid;
      5'b01010:
        casez_tmp_88 = stq_10_valid;
      5'b01011:
        casez_tmp_88 = stq_11_valid;
      5'b01100:
        casez_tmp_88 = stq_12_valid;
      5'b01101:
        casez_tmp_88 = stq_13_valid;
      5'b01110:
        casez_tmp_88 = stq_14_valid;
      5'b01111:
        casez_tmp_88 = stq_15_valid;
      5'b10000:
        casez_tmp_88 = stq_16_valid;
      5'b10001:
        casez_tmp_88 = stq_17_valid;
      5'b10010:
        casez_tmp_88 = stq_18_valid;
      5'b10011:
        casez_tmp_88 = stq_19_valid;
      5'b10100:
        casez_tmp_88 = stq_20_valid;
      5'b10101:
        casez_tmp_88 = stq_21_valid;
      5'b10110:
        casez_tmp_88 = stq_22_valid;
      5'b10111:
        casez_tmp_88 = stq_23_valid;
      5'b11000:
        casez_tmp_88 = stq_24_valid;
      5'b11001:
        casez_tmp_88 = stq_25_valid;
      5'b11010:
        casez_tmp_88 = stq_26_valid;
      5'b11011:
        casez_tmp_88 = stq_27_valid;
      5'b11100:
        casez_tmp_88 = stq_28_valid;
      5'b11101:
        casez_tmp_88 = stq_29_valid;
      5'b11110:
        casez_tmp_88 = stq_30_valid;
      default:
        casez_tmp_88 = stq_31_valid;
    endcase
  end // always @(*)
  wire [4:0]  _GEN_9 = dis_ld_val_1 ? _GEN_7 : _GEN_5;
  wire [4:0]  _GEN_10 = dis_st_val_1 ? _GEN_8 : _GEN_6;
  wire [4:0]  _GEN_11 = _GEN_9 + 5'h1;
  wire [4:0]  _GEN_12 = _GEN_10 + 5'h1;
  wire        dis_ld_val_2 = io_core_dis_uops_2_valid & io_core_dis_uops_2_bits_uses_ldq & ~io_core_dis_uops_2_bits_exception;
  wire        dis_st_val_2 = io_core_dis_uops_2_valid & io_core_dis_uops_2_bits_uses_stq & ~io_core_dis_uops_2_bits_exception;
  reg         casez_tmp_89;
  always @(*) begin
    casez (_GEN_9)
      5'b00000:
        casez_tmp_89 = ldq_0_valid;
      5'b00001:
        casez_tmp_89 = ldq_1_valid;
      5'b00010:
        casez_tmp_89 = ldq_2_valid;
      5'b00011:
        casez_tmp_89 = ldq_3_valid;
      5'b00100:
        casez_tmp_89 = ldq_4_valid;
      5'b00101:
        casez_tmp_89 = ldq_5_valid;
      5'b00110:
        casez_tmp_89 = ldq_6_valid;
      5'b00111:
        casez_tmp_89 = ldq_7_valid;
      5'b01000:
        casez_tmp_89 = ldq_8_valid;
      5'b01001:
        casez_tmp_89 = ldq_9_valid;
      5'b01010:
        casez_tmp_89 = ldq_10_valid;
      5'b01011:
        casez_tmp_89 = ldq_11_valid;
      5'b01100:
        casez_tmp_89 = ldq_12_valid;
      5'b01101:
        casez_tmp_89 = ldq_13_valid;
      5'b01110:
        casez_tmp_89 = ldq_14_valid;
      5'b01111:
        casez_tmp_89 = ldq_15_valid;
      5'b10000:
        casez_tmp_89 = ldq_16_valid;
      5'b10001:
        casez_tmp_89 = ldq_17_valid;
      5'b10010:
        casez_tmp_89 = ldq_18_valid;
      5'b10011:
        casez_tmp_89 = ldq_19_valid;
      5'b10100:
        casez_tmp_89 = ldq_20_valid;
      5'b10101:
        casez_tmp_89 = ldq_21_valid;
      5'b10110:
        casez_tmp_89 = ldq_22_valid;
      5'b10111:
        casez_tmp_89 = ldq_23_valid;
      5'b11000:
        casez_tmp_89 = ldq_24_valid;
      5'b11001:
        casez_tmp_89 = ldq_25_valid;
      5'b11010:
        casez_tmp_89 = ldq_26_valid;
      5'b11011:
        casez_tmp_89 = ldq_27_valid;
      5'b11100:
        casez_tmp_89 = ldq_28_valid;
      5'b11101:
        casez_tmp_89 = ldq_29_valid;
      5'b11110:
        casez_tmp_89 = ldq_30_valid;
      default:
        casez_tmp_89 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_90;
  always @(*) begin
    casez (_GEN_10)
      5'b00000:
        casez_tmp_90 = stq_0_valid;
      5'b00001:
        casez_tmp_90 = stq_1_valid;
      5'b00010:
        casez_tmp_90 = stq_2_valid;
      5'b00011:
        casez_tmp_90 = stq_3_valid;
      5'b00100:
        casez_tmp_90 = stq_4_valid;
      5'b00101:
        casez_tmp_90 = stq_5_valid;
      5'b00110:
        casez_tmp_90 = stq_6_valid;
      5'b00111:
        casez_tmp_90 = stq_7_valid;
      5'b01000:
        casez_tmp_90 = stq_8_valid;
      5'b01001:
        casez_tmp_90 = stq_9_valid;
      5'b01010:
        casez_tmp_90 = stq_10_valid;
      5'b01011:
        casez_tmp_90 = stq_11_valid;
      5'b01100:
        casez_tmp_90 = stq_12_valid;
      5'b01101:
        casez_tmp_90 = stq_13_valid;
      5'b01110:
        casez_tmp_90 = stq_14_valid;
      5'b01111:
        casez_tmp_90 = stq_15_valid;
      5'b10000:
        casez_tmp_90 = stq_16_valid;
      5'b10001:
        casez_tmp_90 = stq_17_valid;
      5'b10010:
        casez_tmp_90 = stq_18_valid;
      5'b10011:
        casez_tmp_90 = stq_19_valid;
      5'b10100:
        casez_tmp_90 = stq_20_valid;
      5'b10101:
        casez_tmp_90 = stq_21_valid;
      5'b10110:
        casez_tmp_90 = stq_22_valid;
      5'b10111:
        casez_tmp_90 = stq_23_valid;
      5'b11000:
        casez_tmp_90 = stq_24_valid;
      5'b11001:
        casez_tmp_90 = stq_25_valid;
      5'b11010:
        casez_tmp_90 = stq_26_valid;
      5'b11011:
        casez_tmp_90 = stq_27_valid;
      5'b11100:
        casez_tmp_90 = stq_28_valid;
      5'b11101:
        casez_tmp_90 = stq_29_valid;
      5'b11110:
        casez_tmp_90 = stq_30_valid;
      default:
        casez_tmp_90 = stq_31_valid;
    endcase
  end // always @(*)
  wire [4:0]  _GEN_13 = dis_ld_val_2 ? _GEN_11 : _GEN_9;
  wire [4:0]  _GEN_14 = dis_st_val_2 ? _GEN_12 : _GEN_10;
  wire [4:0]  _GEN_15 = _GEN_13 + 5'h1;
  wire [4:0]  _GEN_16 = _GEN_14 + 5'h1;
  wire        dis_ld_val_3 = io_core_dis_uops_3_valid & io_core_dis_uops_3_bits_uses_ldq & ~io_core_dis_uops_3_bits_exception;
  wire        dis_st_val_3 = io_core_dis_uops_3_valid & io_core_dis_uops_3_bits_uses_stq & ~io_core_dis_uops_3_bits_exception;
  reg         casez_tmp_91;
  always @(*) begin
    casez (_GEN_13)
      5'b00000:
        casez_tmp_91 = ldq_0_valid;
      5'b00001:
        casez_tmp_91 = ldq_1_valid;
      5'b00010:
        casez_tmp_91 = ldq_2_valid;
      5'b00011:
        casez_tmp_91 = ldq_3_valid;
      5'b00100:
        casez_tmp_91 = ldq_4_valid;
      5'b00101:
        casez_tmp_91 = ldq_5_valid;
      5'b00110:
        casez_tmp_91 = ldq_6_valid;
      5'b00111:
        casez_tmp_91 = ldq_7_valid;
      5'b01000:
        casez_tmp_91 = ldq_8_valid;
      5'b01001:
        casez_tmp_91 = ldq_9_valid;
      5'b01010:
        casez_tmp_91 = ldq_10_valid;
      5'b01011:
        casez_tmp_91 = ldq_11_valid;
      5'b01100:
        casez_tmp_91 = ldq_12_valid;
      5'b01101:
        casez_tmp_91 = ldq_13_valid;
      5'b01110:
        casez_tmp_91 = ldq_14_valid;
      5'b01111:
        casez_tmp_91 = ldq_15_valid;
      5'b10000:
        casez_tmp_91 = ldq_16_valid;
      5'b10001:
        casez_tmp_91 = ldq_17_valid;
      5'b10010:
        casez_tmp_91 = ldq_18_valid;
      5'b10011:
        casez_tmp_91 = ldq_19_valid;
      5'b10100:
        casez_tmp_91 = ldq_20_valid;
      5'b10101:
        casez_tmp_91 = ldq_21_valid;
      5'b10110:
        casez_tmp_91 = ldq_22_valid;
      5'b10111:
        casez_tmp_91 = ldq_23_valid;
      5'b11000:
        casez_tmp_91 = ldq_24_valid;
      5'b11001:
        casez_tmp_91 = ldq_25_valid;
      5'b11010:
        casez_tmp_91 = ldq_26_valid;
      5'b11011:
        casez_tmp_91 = ldq_27_valid;
      5'b11100:
        casez_tmp_91 = ldq_28_valid;
      5'b11101:
        casez_tmp_91 = ldq_29_valid;
      5'b11110:
        casez_tmp_91 = ldq_30_valid;
      default:
        casez_tmp_91 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_92;
  always @(*) begin
    casez (_GEN_14)
      5'b00000:
        casez_tmp_92 = stq_0_valid;
      5'b00001:
        casez_tmp_92 = stq_1_valid;
      5'b00010:
        casez_tmp_92 = stq_2_valid;
      5'b00011:
        casez_tmp_92 = stq_3_valid;
      5'b00100:
        casez_tmp_92 = stq_4_valid;
      5'b00101:
        casez_tmp_92 = stq_5_valid;
      5'b00110:
        casez_tmp_92 = stq_6_valid;
      5'b00111:
        casez_tmp_92 = stq_7_valid;
      5'b01000:
        casez_tmp_92 = stq_8_valid;
      5'b01001:
        casez_tmp_92 = stq_9_valid;
      5'b01010:
        casez_tmp_92 = stq_10_valid;
      5'b01011:
        casez_tmp_92 = stq_11_valid;
      5'b01100:
        casez_tmp_92 = stq_12_valid;
      5'b01101:
        casez_tmp_92 = stq_13_valid;
      5'b01110:
        casez_tmp_92 = stq_14_valid;
      5'b01111:
        casez_tmp_92 = stq_15_valid;
      5'b10000:
        casez_tmp_92 = stq_16_valid;
      5'b10001:
        casez_tmp_92 = stq_17_valid;
      5'b10010:
        casez_tmp_92 = stq_18_valid;
      5'b10011:
        casez_tmp_92 = stq_19_valid;
      5'b10100:
        casez_tmp_92 = stq_20_valid;
      5'b10101:
        casez_tmp_92 = stq_21_valid;
      5'b10110:
        casez_tmp_92 = stq_22_valid;
      5'b10111:
        casez_tmp_92 = stq_23_valid;
      5'b11000:
        casez_tmp_92 = stq_24_valid;
      5'b11001:
        casez_tmp_92 = stq_25_valid;
      5'b11010:
        casez_tmp_92 = stq_26_valid;
      5'b11011:
        casez_tmp_92 = stq_27_valid;
      5'b11100:
        casez_tmp_92 = stq_28_valid;
      5'b11101:
        casez_tmp_92 = stq_29_valid;
      5'b11110:
        casez_tmp_92 = stq_30_valid;
      default:
        casez_tmp_92 = stq_31_valid;
    endcase
  end // always @(*)
  wire [38:0] exe_req_0_bits_sfence_bits_addr = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_bits_addr : io_core_exe_0_req_bits_sfence_bits_addr;
  wire        exe_req_0_bits_sfence_valid = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_valid : io_core_exe_0_req_bits_sfence_valid;
  wire        exe_req_0_bits_mxcpt_valid = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_mxcpt_valid : io_core_exe_0_req_bits_mxcpt_valid;
  wire [39:0] exe_req_0_bits_addr = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_addr : io_core_exe_0_req_bits_addr;
  wire        _mem_incoming_uop_WIRE_0_fp_val = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_fp_val : io_core_exe_0_req_bits_uop_fp_val;
  wire [6:0]  _mem_incoming_uop_WIRE_0_pdst = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_pdst : io_core_exe_0_req_bits_uop_pdst;
  wire [4:0]  _mem_incoming_uop_WIRE_0_stq_idx = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_stq_idx : io_core_exe_0_req_bits_uop_stq_idx;
  wire [4:0]  _mem_incoming_uop_WIRE_0_ldq_idx = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ldq_idx : io_core_exe_0_req_bits_uop_ldq_idx;
  wire [6:0]  _mem_incoming_uop_WIRE_0_rob_idx = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_rob_idx : io_core_exe_0_req_bits_uop_rob_idx;
  wire [19:0] exe_req_0_bits_uop_br_mask = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_br_mask : io_core_exe_0_req_bits_uop_br_mask;
  wire        exe_req_0_bits_uop_ctrl_is_std = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_is_std : io_core_exe_0_req_bits_uop_ctrl_is_std;
  wire        exe_req_0_bits_uop_ctrl_is_sta = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_is_sta : io_core_exe_0_req_bits_uop_ctrl_is_sta;
  wire        exe_req_0_bits_uop_ctrl_is_load = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_is_load : io_core_exe_0_req_bits_uop_ctrl_is_load;
  wire        exe_req_0_valid = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_valid : io_core_exe_0_req_valid;
  wire        _GEN_17 = io_core_exe_1_req_bits_sfence_valid | ~io_core_exe_0_req_bits_sfence_valid;
  wire [38:0] exe_req_1_bits_sfence_bits_addr = _GEN_17 ? io_core_exe_1_req_bits_sfence_bits_addr : io_core_exe_0_req_bits_sfence_bits_addr;
  wire        exe_req_1_bits_sfence_valid = _GEN_17 ? io_core_exe_1_req_bits_sfence_valid : io_core_exe_0_req_bits_sfence_valid;
  wire        exe_req_1_bits_mxcpt_valid = _GEN_17 ? io_core_exe_1_req_bits_mxcpt_valid : io_core_exe_0_req_bits_mxcpt_valid;
  wire [39:0] exe_req_1_bits_addr = _GEN_17 ? io_core_exe_1_req_bits_addr : io_core_exe_0_req_bits_addr;
  wire        _mem_incoming_uop_WIRE_1_fp_val = _GEN_17 ? io_core_exe_1_req_bits_uop_fp_val : io_core_exe_0_req_bits_uop_fp_val;
  wire [6:0]  _mem_incoming_uop_WIRE_1_pdst = _GEN_17 ? io_core_exe_1_req_bits_uop_pdst : io_core_exe_0_req_bits_uop_pdst;
  wire [4:0]  _mem_incoming_uop_WIRE_1_stq_idx = _GEN_17 ? io_core_exe_1_req_bits_uop_stq_idx : io_core_exe_0_req_bits_uop_stq_idx;
  wire [4:0]  _mem_incoming_uop_WIRE_1_ldq_idx = _GEN_17 ? io_core_exe_1_req_bits_uop_ldq_idx : io_core_exe_0_req_bits_uop_ldq_idx;
  wire [6:0]  _mem_incoming_uop_WIRE_1_rob_idx = _GEN_17 ? io_core_exe_1_req_bits_uop_rob_idx : io_core_exe_0_req_bits_uop_rob_idx;
  wire [19:0] exe_req_1_bits_uop_br_mask = _GEN_17 ? io_core_exe_1_req_bits_uop_br_mask : io_core_exe_0_req_bits_uop_br_mask;
  wire        exe_req_1_bits_uop_ctrl_is_std = _GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_is_std : io_core_exe_0_req_bits_uop_ctrl_is_std;
  wire        exe_req_1_bits_uop_ctrl_is_sta = _GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_is_sta : io_core_exe_0_req_bits_uop_ctrl_is_sta;
  wire        exe_req_1_bits_uop_ctrl_is_load = _GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_is_load : io_core_exe_0_req_bits_uop_ctrl_is_load;
  wire        exe_req_1_valid = _GEN_17 ? io_core_exe_1_req_valid : io_core_exe_0_req_valid;
  reg         p1_block_load_mask_0;
  reg         p1_block_load_mask_1;
  reg         p1_block_load_mask_2;
  reg         p1_block_load_mask_3;
  reg         p1_block_load_mask_4;
  reg         p1_block_load_mask_5;
  reg         p1_block_load_mask_6;
  reg         p1_block_load_mask_7;
  reg         p1_block_load_mask_8;
  reg         p1_block_load_mask_9;
  reg         p1_block_load_mask_10;
  reg         p1_block_load_mask_11;
  reg         p1_block_load_mask_12;
  reg         p1_block_load_mask_13;
  reg         p1_block_load_mask_14;
  reg         p1_block_load_mask_15;
  reg         p1_block_load_mask_16;
  reg         p1_block_load_mask_17;
  reg         p1_block_load_mask_18;
  reg         p1_block_load_mask_19;
  reg         p1_block_load_mask_20;
  reg         p1_block_load_mask_21;
  reg         p1_block_load_mask_22;
  reg         p1_block_load_mask_23;
  reg         p1_block_load_mask_24;
  reg         p1_block_load_mask_25;
  reg         p1_block_load_mask_26;
  reg         p1_block_load_mask_27;
  reg         p1_block_load_mask_28;
  reg         p1_block_load_mask_29;
  reg         p1_block_load_mask_30;
  reg         p1_block_load_mask_31;
  reg         p2_block_load_mask_0;
  reg         p2_block_load_mask_1;
  reg         p2_block_load_mask_2;
  reg         p2_block_load_mask_3;
  reg         p2_block_load_mask_4;
  reg         p2_block_load_mask_5;
  reg         p2_block_load_mask_6;
  reg         p2_block_load_mask_7;
  reg         p2_block_load_mask_8;
  reg         p2_block_load_mask_9;
  reg         p2_block_load_mask_10;
  reg         p2_block_load_mask_11;
  reg         p2_block_load_mask_12;
  reg         p2_block_load_mask_13;
  reg         p2_block_load_mask_14;
  reg         p2_block_load_mask_15;
  reg         p2_block_load_mask_16;
  reg         p2_block_load_mask_17;
  reg         p2_block_load_mask_18;
  reg         p2_block_load_mask_19;
  reg         p2_block_load_mask_20;
  reg         p2_block_load_mask_21;
  reg         p2_block_load_mask_22;
  reg         p2_block_load_mask_23;
  reg         p2_block_load_mask_24;
  reg         p2_block_load_mask_25;
  reg         p2_block_load_mask_26;
  reg         p2_block_load_mask_27;
  reg         p2_block_load_mask_28;
  reg         p2_block_load_mask_29;
  reg         p2_block_load_mask_30;
  reg         p2_block_load_mask_31;
  reg  [19:0] casez_tmp_93;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_ldq_idx)
      5'b00000:
        casez_tmp_93 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_93 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_93 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_93 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_93 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_93 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_93 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_93 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_93 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_93 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_93 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_93 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_93 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_93 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_93 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_93 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_93 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_93 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_93 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_93 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_93 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_93 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_93 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_93 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_93 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_93 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_93 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_93 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_93 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_93 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_93 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_93 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_94;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_ldq_idx)
      5'b00000:
        casez_tmp_94 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_94 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_94 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_94 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_94 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_94 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_94 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_94 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_94 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_94 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_94 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_94 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_94 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_94 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_94 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_94 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_94 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_94 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_94 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_94 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_94 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_94 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_94 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_94 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_94 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_94 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_94 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_94 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_94 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_94 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_94 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_94 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_95;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_ldq_idx)
      5'b00000:
        casez_tmp_95 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_95 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_95 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_95 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_95 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_95 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_95 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_95 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_95 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_95 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_95 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_95 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_95 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_95 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_95 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_95 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_95 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_95 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_95 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_95 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_95 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_95 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_95 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_95 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_95 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_95 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_95 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_95 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_95 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_95 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_95 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_95 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_96;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_ldq_idx)
      5'b00000:
        casez_tmp_96 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_96 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_96 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_96 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_96 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_96 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_96 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_96 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_96 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_96 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_96 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_96 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_96 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_96 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_96 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_96 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_96 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_96 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_96 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_96 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_96 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_96 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_96 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_96 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_96 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_96 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_96 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_96 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_96 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_96 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_96 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_96 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_97;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_ldq_idx)
      5'b00000:
        casez_tmp_97 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_97 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_97 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_97 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_97 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_97 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_97 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_97 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_97 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_97 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_97 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_97 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_97 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_97 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_97 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_97 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_97 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_97 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_97 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_97 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_97 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_97 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_97 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_97 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_97 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_97 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_97 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_97 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_97 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_97 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_97 = ldq_30_bits_executed;
      default:
        casez_tmp_97 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_98;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_ldq_idx)
      5'b00000:
        casez_tmp_98 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_98 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_98 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_98 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_98 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_98 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_98 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_98 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_98 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_98 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_98 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_98 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_98 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_98 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_98 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_98 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_98 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_98 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_98 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_98 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_98 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_98 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_98 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_98 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_98 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_98 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_98 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_98 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_98 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_98 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_98 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_98 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_99;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_ldq_idx)
      5'b00000:
        casez_tmp_99 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_99 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_99 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_99 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_99 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_99 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_99 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_99 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_99 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_99 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_99 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_99 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_99 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_99 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_99 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_99 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_99 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_99 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_99 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_99 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_99 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_99 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_99 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_99 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_99 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_99 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_99 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_99 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_99 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_99 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_99 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_99 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_100;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_ldq_idx)
      5'b00000:
        casez_tmp_100 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_100 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_100 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_100 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_100 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_100 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_100 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_100 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_100 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_100 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_100 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_100 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_100 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_100 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_100 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_100 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_100 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_100 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_100 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_100 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_100 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_100 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_100 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_100 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_100 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_100 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_100 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_100 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_100 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_100 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_100 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_100 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_101;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_ldq_idx)
      5'b00000:
        casez_tmp_101 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_101 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_101 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_101 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_101 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_101 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_101 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_101 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_101 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_101 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_101 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_101 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_101 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_101 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_101 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_101 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_101 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_101 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_101 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_101 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_101 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_101 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_101 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_101 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_101 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_101 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_101 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_101 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_101 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_101 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_101 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_101 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_102;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_ldq_idx)
      5'b00000:
        casez_tmp_102 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_102 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_102 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_102 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_102 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_102 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_102 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_102 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_102 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_102 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_102 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_102 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_102 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_102 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_102 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_102 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_102 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_102 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_102 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_102 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_102 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_102 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_102 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_102 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_102 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_102 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_102 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_102 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_102 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_102 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_102 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_102 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_103;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_ldq_idx)
      5'b00000:
        casez_tmp_103 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_103 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_103 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_103 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_103 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_103 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_103 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_103 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_103 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_103 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_103 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_103 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_103 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_103 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_103 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_103 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_103 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_103 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_103 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_103 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_103 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_103 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_103 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_103 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_103 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_103 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_103 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_103 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_103 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_103 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_103 = ldq_30_bits_executed;
      default:
        casez_tmp_103 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_104;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_ldq_idx)
      5'b00000:
        casez_tmp_104 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_104 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_104 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_104 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_104 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_104 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_104 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_104 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_104 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_104 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_104 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_104 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_104 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_104 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_104 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_104 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_104 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_104 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_104 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_104 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_104 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_104 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_104 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_104 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_104 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_104 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_104 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_104 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_104 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_104 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_104 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_104 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  reg         casez_tmp_105;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_105 = stq_0_valid;
      5'b00001:
        casez_tmp_105 = stq_1_valid;
      5'b00010:
        casez_tmp_105 = stq_2_valid;
      5'b00011:
        casez_tmp_105 = stq_3_valid;
      5'b00100:
        casez_tmp_105 = stq_4_valid;
      5'b00101:
        casez_tmp_105 = stq_5_valid;
      5'b00110:
        casez_tmp_105 = stq_6_valid;
      5'b00111:
        casez_tmp_105 = stq_7_valid;
      5'b01000:
        casez_tmp_105 = stq_8_valid;
      5'b01001:
        casez_tmp_105 = stq_9_valid;
      5'b01010:
        casez_tmp_105 = stq_10_valid;
      5'b01011:
        casez_tmp_105 = stq_11_valid;
      5'b01100:
        casez_tmp_105 = stq_12_valid;
      5'b01101:
        casez_tmp_105 = stq_13_valid;
      5'b01110:
        casez_tmp_105 = stq_14_valid;
      5'b01111:
        casez_tmp_105 = stq_15_valid;
      5'b10000:
        casez_tmp_105 = stq_16_valid;
      5'b10001:
        casez_tmp_105 = stq_17_valid;
      5'b10010:
        casez_tmp_105 = stq_18_valid;
      5'b10011:
        casez_tmp_105 = stq_19_valid;
      5'b10100:
        casez_tmp_105 = stq_20_valid;
      5'b10101:
        casez_tmp_105 = stq_21_valid;
      5'b10110:
        casez_tmp_105 = stq_22_valid;
      5'b10111:
        casez_tmp_105 = stq_23_valid;
      5'b11000:
        casez_tmp_105 = stq_24_valid;
      5'b11001:
        casez_tmp_105 = stq_25_valid;
      5'b11010:
        casez_tmp_105 = stq_26_valid;
      5'b11011:
        casez_tmp_105 = stq_27_valid;
      5'b11100:
        casez_tmp_105 = stq_28_valid;
      5'b11101:
        casez_tmp_105 = stq_29_valid;
      5'b11110:
        casez_tmp_105 = stq_30_valid;
      default:
        casez_tmp_105 = stq_31_valid;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_106;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_106 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_106 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_106 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_106 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_106 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_106 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_106 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_106 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_106 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_106 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_106 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_106 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_106 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_106 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_106 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_106 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_106 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_106 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_106 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_106 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_106 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_106 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_106 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_106 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_106 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_106 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_106 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_106 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_106 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_106 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_106 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_106 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_107;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_107 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_107 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_107 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_107 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_107 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_107 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_107 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_107 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_107 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_107 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_107 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_107 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_107 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_107 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_107 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_107 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_107 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_107 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_107 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_107 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_107 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_107 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_107 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_107 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_107 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_107 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_107 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_107 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_107 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_107 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_107 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_107 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_108;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_108 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_108 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_108 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_108 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_108 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_108 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_108 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_108 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_108 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_108 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_108 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_108 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_108 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_108 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_108 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_108 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_108 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_108 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_108 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_108 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_108 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_108 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_108 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_108 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_108 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_108 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_108 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_108 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_108 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_108 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_108 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_108 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_109;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_109 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_109 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_109 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_109 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_109 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_109 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_109 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_109 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_109 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_109 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_109 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_109 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_109 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_109 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_109 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_109 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_109 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_109 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_109 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_109 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_109 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_109 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_109 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_109 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_109 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_109 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_109 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_109 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_109 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_109 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_109 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_109 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_110;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_110 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_110 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_110 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_110 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_110 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_110 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_110 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_110 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_110 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_110 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_110 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_110 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_110 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_110 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_110 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_110 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_110 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_110 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_110 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_110 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_110 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_110 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_110 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_110 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_110 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_110 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_110 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_110 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_110 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_110 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_110 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_110 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_111;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_111 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_111 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_111 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_111 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_111 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_111 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_111 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_111 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_111 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_111 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_111 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_111 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_111 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_111 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_111 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_111 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_111 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_111 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_111 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_111 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_111 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_111 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_111 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_111 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_111 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_111 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_111 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_111 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_111 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_111 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_111 = stq_30_bits_addr_valid;
      default:
        casez_tmp_111 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_112;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_112 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_112 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_112 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_112 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_112 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_112 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_112 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_112 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_112 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_112 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_112 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_112 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_112 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_112 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_112 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_112 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_112 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_112 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_112 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_112 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_112 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_112 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_112 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_112 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_112 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_112 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_112 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_112 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_112 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_112 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_112 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_112 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         casez_tmp_113;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_0_stq_idx)
      5'b00000:
        casez_tmp_113 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_113 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_113 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_113 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_113 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_113 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_113 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_113 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_113 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_113 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_113 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_113 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_113 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_113 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_113 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_113 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_113 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_113 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_113 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_113 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_113 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_113 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_113 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_113 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_113 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_113 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_113 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_113 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_113 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_113 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_113 = stq_30_bits_data_valid;
      default:
        casez_tmp_113 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_114;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_114 = stq_0_valid;
      5'b00001:
        casez_tmp_114 = stq_1_valid;
      5'b00010:
        casez_tmp_114 = stq_2_valid;
      5'b00011:
        casez_tmp_114 = stq_3_valid;
      5'b00100:
        casez_tmp_114 = stq_4_valid;
      5'b00101:
        casez_tmp_114 = stq_5_valid;
      5'b00110:
        casez_tmp_114 = stq_6_valid;
      5'b00111:
        casez_tmp_114 = stq_7_valid;
      5'b01000:
        casez_tmp_114 = stq_8_valid;
      5'b01001:
        casez_tmp_114 = stq_9_valid;
      5'b01010:
        casez_tmp_114 = stq_10_valid;
      5'b01011:
        casez_tmp_114 = stq_11_valid;
      5'b01100:
        casez_tmp_114 = stq_12_valid;
      5'b01101:
        casez_tmp_114 = stq_13_valid;
      5'b01110:
        casez_tmp_114 = stq_14_valid;
      5'b01111:
        casez_tmp_114 = stq_15_valid;
      5'b10000:
        casez_tmp_114 = stq_16_valid;
      5'b10001:
        casez_tmp_114 = stq_17_valid;
      5'b10010:
        casez_tmp_114 = stq_18_valid;
      5'b10011:
        casez_tmp_114 = stq_19_valid;
      5'b10100:
        casez_tmp_114 = stq_20_valid;
      5'b10101:
        casez_tmp_114 = stq_21_valid;
      5'b10110:
        casez_tmp_114 = stq_22_valid;
      5'b10111:
        casez_tmp_114 = stq_23_valid;
      5'b11000:
        casez_tmp_114 = stq_24_valid;
      5'b11001:
        casez_tmp_114 = stq_25_valid;
      5'b11010:
        casez_tmp_114 = stq_26_valid;
      5'b11011:
        casez_tmp_114 = stq_27_valid;
      5'b11100:
        casez_tmp_114 = stq_28_valid;
      5'b11101:
        casez_tmp_114 = stq_29_valid;
      5'b11110:
        casez_tmp_114 = stq_30_valid;
      default:
        casez_tmp_114 = stq_31_valid;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_115;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_115 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_115 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_115 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_115 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_115 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_115 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_115 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_115 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_115 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_115 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_115 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_115 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_115 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_115 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_115 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_115 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_115 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_115 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_115 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_115 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_115 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_115 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_115 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_115 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_115 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_115 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_115 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_115 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_115 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_115 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_115 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_115 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_116;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_116 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_116 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_116 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_116 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_116 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_116 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_116 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_116 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_116 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_116 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_116 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_116 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_116 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_116 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_116 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_116 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_116 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_116 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_116 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_116 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_116 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_116 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_116 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_116 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_116 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_116 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_116 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_116 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_116 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_116 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_116 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_116 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_117;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_117 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_117 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_117 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_117 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_117 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_117 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_117 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_117 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_117 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_117 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_117 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_117 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_117 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_117 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_117 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_117 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_117 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_117 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_117 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_117 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_117 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_117 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_117 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_117 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_117 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_117 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_117 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_117 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_117 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_117 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_117 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_117 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_118;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_118 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_118 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_118 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_118 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_118 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_118 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_118 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_118 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_118 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_118 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_118 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_118 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_118 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_118 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_118 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_118 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_118 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_118 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_118 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_118 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_118 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_118 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_118 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_118 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_118 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_118 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_118 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_118 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_118 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_118 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_118 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_118 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_119;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_119 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_119 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_119 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_119 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_119 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_119 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_119 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_119 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_119 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_119 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_119 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_119 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_119 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_119 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_119 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_119 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_119 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_119 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_119 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_119 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_119 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_119 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_119 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_119 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_119 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_119 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_119 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_119 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_119 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_119 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_119 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_119 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_120;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_120 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_120 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_120 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_120 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_120 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_120 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_120 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_120 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_120 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_120 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_120 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_120 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_120 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_120 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_120 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_120 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_120 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_120 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_120 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_120 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_120 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_120 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_120 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_120 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_120 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_120 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_120 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_120 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_120 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_120 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_120 = stq_30_bits_addr_valid;
      default:
        casez_tmp_120 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_121;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_121 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_121 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_121 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_121 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_121 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_121 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_121 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_121 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_121 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_121 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_121 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_121 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_121 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_121 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_121 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_121 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_121 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_121 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_121 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_121 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_121 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_121 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_121 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_121 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_121 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_121 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_121 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_121 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_121 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_121 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_121 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_121 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         casez_tmp_122;
  always @(*) begin
    casez (_mem_incoming_uop_WIRE_1_stq_idx)
      5'b00000:
        casez_tmp_122 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_122 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_122 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_122 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_122 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_122 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_122 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_122 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_122 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_122 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_122 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_122 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_122 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_122 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_122 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_122 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_122 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_122 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_122 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_122 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_122 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_122 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_122 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_122 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_122 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_122 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_122 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_122 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_122 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_122 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_122 = stq_30_bits_data_valid;
      default:
        casez_tmp_122 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  wire        _temp_bits_T = ldq_head == 5'h0;
  wire        _temp_bits_T_2 = ldq_head < 5'h2;
  wire        _temp_bits_T_4 = ldq_head < 5'h3;
  wire        _temp_bits_T_6 = ldq_head < 5'h4;
  wire        _temp_bits_T_8 = ldq_head < 5'h5;
  wire        _temp_bits_T_10 = ldq_head < 5'h6;
  wire        _temp_bits_T_12 = ldq_head < 5'h7;
  wire        _temp_bits_T_14 = ldq_head < 5'h8;
  wire        _temp_bits_T_16 = ldq_head < 5'h9;
  wire        _temp_bits_T_18 = ldq_head < 5'hA;
  wire        _temp_bits_T_20 = ldq_head < 5'hB;
  wire        _temp_bits_T_22 = ldq_head < 5'hC;
  wire        _temp_bits_T_24 = ldq_head < 5'hD;
  wire        _temp_bits_T_26 = ldq_head < 5'hE;
  wire        _temp_bits_T_28 = ldq_head < 5'hF;
  wire        _temp_bits_T_32 = ldq_head < 5'h11;
  wire        _temp_bits_T_34 = ldq_head < 5'h12;
  wire        _temp_bits_T_36 = ldq_head < 5'h13;
  wire        _temp_bits_T_38 = ldq_head < 5'h14;
  wire        _temp_bits_T_40 = ldq_head < 5'h15;
  wire        _temp_bits_T_42 = ldq_head < 5'h16;
  wire        _temp_bits_T_44 = ldq_head < 5'h17;
  wire        _temp_bits_T_46 = ldq_head[4:3] != 2'h3;
  wire        _temp_bits_T_48 = ldq_head < 5'h19;
  wire        _temp_bits_T_50 = ldq_head < 5'h1A;
  wire        _temp_bits_T_52 = ldq_head < 5'h1B;
  wire        _temp_bits_T_54 = ldq_head[4:2] != 3'h7;
  wire        _temp_bits_T_56 = ldq_head < 5'h1D;
  wire        _temp_bits_T_58 = ldq_head[4:1] != 4'hF;
  wire        _temp_bits_T_60 = ldq_head != 5'h1F;
  reg  [4:0]  ldq_retry_idx;
  reg  [4:0]  stq_retry_idx;
  reg  [4:0]  ldq_wakeup_idx;
  wire        will_fire_load_incoming_0_will_fire = exe_req_0_valid & exe_req_0_bits_uop_ctrl_is_load;
  wire        will_fire_load_incoming_1_will_fire = exe_req_1_valid & exe_req_1_bits_uop_ctrl_is_load;
  wire        _can_fire_sta_incoming_T = exe_req_0_valid & exe_req_0_bits_uop_ctrl_is_sta;
  wire        _can_fire_sta_incoming_T_3 = exe_req_1_valid & exe_req_1_bits_uop_ctrl_is_sta;
  wire        can_fire_std_incoming_0 = exe_req_0_valid & exe_req_0_bits_uop_ctrl_is_std & ~exe_req_0_bits_uop_ctrl_is_sta;
  wire        will_fire_release_1_will_fire;
  reg         casez_tmp_123;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_123 = ldq_0_valid;
      5'b00001:
        casez_tmp_123 = ldq_1_valid;
      5'b00010:
        casez_tmp_123 = ldq_2_valid;
      5'b00011:
        casez_tmp_123 = ldq_3_valid;
      5'b00100:
        casez_tmp_123 = ldq_4_valid;
      5'b00101:
        casez_tmp_123 = ldq_5_valid;
      5'b00110:
        casez_tmp_123 = ldq_6_valid;
      5'b00111:
        casez_tmp_123 = ldq_7_valid;
      5'b01000:
        casez_tmp_123 = ldq_8_valid;
      5'b01001:
        casez_tmp_123 = ldq_9_valid;
      5'b01010:
        casez_tmp_123 = ldq_10_valid;
      5'b01011:
        casez_tmp_123 = ldq_11_valid;
      5'b01100:
        casez_tmp_123 = ldq_12_valid;
      5'b01101:
        casez_tmp_123 = ldq_13_valid;
      5'b01110:
        casez_tmp_123 = ldq_14_valid;
      5'b01111:
        casez_tmp_123 = ldq_15_valid;
      5'b10000:
        casez_tmp_123 = ldq_16_valid;
      5'b10001:
        casez_tmp_123 = ldq_17_valid;
      5'b10010:
        casez_tmp_123 = ldq_18_valid;
      5'b10011:
        casez_tmp_123 = ldq_19_valid;
      5'b10100:
        casez_tmp_123 = ldq_20_valid;
      5'b10101:
        casez_tmp_123 = ldq_21_valid;
      5'b10110:
        casez_tmp_123 = ldq_22_valid;
      5'b10111:
        casez_tmp_123 = ldq_23_valid;
      5'b11000:
        casez_tmp_123 = ldq_24_valid;
      5'b11001:
        casez_tmp_123 = ldq_25_valid;
      5'b11010:
        casez_tmp_123 = ldq_26_valid;
      5'b11011:
        casez_tmp_123 = ldq_27_valid;
      5'b11100:
        casez_tmp_123 = ldq_28_valid;
      5'b11101:
        casez_tmp_123 = ldq_29_valid;
      5'b11110:
        casez_tmp_123 = ldq_30_valid;
      default:
        casez_tmp_123 = ldq_31_valid;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_124;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_124 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_124 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_124 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_124 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_124 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_124 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_124 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_124 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_124 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_124 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_124 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_124 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_124 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_124 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_124 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_124 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_124 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_124 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_124 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_124 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_124 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_124 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_124 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_124 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_124 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_124 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_124 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_124 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_124 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_124 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_124 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_124 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_125;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_125 = ldq_0_bits_uop_inst;
      5'b00001:
        casez_tmp_125 = ldq_1_bits_uop_inst;
      5'b00010:
        casez_tmp_125 = ldq_2_bits_uop_inst;
      5'b00011:
        casez_tmp_125 = ldq_3_bits_uop_inst;
      5'b00100:
        casez_tmp_125 = ldq_4_bits_uop_inst;
      5'b00101:
        casez_tmp_125 = ldq_5_bits_uop_inst;
      5'b00110:
        casez_tmp_125 = ldq_6_bits_uop_inst;
      5'b00111:
        casez_tmp_125 = ldq_7_bits_uop_inst;
      5'b01000:
        casez_tmp_125 = ldq_8_bits_uop_inst;
      5'b01001:
        casez_tmp_125 = ldq_9_bits_uop_inst;
      5'b01010:
        casez_tmp_125 = ldq_10_bits_uop_inst;
      5'b01011:
        casez_tmp_125 = ldq_11_bits_uop_inst;
      5'b01100:
        casez_tmp_125 = ldq_12_bits_uop_inst;
      5'b01101:
        casez_tmp_125 = ldq_13_bits_uop_inst;
      5'b01110:
        casez_tmp_125 = ldq_14_bits_uop_inst;
      5'b01111:
        casez_tmp_125 = ldq_15_bits_uop_inst;
      5'b10000:
        casez_tmp_125 = ldq_16_bits_uop_inst;
      5'b10001:
        casez_tmp_125 = ldq_17_bits_uop_inst;
      5'b10010:
        casez_tmp_125 = ldq_18_bits_uop_inst;
      5'b10011:
        casez_tmp_125 = ldq_19_bits_uop_inst;
      5'b10100:
        casez_tmp_125 = ldq_20_bits_uop_inst;
      5'b10101:
        casez_tmp_125 = ldq_21_bits_uop_inst;
      5'b10110:
        casez_tmp_125 = ldq_22_bits_uop_inst;
      5'b10111:
        casez_tmp_125 = ldq_23_bits_uop_inst;
      5'b11000:
        casez_tmp_125 = ldq_24_bits_uop_inst;
      5'b11001:
        casez_tmp_125 = ldq_25_bits_uop_inst;
      5'b11010:
        casez_tmp_125 = ldq_26_bits_uop_inst;
      5'b11011:
        casez_tmp_125 = ldq_27_bits_uop_inst;
      5'b11100:
        casez_tmp_125 = ldq_28_bits_uop_inst;
      5'b11101:
        casez_tmp_125 = ldq_29_bits_uop_inst;
      5'b11110:
        casez_tmp_125 = ldq_30_bits_uop_inst;
      default:
        casez_tmp_125 = ldq_31_bits_uop_inst;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_126;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_126 = ldq_0_bits_uop_debug_inst;
      5'b00001:
        casez_tmp_126 = ldq_1_bits_uop_debug_inst;
      5'b00010:
        casez_tmp_126 = ldq_2_bits_uop_debug_inst;
      5'b00011:
        casez_tmp_126 = ldq_3_bits_uop_debug_inst;
      5'b00100:
        casez_tmp_126 = ldq_4_bits_uop_debug_inst;
      5'b00101:
        casez_tmp_126 = ldq_5_bits_uop_debug_inst;
      5'b00110:
        casez_tmp_126 = ldq_6_bits_uop_debug_inst;
      5'b00111:
        casez_tmp_126 = ldq_7_bits_uop_debug_inst;
      5'b01000:
        casez_tmp_126 = ldq_8_bits_uop_debug_inst;
      5'b01001:
        casez_tmp_126 = ldq_9_bits_uop_debug_inst;
      5'b01010:
        casez_tmp_126 = ldq_10_bits_uop_debug_inst;
      5'b01011:
        casez_tmp_126 = ldq_11_bits_uop_debug_inst;
      5'b01100:
        casez_tmp_126 = ldq_12_bits_uop_debug_inst;
      5'b01101:
        casez_tmp_126 = ldq_13_bits_uop_debug_inst;
      5'b01110:
        casez_tmp_126 = ldq_14_bits_uop_debug_inst;
      5'b01111:
        casez_tmp_126 = ldq_15_bits_uop_debug_inst;
      5'b10000:
        casez_tmp_126 = ldq_16_bits_uop_debug_inst;
      5'b10001:
        casez_tmp_126 = ldq_17_bits_uop_debug_inst;
      5'b10010:
        casez_tmp_126 = ldq_18_bits_uop_debug_inst;
      5'b10011:
        casez_tmp_126 = ldq_19_bits_uop_debug_inst;
      5'b10100:
        casez_tmp_126 = ldq_20_bits_uop_debug_inst;
      5'b10101:
        casez_tmp_126 = ldq_21_bits_uop_debug_inst;
      5'b10110:
        casez_tmp_126 = ldq_22_bits_uop_debug_inst;
      5'b10111:
        casez_tmp_126 = ldq_23_bits_uop_debug_inst;
      5'b11000:
        casez_tmp_126 = ldq_24_bits_uop_debug_inst;
      5'b11001:
        casez_tmp_126 = ldq_25_bits_uop_debug_inst;
      5'b11010:
        casez_tmp_126 = ldq_26_bits_uop_debug_inst;
      5'b11011:
        casez_tmp_126 = ldq_27_bits_uop_debug_inst;
      5'b11100:
        casez_tmp_126 = ldq_28_bits_uop_debug_inst;
      5'b11101:
        casez_tmp_126 = ldq_29_bits_uop_debug_inst;
      5'b11110:
        casez_tmp_126 = ldq_30_bits_uop_debug_inst;
      default:
        casez_tmp_126 = ldq_31_bits_uop_debug_inst;
    endcase
  end // always @(*)
  reg         casez_tmp_127;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_127 = ldq_0_bits_uop_is_rvc;
      5'b00001:
        casez_tmp_127 = ldq_1_bits_uop_is_rvc;
      5'b00010:
        casez_tmp_127 = ldq_2_bits_uop_is_rvc;
      5'b00011:
        casez_tmp_127 = ldq_3_bits_uop_is_rvc;
      5'b00100:
        casez_tmp_127 = ldq_4_bits_uop_is_rvc;
      5'b00101:
        casez_tmp_127 = ldq_5_bits_uop_is_rvc;
      5'b00110:
        casez_tmp_127 = ldq_6_bits_uop_is_rvc;
      5'b00111:
        casez_tmp_127 = ldq_7_bits_uop_is_rvc;
      5'b01000:
        casez_tmp_127 = ldq_8_bits_uop_is_rvc;
      5'b01001:
        casez_tmp_127 = ldq_9_bits_uop_is_rvc;
      5'b01010:
        casez_tmp_127 = ldq_10_bits_uop_is_rvc;
      5'b01011:
        casez_tmp_127 = ldq_11_bits_uop_is_rvc;
      5'b01100:
        casez_tmp_127 = ldq_12_bits_uop_is_rvc;
      5'b01101:
        casez_tmp_127 = ldq_13_bits_uop_is_rvc;
      5'b01110:
        casez_tmp_127 = ldq_14_bits_uop_is_rvc;
      5'b01111:
        casez_tmp_127 = ldq_15_bits_uop_is_rvc;
      5'b10000:
        casez_tmp_127 = ldq_16_bits_uop_is_rvc;
      5'b10001:
        casez_tmp_127 = ldq_17_bits_uop_is_rvc;
      5'b10010:
        casez_tmp_127 = ldq_18_bits_uop_is_rvc;
      5'b10011:
        casez_tmp_127 = ldq_19_bits_uop_is_rvc;
      5'b10100:
        casez_tmp_127 = ldq_20_bits_uop_is_rvc;
      5'b10101:
        casez_tmp_127 = ldq_21_bits_uop_is_rvc;
      5'b10110:
        casez_tmp_127 = ldq_22_bits_uop_is_rvc;
      5'b10111:
        casez_tmp_127 = ldq_23_bits_uop_is_rvc;
      5'b11000:
        casez_tmp_127 = ldq_24_bits_uop_is_rvc;
      5'b11001:
        casez_tmp_127 = ldq_25_bits_uop_is_rvc;
      5'b11010:
        casez_tmp_127 = ldq_26_bits_uop_is_rvc;
      5'b11011:
        casez_tmp_127 = ldq_27_bits_uop_is_rvc;
      5'b11100:
        casez_tmp_127 = ldq_28_bits_uop_is_rvc;
      5'b11101:
        casez_tmp_127 = ldq_29_bits_uop_is_rvc;
      5'b11110:
        casez_tmp_127 = ldq_30_bits_uop_is_rvc;
      default:
        casez_tmp_127 = ldq_31_bits_uop_is_rvc;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_128;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_128 = ldq_0_bits_uop_debug_pc;
      5'b00001:
        casez_tmp_128 = ldq_1_bits_uop_debug_pc;
      5'b00010:
        casez_tmp_128 = ldq_2_bits_uop_debug_pc;
      5'b00011:
        casez_tmp_128 = ldq_3_bits_uop_debug_pc;
      5'b00100:
        casez_tmp_128 = ldq_4_bits_uop_debug_pc;
      5'b00101:
        casez_tmp_128 = ldq_5_bits_uop_debug_pc;
      5'b00110:
        casez_tmp_128 = ldq_6_bits_uop_debug_pc;
      5'b00111:
        casez_tmp_128 = ldq_7_bits_uop_debug_pc;
      5'b01000:
        casez_tmp_128 = ldq_8_bits_uop_debug_pc;
      5'b01001:
        casez_tmp_128 = ldq_9_bits_uop_debug_pc;
      5'b01010:
        casez_tmp_128 = ldq_10_bits_uop_debug_pc;
      5'b01011:
        casez_tmp_128 = ldq_11_bits_uop_debug_pc;
      5'b01100:
        casez_tmp_128 = ldq_12_bits_uop_debug_pc;
      5'b01101:
        casez_tmp_128 = ldq_13_bits_uop_debug_pc;
      5'b01110:
        casez_tmp_128 = ldq_14_bits_uop_debug_pc;
      5'b01111:
        casez_tmp_128 = ldq_15_bits_uop_debug_pc;
      5'b10000:
        casez_tmp_128 = ldq_16_bits_uop_debug_pc;
      5'b10001:
        casez_tmp_128 = ldq_17_bits_uop_debug_pc;
      5'b10010:
        casez_tmp_128 = ldq_18_bits_uop_debug_pc;
      5'b10011:
        casez_tmp_128 = ldq_19_bits_uop_debug_pc;
      5'b10100:
        casez_tmp_128 = ldq_20_bits_uop_debug_pc;
      5'b10101:
        casez_tmp_128 = ldq_21_bits_uop_debug_pc;
      5'b10110:
        casez_tmp_128 = ldq_22_bits_uop_debug_pc;
      5'b10111:
        casez_tmp_128 = ldq_23_bits_uop_debug_pc;
      5'b11000:
        casez_tmp_128 = ldq_24_bits_uop_debug_pc;
      5'b11001:
        casez_tmp_128 = ldq_25_bits_uop_debug_pc;
      5'b11010:
        casez_tmp_128 = ldq_26_bits_uop_debug_pc;
      5'b11011:
        casez_tmp_128 = ldq_27_bits_uop_debug_pc;
      5'b11100:
        casez_tmp_128 = ldq_28_bits_uop_debug_pc;
      5'b11101:
        casez_tmp_128 = ldq_29_bits_uop_debug_pc;
      5'b11110:
        casez_tmp_128 = ldq_30_bits_uop_debug_pc;
      default:
        casez_tmp_128 = ldq_31_bits_uop_debug_pc;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_129;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_129 = ldq_0_bits_uop_iq_type;
      5'b00001:
        casez_tmp_129 = ldq_1_bits_uop_iq_type;
      5'b00010:
        casez_tmp_129 = ldq_2_bits_uop_iq_type;
      5'b00011:
        casez_tmp_129 = ldq_3_bits_uop_iq_type;
      5'b00100:
        casez_tmp_129 = ldq_4_bits_uop_iq_type;
      5'b00101:
        casez_tmp_129 = ldq_5_bits_uop_iq_type;
      5'b00110:
        casez_tmp_129 = ldq_6_bits_uop_iq_type;
      5'b00111:
        casez_tmp_129 = ldq_7_bits_uop_iq_type;
      5'b01000:
        casez_tmp_129 = ldq_8_bits_uop_iq_type;
      5'b01001:
        casez_tmp_129 = ldq_9_bits_uop_iq_type;
      5'b01010:
        casez_tmp_129 = ldq_10_bits_uop_iq_type;
      5'b01011:
        casez_tmp_129 = ldq_11_bits_uop_iq_type;
      5'b01100:
        casez_tmp_129 = ldq_12_bits_uop_iq_type;
      5'b01101:
        casez_tmp_129 = ldq_13_bits_uop_iq_type;
      5'b01110:
        casez_tmp_129 = ldq_14_bits_uop_iq_type;
      5'b01111:
        casez_tmp_129 = ldq_15_bits_uop_iq_type;
      5'b10000:
        casez_tmp_129 = ldq_16_bits_uop_iq_type;
      5'b10001:
        casez_tmp_129 = ldq_17_bits_uop_iq_type;
      5'b10010:
        casez_tmp_129 = ldq_18_bits_uop_iq_type;
      5'b10011:
        casez_tmp_129 = ldq_19_bits_uop_iq_type;
      5'b10100:
        casez_tmp_129 = ldq_20_bits_uop_iq_type;
      5'b10101:
        casez_tmp_129 = ldq_21_bits_uop_iq_type;
      5'b10110:
        casez_tmp_129 = ldq_22_bits_uop_iq_type;
      5'b10111:
        casez_tmp_129 = ldq_23_bits_uop_iq_type;
      5'b11000:
        casez_tmp_129 = ldq_24_bits_uop_iq_type;
      5'b11001:
        casez_tmp_129 = ldq_25_bits_uop_iq_type;
      5'b11010:
        casez_tmp_129 = ldq_26_bits_uop_iq_type;
      5'b11011:
        casez_tmp_129 = ldq_27_bits_uop_iq_type;
      5'b11100:
        casez_tmp_129 = ldq_28_bits_uop_iq_type;
      5'b11101:
        casez_tmp_129 = ldq_29_bits_uop_iq_type;
      5'b11110:
        casez_tmp_129 = ldq_30_bits_uop_iq_type;
      default:
        casez_tmp_129 = ldq_31_bits_uop_iq_type;
    endcase
  end // always @(*)
  reg  [9:0]  casez_tmp_130;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_130 = ldq_0_bits_uop_fu_code;
      5'b00001:
        casez_tmp_130 = ldq_1_bits_uop_fu_code;
      5'b00010:
        casez_tmp_130 = ldq_2_bits_uop_fu_code;
      5'b00011:
        casez_tmp_130 = ldq_3_bits_uop_fu_code;
      5'b00100:
        casez_tmp_130 = ldq_4_bits_uop_fu_code;
      5'b00101:
        casez_tmp_130 = ldq_5_bits_uop_fu_code;
      5'b00110:
        casez_tmp_130 = ldq_6_bits_uop_fu_code;
      5'b00111:
        casez_tmp_130 = ldq_7_bits_uop_fu_code;
      5'b01000:
        casez_tmp_130 = ldq_8_bits_uop_fu_code;
      5'b01001:
        casez_tmp_130 = ldq_9_bits_uop_fu_code;
      5'b01010:
        casez_tmp_130 = ldq_10_bits_uop_fu_code;
      5'b01011:
        casez_tmp_130 = ldq_11_bits_uop_fu_code;
      5'b01100:
        casez_tmp_130 = ldq_12_bits_uop_fu_code;
      5'b01101:
        casez_tmp_130 = ldq_13_bits_uop_fu_code;
      5'b01110:
        casez_tmp_130 = ldq_14_bits_uop_fu_code;
      5'b01111:
        casez_tmp_130 = ldq_15_bits_uop_fu_code;
      5'b10000:
        casez_tmp_130 = ldq_16_bits_uop_fu_code;
      5'b10001:
        casez_tmp_130 = ldq_17_bits_uop_fu_code;
      5'b10010:
        casez_tmp_130 = ldq_18_bits_uop_fu_code;
      5'b10011:
        casez_tmp_130 = ldq_19_bits_uop_fu_code;
      5'b10100:
        casez_tmp_130 = ldq_20_bits_uop_fu_code;
      5'b10101:
        casez_tmp_130 = ldq_21_bits_uop_fu_code;
      5'b10110:
        casez_tmp_130 = ldq_22_bits_uop_fu_code;
      5'b10111:
        casez_tmp_130 = ldq_23_bits_uop_fu_code;
      5'b11000:
        casez_tmp_130 = ldq_24_bits_uop_fu_code;
      5'b11001:
        casez_tmp_130 = ldq_25_bits_uop_fu_code;
      5'b11010:
        casez_tmp_130 = ldq_26_bits_uop_fu_code;
      5'b11011:
        casez_tmp_130 = ldq_27_bits_uop_fu_code;
      5'b11100:
        casez_tmp_130 = ldq_28_bits_uop_fu_code;
      5'b11101:
        casez_tmp_130 = ldq_29_bits_uop_fu_code;
      5'b11110:
        casez_tmp_130 = ldq_30_bits_uop_fu_code;
      default:
        casez_tmp_130 = ldq_31_bits_uop_fu_code;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_131;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_131 = ldq_0_bits_uop_ctrl_br_type;
      5'b00001:
        casez_tmp_131 = ldq_1_bits_uop_ctrl_br_type;
      5'b00010:
        casez_tmp_131 = ldq_2_bits_uop_ctrl_br_type;
      5'b00011:
        casez_tmp_131 = ldq_3_bits_uop_ctrl_br_type;
      5'b00100:
        casez_tmp_131 = ldq_4_bits_uop_ctrl_br_type;
      5'b00101:
        casez_tmp_131 = ldq_5_bits_uop_ctrl_br_type;
      5'b00110:
        casez_tmp_131 = ldq_6_bits_uop_ctrl_br_type;
      5'b00111:
        casez_tmp_131 = ldq_7_bits_uop_ctrl_br_type;
      5'b01000:
        casez_tmp_131 = ldq_8_bits_uop_ctrl_br_type;
      5'b01001:
        casez_tmp_131 = ldq_9_bits_uop_ctrl_br_type;
      5'b01010:
        casez_tmp_131 = ldq_10_bits_uop_ctrl_br_type;
      5'b01011:
        casez_tmp_131 = ldq_11_bits_uop_ctrl_br_type;
      5'b01100:
        casez_tmp_131 = ldq_12_bits_uop_ctrl_br_type;
      5'b01101:
        casez_tmp_131 = ldq_13_bits_uop_ctrl_br_type;
      5'b01110:
        casez_tmp_131 = ldq_14_bits_uop_ctrl_br_type;
      5'b01111:
        casez_tmp_131 = ldq_15_bits_uop_ctrl_br_type;
      5'b10000:
        casez_tmp_131 = ldq_16_bits_uop_ctrl_br_type;
      5'b10001:
        casez_tmp_131 = ldq_17_bits_uop_ctrl_br_type;
      5'b10010:
        casez_tmp_131 = ldq_18_bits_uop_ctrl_br_type;
      5'b10011:
        casez_tmp_131 = ldq_19_bits_uop_ctrl_br_type;
      5'b10100:
        casez_tmp_131 = ldq_20_bits_uop_ctrl_br_type;
      5'b10101:
        casez_tmp_131 = ldq_21_bits_uop_ctrl_br_type;
      5'b10110:
        casez_tmp_131 = ldq_22_bits_uop_ctrl_br_type;
      5'b10111:
        casez_tmp_131 = ldq_23_bits_uop_ctrl_br_type;
      5'b11000:
        casez_tmp_131 = ldq_24_bits_uop_ctrl_br_type;
      5'b11001:
        casez_tmp_131 = ldq_25_bits_uop_ctrl_br_type;
      5'b11010:
        casez_tmp_131 = ldq_26_bits_uop_ctrl_br_type;
      5'b11011:
        casez_tmp_131 = ldq_27_bits_uop_ctrl_br_type;
      5'b11100:
        casez_tmp_131 = ldq_28_bits_uop_ctrl_br_type;
      5'b11101:
        casez_tmp_131 = ldq_29_bits_uop_ctrl_br_type;
      5'b11110:
        casez_tmp_131 = ldq_30_bits_uop_ctrl_br_type;
      default:
        casez_tmp_131 = ldq_31_bits_uop_ctrl_br_type;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_132;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_132 = ldq_0_bits_uop_ctrl_op1_sel;
      5'b00001:
        casez_tmp_132 = ldq_1_bits_uop_ctrl_op1_sel;
      5'b00010:
        casez_tmp_132 = ldq_2_bits_uop_ctrl_op1_sel;
      5'b00011:
        casez_tmp_132 = ldq_3_bits_uop_ctrl_op1_sel;
      5'b00100:
        casez_tmp_132 = ldq_4_bits_uop_ctrl_op1_sel;
      5'b00101:
        casez_tmp_132 = ldq_5_bits_uop_ctrl_op1_sel;
      5'b00110:
        casez_tmp_132 = ldq_6_bits_uop_ctrl_op1_sel;
      5'b00111:
        casez_tmp_132 = ldq_7_bits_uop_ctrl_op1_sel;
      5'b01000:
        casez_tmp_132 = ldq_8_bits_uop_ctrl_op1_sel;
      5'b01001:
        casez_tmp_132 = ldq_9_bits_uop_ctrl_op1_sel;
      5'b01010:
        casez_tmp_132 = ldq_10_bits_uop_ctrl_op1_sel;
      5'b01011:
        casez_tmp_132 = ldq_11_bits_uop_ctrl_op1_sel;
      5'b01100:
        casez_tmp_132 = ldq_12_bits_uop_ctrl_op1_sel;
      5'b01101:
        casez_tmp_132 = ldq_13_bits_uop_ctrl_op1_sel;
      5'b01110:
        casez_tmp_132 = ldq_14_bits_uop_ctrl_op1_sel;
      5'b01111:
        casez_tmp_132 = ldq_15_bits_uop_ctrl_op1_sel;
      5'b10000:
        casez_tmp_132 = ldq_16_bits_uop_ctrl_op1_sel;
      5'b10001:
        casez_tmp_132 = ldq_17_bits_uop_ctrl_op1_sel;
      5'b10010:
        casez_tmp_132 = ldq_18_bits_uop_ctrl_op1_sel;
      5'b10011:
        casez_tmp_132 = ldq_19_bits_uop_ctrl_op1_sel;
      5'b10100:
        casez_tmp_132 = ldq_20_bits_uop_ctrl_op1_sel;
      5'b10101:
        casez_tmp_132 = ldq_21_bits_uop_ctrl_op1_sel;
      5'b10110:
        casez_tmp_132 = ldq_22_bits_uop_ctrl_op1_sel;
      5'b10111:
        casez_tmp_132 = ldq_23_bits_uop_ctrl_op1_sel;
      5'b11000:
        casez_tmp_132 = ldq_24_bits_uop_ctrl_op1_sel;
      5'b11001:
        casez_tmp_132 = ldq_25_bits_uop_ctrl_op1_sel;
      5'b11010:
        casez_tmp_132 = ldq_26_bits_uop_ctrl_op1_sel;
      5'b11011:
        casez_tmp_132 = ldq_27_bits_uop_ctrl_op1_sel;
      5'b11100:
        casez_tmp_132 = ldq_28_bits_uop_ctrl_op1_sel;
      5'b11101:
        casez_tmp_132 = ldq_29_bits_uop_ctrl_op1_sel;
      5'b11110:
        casez_tmp_132 = ldq_30_bits_uop_ctrl_op1_sel;
      default:
        casez_tmp_132 = ldq_31_bits_uop_ctrl_op1_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_133;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_133 = ldq_0_bits_uop_ctrl_op2_sel;
      5'b00001:
        casez_tmp_133 = ldq_1_bits_uop_ctrl_op2_sel;
      5'b00010:
        casez_tmp_133 = ldq_2_bits_uop_ctrl_op2_sel;
      5'b00011:
        casez_tmp_133 = ldq_3_bits_uop_ctrl_op2_sel;
      5'b00100:
        casez_tmp_133 = ldq_4_bits_uop_ctrl_op2_sel;
      5'b00101:
        casez_tmp_133 = ldq_5_bits_uop_ctrl_op2_sel;
      5'b00110:
        casez_tmp_133 = ldq_6_bits_uop_ctrl_op2_sel;
      5'b00111:
        casez_tmp_133 = ldq_7_bits_uop_ctrl_op2_sel;
      5'b01000:
        casez_tmp_133 = ldq_8_bits_uop_ctrl_op2_sel;
      5'b01001:
        casez_tmp_133 = ldq_9_bits_uop_ctrl_op2_sel;
      5'b01010:
        casez_tmp_133 = ldq_10_bits_uop_ctrl_op2_sel;
      5'b01011:
        casez_tmp_133 = ldq_11_bits_uop_ctrl_op2_sel;
      5'b01100:
        casez_tmp_133 = ldq_12_bits_uop_ctrl_op2_sel;
      5'b01101:
        casez_tmp_133 = ldq_13_bits_uop_ctrl_op2_sel;
      5'b01110:
        casez_tmp_133 = ldq_14_bits_uop_ctrl_op2_sel;
      5'b01111:
        casez_tmp_133 = ldq_15_bits_uop_ctrl_op2_sel;
      5'b10000:
        casez_tmp_133 = ldq_16_bits_uop_ctrl_op2_sel;
      5'b10001:
        casez_tmp_133 = ldq_17_bits_uop_ctrl_op2_sel;
      5'b10010:
        casez_tmp_133 = ldq_18_bits_uop_ctrl_op2_sel;
      5'b10011:
        casez_tmp_133 = ldq_19_bits_uop_ctrl_op2_sel;
      5'b10100:
        casez_tmp_133 = ldq_20_bits_uop_ctrl_op2_sel;
      5'b10101:
        casez_tmp_133 = ldq_21_bits_uop_ctrl_op2_sel;
      5'b10110:
        casez_tmp_133 = ldq_22_bits_uop_ctrl_op2_sel;
      5'b10111:
        casez_tmp_133 = ldq_23_bits_uop_ctrl_op2_sel;
      5'b11000:
        casez_tmp_133 = ldq_24_bits_uop_ctrl_op2_sel;
      5'b11001:
        casez_tmp_133 = ldq_25_bits_uop_ctrl_op2_sel;
      5'b11010:
        casez_tmp_133 = ldq_26_bits_uop_ctrl_op2_sel;
      5'b11011:
        casez_tmp_133 = ldq_27_bits_uop_ctrl_op2_sel;
      5'b11100:
        casez_tmp_133 = ldq_28_bits_uop_ctrl_op2_sel;
      5'b11101:
        casez_tmp_133 = ldq_29_bits_uop_ctrl_op2_sel;
      5'b11110:
        casez_tmp_133 = ldq_30_bits_uop_ctrl_op2_sel;
      default:
        casez_tmp_133 = ldq_31_bits_uop_ctrl_op2_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_134;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_134 = ldq_0_bits_uop_ctrl_imm_sel;
      5'b00001:
        casez_tmp_134 = ldq_1_bits_uop_ctrl_imm_sel;
      5'b00010:
        casez_tmp_134 = ldq_2_bits_uop_ctrl_imm_sel;
      5'b00011:
        casez_tmp_134 = ldq_3_bits_uop_ctrl_imm_sel;
      5'b00100:
        casez_tmp_134 = ldq_4_bits_uop_ctrl_imm_sel;
      5'b00101:
        casez_tmp_134 = ldq_5_bits_uop_ctrl_imm_sel;
      5'b00110:
        casez_tmp_134 = ldq_6_bits_uop_ctrl_imm_sel;
      5'b00111:
        casez_tmp_134 = ldq_7_bits_uop_ctrl_imm_sel;
      5'b01000:
        casez_tmp_134 = ldq_8_bits_uop_ctrl_imm_sel;
      5'b01001:
        casez_tmp_134 = ldq_9_bits_uop_ctrl_imm_sel;
      5'b01010:
        casez_tmp_134 = ldq_10_bits_uop_ctrl_imm_sel;
      5'b01011:
        casez_tmp_134 = ldq_11_bits_uop_ctrl_imm_sel;
      5'b01100:
        casez_tmp_134 = ldq_12_bits_uop_ctrl_imm_sel;
      5'b01101:
        casez_tmp_134 = ldq_13_bits_uop_ctrl_imm_sel;
      5'b01110:
        casez_tmp_134 = ldq_14_bits_uop_ctrl_imm_sel;
      5'b01111:
        casez_tmp_134 = ldq_15_bits_uop_ctrl_imm_sel;
      5'b10000:
        casez_tmp_134 = ldq_16_bits_uop_ctrl_imm_sel;
      5'b10001:
        casez_tmp_134 = ldq_17_bits_uop_ctrl_imm_sel;
      5'b10010:
        casez_tmp_134 = ldq_18_bits_uop_ctrl_imm_sel;
      5'b10011:
        casez_tmp_134 = ldq_19_bits_uop_ctrl_imm_sel;
      5'b10100:
        casez_tmp_134 = ldq_20_bits_uop_ctrl_imm_sel;
      5'b10101:
        casez_tmp_134 = ldq_21_bits_uop_ctrl_imm_sel;
      5'b10110:
        casez_tmp_134 = ldq_22_bits_uop_ctrl_imm_sel;
      5'b10111:
        casez_tmp_134 = ldq_23_bits_uop_ctrl_imm_sel;
      5'b11000:
        casez_tmp_134 = ldq_24_bits_uop_ctrl_imm_sel;
      5'b11001:
        casez_tmp_134 = ldq_25_bits_uop_ctrl_imm_sel;
      5'b11010:
        casez_tmp_134 = ldq_26_bits_uop_ctrl_imm_sel;
      5'b11011:
        casez_tmp_134 = ldq_27_bits_uop_ctrl_imm_sel;
      5'b11100:
        casez_tmp_134 = ldq_28_bits_uop_ctrl_imm_sel;
      5'b11101:
        casez_tmp_134 = ldq_29_bits_uop_ctrl_imm_sel;
      5'b11110:
        casez_tmp_134 = ldq_30_bits_uop_ctrl_imm_sel;
      default:
        casez_tmp_134 = ldq_31_bits_uop_ctrl_imm_sel;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_135;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_135 = ldq_0_bits_uop_ctrl_op_fcn;
      5'b00001:
        casez_tmp_135 = ldq_1_bits_uop_ctrl_op_fcn;
      5'b00010:
        casez_tmp_135 = ldq_2_bits_uop_ctrl_op_fcn;
      5'b00011:
        casez_tmp_135 = ldq_3_bits_uop_ctrl_op_fcn;
      5'b00100:
        casez_tmp_135 = ldq_4_bits_uop_ctrl_op_fcn;
      5'b00101:
        casez_tmp_135 = ldq_5_bits_uop_ctrl_op_fcn;
      5'b00110:
        casez_tmp_135 = ldq_6_bits_uop_ctrl_op_fcn;
      5'b00111:
        casez_tmp_135 = ldq_7_bits_uop_ctrl_op_fcn;
      5'b01000:
        casez_tmp_135 = ldq_8_bits_uop_ctrl_op_fcn;
      5'b01001:
        casez_tmp_135 = ldq_9_bits_uop_ctrl_op_fcn;
      5'b01010:
        casez_tmp_135 = ldq_10_bits_uop_ctrl_op_fcn;
      5'b01011:
        casez_tmp_135 = ldq_11_bits_uop_ctrl_op_fcn;
      5'b01100:
        casez_tmp_135 = ldq_12_bits_uop_ctrl_op_fcn;
      5'b01101:
        casez_tmp_135 = ldq_13_bits_uop_ctrl_op_fcn;
      5'b01110:
        casez_tmp_135 = ldq_14_bits_uop_ctrl_op_fcn;
      5'b01111:
        casez_tmp_135 = ldq_15_bits_uop_ctrl_op_fcn;
      5'b10000:
        casez_tmp_135 = ldq_16_bits_uop_ctrl_op_fcn;
      5'b10001:
        casez_tmp_135 = ldq_17_bits_uop_ctrl_op_fcn;
      5'b10010:
        casez_tmp_135 = ldq_18_bits_uop_ctrl_op_fcn;
      5'b10011:
        casez_tmp_135 = ldq_19_bits_uop_ctrl_op_fcn;
      5'b10100:
        casez_tmp_135 = ldq_20_bits_uop_ctrl_op_fcn;
      5'b10101:
        casez_tmp_135 = ldq_21_bits_uop_ctrl_op_fcn;
      5'b10110:
        casez_tmp_135 = ldq_22_bits_uop_ctrl_op_fcn;
      5'b10111:
        casez_tmp_135 = ldq_23_bits_uop_ctrl_op_fcn;
      5'b11000:
        casez_tmp_135 = ldq_24_bits_uop_ctrl_op_fcn;
      5'b11001:
        casez_tmp_135 = ldq_25_bits_uop_ctrl_op_fcn;
      5'b11010:
        casez_tmp_135 = ldq_26_bits_uop_ctrl_op_fcn;
      5'b11011:
        casez_tmp_135 = ldq_27_bits_uop_ctrl_op_fcn;
      5'b11100:
        casez_tmp_135 = ldq_28_bits_uop_ctrl_op_fcn;
      5'b11101:
        casez_tmp_135 = ldq_29_bits_uop_ctrl_op_fcn;
      5'b11110:
        casez_tmp_135 = ldq_30_bits_uop_ctrl_op_fcn;
      default:
        casez_tmp_135 = ldq_31_bits_uop_ctrl_op_fcn;
    endcase
  end // always @(*)
  reg         casez_tmp_136;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_136 = ldq_0_bits_uop_ctrl_fcn_dw;
      5'b00001:
        casez_tmp_136 = ldq_1_bits_uop_ctrl_fcn_dw;
      5'b00010:
        casez_tmp_136 = ldq_2_bits_uop_ctrl_fcn_dw;
      5'b00011:
        casez_tmp_136 = ldq_3_bits_uop_ctrl_fcn_dw;
      5'b00100:
        casez_tmp_136 = ldq_4_bits_uop_ctrl_fcn_dw;
      5'b00101:
        casez_tmp_136 = ldq_5_bits_uop_ctrl_fcn_dw;
      5'b00110:
        casez_tmp_136 = ldq_6_bits_uop_ctrl_fcn_dw;
      5'b00111:
        casez_tmp_136 = ldq_7_bits_uop_ctrl_fcn_dw;
      5'b01000:
        casez_tmp_136 = ldq_8_bits_uop_ctrl_fcn_dw;
      5'b01001:
        casez_tmp_136 = ldq_9_bits_uop_ctrl_fcn_dw;
      5'b01010:
        casez_tmp_136 = ldq_10_bits_uop_ctrl_fcn_dw;
      5'b01011:
        casez_tmp_136 = ldq_11_bits_uop_ctrl_fcn_dw;
      5'b01100:
        casez_tmp_136 = ldq_12_bits_uop_ctrl_fcn_dw;
      5'b01101:
        casez_tmp_136 = ldq_13_bits_uop_ctrl_fcn_dw;
      5'b01110:
        casez_tmp_136 = ldq_14_bits_uop_ctrl_fcn_dw;
      5'b01111:
        casez_tmp_136 = ldq_15_bits_uop_ctrl_fcn_dw;
      5'b10000:
        casez_tmp_136 = ldq_16_bits_uop_ctrl_fcn_dw;
      5'b10001:
        casez_tmp_136 = ldq_17_bits_uop_ctrl_fcn_dw;
      5'b10010:
        casez_tmp_136 = ldq_18_bits_uop_ctrl_fcn_dw;
      5'b10011:
        casez_tmp_136 = ldq_19_bits_uop_ctrl_fcn_dw;
      5'b10100:
        casez_tmp_136 = ldq_20_bits_uop_ctrl_fcn_dw;
      5'b10101:
        casez_tmp_136 = ldq_21_bits_uop_ctrl_fcn_dw;
      5'b10110:
        casez_tmp_136 = ldq_22_bits_uop_ctrl_fcn_dw;
      5'b10111:
        casez_tmp_136 = ldq_23_bits_uop_ctrl_fcn_dw;
      5'b11000:
        casez_tmp_136 = ldq_24_bits_uop_ctrl_fcn_dw;
      5'b11001:
        casez_tmp_136 = ldq_25_bits_uop_ctrl_fcn_dw;
      5'b11010:
        casez_tmp_136 = ldq_26_bits_uop_ctrl_fcn_dw;
      5'b11011:
        casez_tmp_136 = ldq_27_bits_uop_ctrl_fcn_dw;
      5'b11100:
        casez_tmp_136 = ldq_28_bits_uop_ctrl_fcn_dw;
      5'b11101:
        casez_tmp_136 = ldq_29_bits_uop_ctrl_fcn_dw;
      5'b11110:
        casez_tmp_136 = ldq_30_bits_uop_ctrl_fcn_dw;
      default:
        casez_tmp_136 = ldq_31_bits_uop_ctrl_fcn_dw;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_137;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_137 = ldq_0_bits_uop_ctrl_csr_cmd;
      5'b00001:
        casez_tmp_137 = ldq_1_bits_uop_ctrl_csr_cmd;
      5'b00010:
        casez_tmp_137 = ldq_2_bits_uop_ctrl_csr_cmd;
      5'b00011:
        casez_tmp_137 = ldq_3_bits_uop_ctrl_csr_cmd;
      5'b00100:
        casez_tmp_137 = ldq_4_bits_uop_ctrl_csr_cmd;
      5'b00101:
        casez_tmp_137 = ldq_5_bits_uop_ctrl_csr_cmd;
      5'b00110:
        casez_tmp_137 = ldq_6_bits_uop_ctrl_csr_cmd;
      5'b00111:
        casez_tmp_137 = ldq_7_bits_uop_ctrl_csr_cmd;
      5'b01000:
        casez_tmp_137 = ldq_8_bits_uop_ctrl_csr_cmd;
      5'b01001:
        casez_tmp_137 = ldq_9_bits_uop_ctrl_csr_cmd;
      5'b01010:
        casez_tmp_137 = ldq_10_bits_uop_ctrl_csr_cmd;
      5'b01011:
        casez_tmp_137 = ldq_11_bits_uop_ctrl_csr_cmd;
      5'b01100:
        casez_tmp_137 = ldq_12_bits_uop_ctrl_csr_cmd;
      5'b01101:
        casez_tmp_137 = ldq_13_bits_uop_ctrl_csr_cmd;
      5'b01110:
        casez_tmp_137 = ldq_14_bits_uop_ctrl_csr_cmd;
      5'b01111:
        casez_tmp_137 = ldq_15_bits_uop_ctrl_csr_cmd;
      5'b10000:
        casez_tmp_137 = ldq_16_bits_uop_ctrl_csr_cmd;
      5'b10001:
        casez_tmp_137 = ldq_17_bits_uop_ctrl_csr_cmd;
      5'b10010:
        casez_tmp_137 = ldq_18_bits_uop_ctrl_csr_cmd;
      5'b10011:
        casez_tmp_137 = ldq_19_bits_uop_ctrl_csr_cmd;
      5'b10100:
        casez_tmp_137 = ldq_20_bits_uop_ctrl_csr_cmd;
      5'b10101:
        casez_tmp_137 = ldq_21_bits_uop_ctrl_csr_cmd;
      5'b10110:
        casez_tmp_137 = ldq_22_bits_uop_ctrl_csr_cmd;
      5'b10111:
        casez_tmp_137 = ldq_23_bits_uop_ctrl_csr_cmd;
      5'b11000:
        casez_tmp_137 = ldq_24_bits_uop_ctrl_csr_cmd;
      5'b11001:
        casez_tmp_137 = ldq_25_bits_uop_ctrl_csr_cmd;
      5'b11010:
        casez_tmp_137 = ldq_26_bits_uop_ctrl_csr_cmd;
      5'b11011:
        casez_tmp_137 = ldq_27_bits_uop_ctrl_csr_cmd;
      5'b11100:
        casez_tmp_137 = ldq_28_bits_uop_ctrl_csr_cmd;
      5'b11101:
        casez_tmp_137 = ldq_29_bits_uop_ctrl_csr_cmd;
      5'b11110:
        casez_tmp_137 = ldq_30_bits_uop_ctrl_csr_cmd;
      default:
        casez_tmp_137 = ldq_31_bits_uop_ctrl_csr_cmd;
    endcase
  end // always @(*)
  reg         casez_tmp_138;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_138 = ldq_0_bits_uop_ctrl_is_load;
      5'b00001:
        casez_tmp_138 = ldq_1_bits_uop_ctrl_is_load;
      5'b00010:
        casez_tmp_138 = ldq_2_bits_uop_ctrl_is_load;
      5'b00011:
        casez_tmp_138 = ldq_3_bits_uop_ctrl_is_load;
      5'b00100:
        casez_tmp_138 = ldq_4_bits_uop_ctrl_is_load;
      5'b00101:
        casez_tmp_138 = ldq_5_bits_uop_ctrl_is_load;
      5'b00110:
        casez_tmp_138 = ldq_6_bits_uop_ctrl_is_load;
      5'b00111:
        casez_tmp_138 = ldq_7_bits_uop_ctrl_is_load;
      5'b01000:
        casez_tmp_138 = ldq_8_bits_uop_ctrl_is_load;
      5'b01001:
        casez_tmp_138 = ldq_9_bits_uop_ctrl_is_load;
      5'b01010:
        casez_tmp_138 = ldq_10_bits_uop_ctrl_is_load;
      5'b01011:
        casez_tmp_138 = ldq_11_bits_uop_ctrl_is_load;
      5'b01100:
        casez_tmp_138 = ldq_12_bits_uop_ctrl_is_load;
      5'b01101:
        casez_tmp_138 = ldq_13_bits_uop_ctrl_is_load;
      5'b01110:
        casez_tmp_138 = ldq_14_bits_uop_ctrl_is_load;
      5'b01111:
        casez_tmp_138 = ldq_15_bits_uop_ctrl_is_load;
      5'b10000:
        casez_tmp_138 = ldq_16_bits_uop_ctrl_is_load;
      5'b10001:
        casez_tmp_138 = ldq_17_bits_uop_ctrl_is_load;
      5'b10010:
        casez_tmp_138 = ldq_18_bits_uop_ctrl_is_load;
      5'b10011:
        casez_tmp_138 = ldq_19_bits_uop_ctrl_is_load;
      5'b10100:
        casez_tmp_138 = ldq_20_bits_uop_ctrl_is_load;
      5'b10101:
        casez_tmp_138 = ldq_21_bits_uop_ctrl_is_load;
      5'b10110:
        casez_tmp_138 = ldq_22_bits_uop_ctrl_is_load;
      5'b10111:
        casez_tmp_138 = ldq_23_bits_uop_ctrl_is_load;
      5'b11000:
        casez_tmp_138 = ldq_24_bits_uop_ctrl_is_load;
      5'b11001:
        casez_tmp_138 = ldq_25_bits_uop_ctrl_is_load;
      5'b11010:
        casez_tmp_138 = ldq_26_bits_uop_ctrl_is_load;
      5'b11011:
        casez_tmp_138 = ldq_27_bits_uop_ctrl_is_load;
      5'b11100:
        casez_tmp_138 = ldq_28_bits_uop_ctrl_is_load;
      5'b11101:
        casez_tmp_138 = ldq_29_bits_uop_ctrl_is_load;
      5'b11110:
        casez_tmp_138 = ldq_30_bits_uop_ctrl_is_load;
      default:
        casez_tmp_138 = ldq_31_bits_uop_ctrl_is_load;
    endcase
  end // always @(*)
  reg         casez_tmp_139;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_139 = ldq_0_bits_uop_ctrl_is_sta;
      5'b00001:
        casez_tmp_139 = ldq_1_bits_uop_ctrl_is_sta;
      5'b00010:
        casez_tmp_139 = ldq_2_bits_uop_ctrl_is_sta;
      5'b00011:
        casez_tmp_139 = ldq_3_bits_uop_ctrl_is_sta;
      5'b00100:
        casez_tmp_139 = ldq_4_bits_uop_ctrl_is_sta;
      5'b00101:
        casez_tmp_139 = ldq_5_bits_uop_ctrl_is_sta;
      5'b00110:
        casez_tmp_139 = ldq_6_bits_uop_ctrl_is_sta;
      5'b00111:
        casez_tmp_139 = ldq_7_bits_uop_ctrl_is_sta;
      5'b01000:
        casez_tmp_139 = ldq_8_bits_uop_ctrl_is_sta;
      5'b01001:
        casez_tmp_139 = ldq_9_bits_uop_ctrl_is_sta;
      5'b01010:
        casez_tmp_139 = ldq_10_bits_uop_ctrl_is_sta;
      5'b01011:
        casez_tmp_139 = ldq_11_bits_uop_ctrl_is_sta;
      5'b01100:
        casez_tmp_139 = ldq_12_bits_uop_ctrl_is_sta;
      5'b01101:
        casez_tmp_139 = ldq_13_bits_uop_ctrl_is_sta;
      5'b01110:
        casez_tmp_139 = ldq_14_bits_uop_ctrl_is_sta;
      5'b01111:
        casez_tmp_139 = ldq_15_bits_uop_ctrl_is_sta;
      5'b10000:
        casez_tmp_139 = ldq_16_bits_uop_ctrl_is_sta;
      5'b10001:
        casez_tmp_139 = ldq_17_bits_uop_ctrl_is_sta;
      5'b10010:
        casez_tmp_139 = ldq_18_bits_uop_ctrl_is_sta;
      5'b10011:
        casez_tmp_139 = ldq_19_bits_uop_ctrl_is_sta;
      5'b10100:
        casez_tmp_139 = ldq_20_bits_uop_ctrl_is_sta;
      5'b10101:
        casez_tmp_139 = ldq_21_bits_uop_ctrl_is_sta;
      5'b10110:
        casez_tmp_139 = ldq_22_bits_uop_ctrl_is_sta;
      5'b10111:
        casez_tmp_139 = ldq_23_bits_uop_ctrl_is_sta;
      5'b11000:
        casez_tmp_139 = ldq_24_bits_uop_ctrl_is_sta;
      5'b11001:
        casez_tmp_139 = ldq_25_bits_uop_ctrl_is_sta;
      5'b11010:
        casez_tmp_139 = ldq_26_bits_uop_ctrl_is_sta;
      5'b11011:
        casez_tmp_139 = ldq_27_bits_uop_ctrl_is_sta;
      5'b11100:
        casez_tmp_139 = ldq_28_bits_uop_ctrl_is_sta;
      5'b11101:
        casez_tmp_139 = ldq_29_bits_uop_ctrl_is_sta;
      5'b11110:
        casez_tmp_139 = ldq_30_bits_uop_ctrl_is_sta;
      default:
        casez_tmp_139 = ldq_31_bits_uop_ctrl_is_sta;
    endcase
  end // always @(*)
  reg         casez_tmp_140;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_140 = ldq_0_bits_uop_ctrl_is_std;
      5'b00001:
        casez_tmp_140 = ldq_1_bits_uop_ctrl_is_std;
      5'b00010:
        casez_tmp_140 = ldq_2_bits_uop_ctrl_is_std;
      5'b00011:
        casez_tmp_140 = ldq_3_bits_uop_ctrl_is_std;
      5'b00100:
        casez_tmp_140 = ldq_4_bits_uop_ctrl_is_std;
      5'b00101:
        casez_tmp_140 = ldq_5_bits_uop_ctrl_is_std;
      5'b00110:
        casez_tmp_140 = ldq_6_bits_uop_ctrl_is_std;
      5'b00111:
        casez_tmp_140 = ldq_7_bits_uop_ctrl_is_std;
      5'b01000:
        casez_tmp_140 = ldq_8_bits_uop_ctrl_is_std;
      5'b01001:
        casez_tmp_140 = ldq_9_bits_uop_ctrl_is_std;
      5'b01010:
        casez_tmp_140 = ldq_10_bits_uop_ctrl_is_std;
      5'b01011:
        casez_tmp_140 = ldq_11_bits_uop_ctrl_is_std;
      5'b01100:
        casez_tmp_140 = ldq_12_bits_uop_ctrl_is_std;
      5'b01101:
        casez_tmp_140 = ldq_13_bits_uop_ctrl_is_std;
      5'b01110:
        casez_tmp_140 = ldq_14_bits_uop_ctrl_is_std;
      5'b01111:
        casez_tmp_140 = ldq_15_bits_uop_ctrl_is_std;
      5'b10000:
        casez_tmp_140 = ldq_16_bits_uop_ctrl_is_std;
      5'b10001:
        casez_tmp_140 = ldq_17_bits_uop_ctrl_is_std;
      5'b10010:
        casez_tmp_140 = ldq_18_bits_uop_ctrl_is_std;
      5'b10011:
        casez_tmp_140 = ldq_19_bits_uop_ctrl_is_std;
      5'b10100:
        casez_tmp_140 = ldq_20_bits_uop_ctrl_is_std;
      5'b10101:
        casez_tmp_140 = ldq_21_bits_uop_ctrl_is_std;
      5'b10110:
        casez_tmp_140 = ldq_22_bits_uop_ctrl_is_std;
      5'b10111:
        casez_tmp_140 = ldq_23_bits_uop_ctrl_is_std;
      5'b11000:
        casez_tmp_140 = ldq_24_bits_uop_ctrl_is_std;
      5'b11001:
        casez_tmp_140 = ldq_25_bits_uop_ctrl_is_std;
      5'b11010:
        casez_tmp_140 = ldq_26_bits_uop_ctrl_is_std;
      5'b11011:
        casez_tmp_140 = ldq_27_bits_uop_ctrl_is_std;
      5'b11100:
        casez_tmp_140 = ldq_28_bits_uop_ctrl_is_std;
      5'b11101:
        casez_tmp_140 = ldq_29_bits_uop_ctrl_is_std;
      5'b11110:
        casez_tmp_140 = ldq_30_bits_uop_ctrl_is_std;
      default:
        casez_tmp_140 = ldq_31_bits_uop_ctrl_is_std;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_141;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_141 = ldq_0_bits_uop_iw_state;
      5'b00001:
        casez_tmp_141 = ldq_1_bits_uop_iw_state;
      5'b00010:
        casez_tmp_141 = ldq_2_bits_uop_iw_state;
      5'b00011:
        casez_tmp_141 = ldq_3_bits_uop_iw_state;
      5'b00100:
        casez_tmp_141 = ldq_4_bits_uop_iw_state;
      5'b00101:
        casez_tmp_141 = ldq_5_bits_uop_iw_state;
      5'b00110:
        casez_tmp_141 = ldq_6_bits_uop_iw_state;
      5'b00111:
        casez_tmp_141 = ldq_7_bits_uop_iw_state;
      5'b01000:
        casez_tmp_141 = ldq_8_bits_uop_iw_state;
      5'b01001:
        casez_tmp_141 = ldq_9_bits_uop_iw_state;
      5'b01010:
        casez_tmp_141 = ldq_10_bits_uop_iw_state;
      5'b01011:
        casez_tmp_141 = ldq_11_bits_uop_iw_state;
      5'b01100:
        casez_tmp_141 = ldq_12_bits_uop_iw_state;
      5'b01101:
        casez_tmp_141 = ldq_13_bits_uop_iw_state;
      5'b01110:
        casez_tmp_141 = ldq_14_bits_uop_iw_state;
      5'b01111:
        casez_tmp_141 = ldq_15_bits_uop_iw_state;
      5'b10000:
        casez_tmp_141 = ldq_16_bits_uop_iw_state;
      5'b10001:
        casez_tmp_141 = ldq_17_bits_uop_iw_state;
      5'b10010:
        casez_tmp_141 = ldq_18_bits_uop_iw_state;
      5'b10011:
        casez_tmp_141 = ldq_19_bits_uop_iw_state;
      5'b10100:
        casez_tmp_141 = ldq_20_bits_uop_iw_state;
      5'b10101:
        casez_tmp_141 = ldq_21_bits_uop_iw_state;
      5'b10110:
        casez_tmp_141 = ldq_22_bits_uop_iw_state;
      5'b10111:
        casez_tmp_141 = ldq_23_bits_uop_iw_state;
      5'b11000:
        casez_tmp_141 = ldq_24_bits_uop_iw_state;
      5'b11001:
        casez_tmp_141 = ldq_25_bits_uop_iw_state;
      5'b11010:
        casez_tmp_141 = ldq_26_bits_uop_iw_state;
      5'b11011:
        casez_tmp_141 = ldq_27_bits_uop_iw_state;
      5'b11100:
        casez_tmp_141 = ldq_28_bits_uop_iw_state;
      5'b11101:
        casez_tmp_141 = ldq_29_bits_uop_iw_state;
      5'b11110:
        casez_tmp_141 = ldq_30_bits_uop_iw_state;
      default:
        casez_tmp_141 = ldq_31_bits_uop_iw_state;
    endcase
  end // always @(*)
  reg         casez_tmp_142;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_142 = ldq_0_bits_uop_iw_p1_poisoned;
      5'b00001:
        casez_tmp_142 = ldq_1_bits_uop_iw_p1_poisoned;
      5'b00010:
        casez_tmp_142 = ldq_2_bits_uop_iw_p1_poisoned;
      5'b00011:
        casez_tmp_142 = ldq_3_bits_uop_iw_p1_poisoned;
      5'b00100:
        casez_tmp_142 = ldq_4_bits_uop_iw_p1_poisoned;
      5'b00101:
        casez_tmp_142 = ldq_5_bits_uop_iw_p1_poisoned;
      5'b00110:
        casez_tmp_142 = ldq_6_bits_uop_iw_p1_poisoned;
      5'b00111:
        casez_tmp_142 = ldq_7_bits_uop_iw_p1_poisoned;
      5'b01000:
        casez_tmp_142 = ldq_8_bits_uop_iw_p1_poisoned;
      5'b01001:
        casez_tmp_142 = ldq_9_bits_uop_iw_p1_poisoned;
      5'b01010:
        casez_tmp_142 = ldq_10_bits_uop_iw_p1_poisoned;
      5'b01011:
        casez_tmp_142 = ldq_11_bits_uop_iw_p1_poisoned;
      5'b01100:
        casez_tmp_142 = ldq_12_bits_uop_iw_p1_poisoned;
      5'b01101:
        casez_tmp_142 = ldq_13_bits_uop_iw_p1_poisoned;
      5'b01110:
        casez_tmp_142 = ldq_14_bits_uop_iw_p1_poisoned;
      5'b01111:
        casez_tmp_142 = ldq_15_bits_uop_iw_p1_poisoned;
      5'b10000:
        casez_tmp_142 = ldq_16_bits_uop_iw_p1_poisoned;
      5'b10001:
        casez_tmp_142 = ldq_17_bits_uop_iw_p1_poisoned;
      5'b10010:
        casez_tmp_142 = ldq_18_bits_uop_iw_p1_poisoned;
      5'b10011:
        casez_tmp_142 = ldq_19_bits_uop_iw_p1_poisoned;
      5'b10100:
        casez_tmp_142 = ldq_20_bits_uop_iw_p1_poisoned;
      5'b10101:
        casez_tmp_142 = ldq_21_bits_uop_iw_p1_poisoned;
      5'b10110:
        casez_tmp_142 = ldq_22_bits_uop_iw_p1_poisoned;
      5'b10111:
        casez_tmp_142 = ldq_23_bits_uop_iw_p1_poisoned;
      5'b11000:
        casez_tmp_142 = ldq_24_bits_uop_iw_p1_poisoned;
      5'b11001:
        casez_tmp_142 = ldq_25_bits_uop_iw_p1_poisoned;
      5'b11010:
        casez_tmp_142 = ldq_26_bits_uop_iw_p1_poisoned;
      5'b11011:
        casez_tmp_142 = ldq_27_bits_uop_iw_p1_poisoned;
      5'b11100:
        casez_tmp_142 = ldq_28_bits_uop_iw_p1_poisoned;
      5'b11101:
        casez_tmp_142 = ldq_29_bits_uop_iw_p1_poisoned;
      5'b11110:
        casez_tmp_142 = ldq_30_bits_uop_iw_p1_poisoned;
      default:
        casez_tmp_142 = ldq_31_bits_uop_iw_p1_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_143;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_143 = ldq_0_bits_uop_iw_p2_poisoned;
      5'b00001:
        casez_tmp_143 = ldq_1_bits_uop_iw_p2_poisoned;
      5'b00010:
        casez_tmp_143 = ldq_2_bits_uop_iw_p2_poisoned;
      5'b00011:
        casez_tmp_143 = ldq_3_bits_uop_iw_p2_poisoned;
      5'b00100:
        casez_tmp_143 = ldq_4_bits_uop_iw_p2_poisoned;
      5'b00101:
        casez_tmp_143 = ldq_5_bits_uop_iw_p2_poisoned;
      5'b00110:
        casez_tmp_143 = ldq_6_bits_uop_iw_p2_poisoned;
      5'b00111:
        casez_tmp_143 = ldq_7_bits_uop_iw_p2_poisoned;
      5'b01000:
        casez_tmp_143 = ldq_8_bits_uop_iw_p2_poisoned;
      5'b01001:
        casez_tmp_143 = ldq_9_bits_uop_iw_p2_poisoned;
      5'b01010:
        casez_tmp_143 = ldq_10_bits_uop_iw_p2_poisoned;
      5'b01011:
        casez_tmp_143 = ldq_11_bits_uop_iw_p2_poisoned;
      5'b01100:
        casez_tmp_143 = ldq_12_bits_uop_iw_p2_poisoned;
      5'b01101:
        casez_tmp_143 = ldq_13_bits_uop_iw_p2_poisoned;
      5'b01110:
        casez_tmp_143 = ldq_14_bits_uop_iw_p2_poisoned;
      5'b01111:
        casez_tmp_143 = ldq_15_bits_uop_iw_p2_poisoned;
      5'b10000:
        casez_tmp_143 = ldq_16_bits_uop_iw_p2_poisoned;
      5'b10001:
        casez_tmp_143 = ldq_17_bits_uop_iw_p2_poisoned;
      5'b10010:
        casez_tmp_143 = ldq_18_bits_uop_iw_p2_poisoned;
      5'b10011:
        casez_tmp_143 = ldq_19_bits_uop_iw_p2_poisoned;
      5'b10100:
        casez_tmp_143 = ldq_20_bits_uop_iw_p2_poisoned;
      5'b10101:
        casez_tmp_143 = ldq_21_bits_uop_iw_p2_poisoned;
      5'b10110:
        casez_tmp_143 = ldq_22_bits_uop_iw_p2_poisoned;
      5'b10111:
        casez_tmp_143 = ldq_23_bits_uop_iw_p2_poisoned;
      5'b11000:
        casez_tmp_143 = ldq_24_bits_uop_iw_p2_poisoned;
      5'b11001:
        casez_tmp_143 = ldq_25_bits_uop_iw_p2_poisoned;
      5'b11010:
        casez_tmp_143 = ldq_26_bits_uop_iw_p2_poisoned;
      5'b11011:
        casez_tmp_143 = ldq_27_bits_uop_iw_p2_poisoned;
      5'b11100:
        casez_tmp_143 = ldq_28_bits_uop_iw_p2_poisoned;
      5'b11101:
        casez_tmp_143 = ldq_29_bits_uop_iw_p2_poisoned;
      5'b11110:
        casez_tmp_143 = ldq_30_bits_uop_iw_p2_poisoned;
      default:
        casez_tmp_143 = ldq_31_bits_uop_iw_p2_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_144;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_144 = ldq_0_bits_uop_is_br;
      5'b00001:
        casez_tmp_144 = ldq_1_bits_uop_is_br;
      5'b00010:
        casez_tmp_144 = ldq_2_bits_uop_is_br;
      5'b00011:
        casez_tmp_144 = ldq_3_bits_uop_is_br;
      5'b00100:
        casez_tmp_144 = ldq_4_bits_uop_is_br;
      5'b00101:
        casez_tmp_144 = ldq_5_bits_uop_is_br;
      5'b00110:
        casez_tmp_144 = ldq_6_bits_uop_is_br;
      5'b00111:
        casez_tmp_144 = ldq_7_bits_uop_is_br;
      5'b01000:
        casez_tmp_144 = ldq_8_bits_uop_is_br;
      5'b01001:
        casez_tmp_144 = ldq_9_bits_uop_is_br;
      5'b01010:
        casez_tmp_144 = ldq_10_bits_uop_is_br;
      5'b01011:
        casez_tmp_144 = ldq_11_bits_uop_is_br;
      5'b01100:
        casez_tmp_144 = ldq_12_bits_uop_is_br;
      5'b01101:
        casez_tmp_144 = ldq_13_bits_uop_is_br;
      5'b01110:
        casez_tmp_144 = ldq_14_bits_uop_is_br;
      5'b01111:
        casez_tmp_144 = ldq_15_bits_uop_is_br;
      5'b10000:
        casez_tmp_144 = ldq_16_bits_uop_is_br;
      5'b10001:
        casez_tmp_144 = ldq_17_bits_uop_is_br;
      5'b10010:
        casez_tmp_144 = ldq_18_bits_uop_is_br;
      5'b10011:
        casez_tmp_144 = ldq_19_bits_uop_is_br;
      5'b10100:
        casez_tmp_144 = ldq_20_bits_uop_is_br;
      5'b10101:
        casez_tmp_144 = ldq_21_bits_uop_is_br;
      5'b10110:
        casez_tmp_144 = ldq_22_bits_uop_is_br;
      5'b10111:
        casez_tmp_144 = ldq_23_bits_uop_is_br;
      5'b11000:
        casez_tmp_144 = ldq_24_bits_uop_is_br;
      5'b11001:
        casez_tmp_144 = ldq_25_bits_uop_is_br;
      5'b11010:
        casez_tmp_144 = ldq_26_bits_uop_is_br;
      5'b11011:
        casez_tmp_144 = ldq_27_bits_uop_is_br;
      5'b11100:
        casez_tmp_144 = ldq_28_bits_uop_is_br;
      5'b11101:
        casez_tmp_144 = ldq_29_bits_uop_is_br;
      5'b11110:
        casez_tmp_144 = ldq_30_bits_uop_is_br;
      default:
        casez_tmp_144 = ldq_31_bits_uop_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_145;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_145 = ldq_0_bits_uop_is_jalr;
      5'b00001:
        casez_tmp_145 = ldq_1_bits_uop_is_jalr;
      5'b00010:
        casez_tmp_145 = ldq_2_bits_uop_is_jalr;
      5'b00011:
        casez_tmp_145 = ldq_3_bits_uop_is_jalr;
      5'b00100:
        casez_tmp_145 = ldq_4_bits_uop_is_jalr;
      5'b00101:
        casez_tmp_145 = ldq_5_bits_uop_is_jalr;
      5'b00110:
        casez_tmp_145 = ldq_6_bits_uop_is_jalr;
      5'b00111:
        casez_tmp_145 = ldq_7_bits_uop_is_jalr;
      5'b01000:
        casez_tmp_145 = ldq_8_bits_uop_is_jalr;
      5'b01001:
        casez_tmp_145 = ldq_9_bits_uop_is_jalr;
      5'b01010:
        casez_tmp_145 = ldq_10_bits_uop_is_jalr;
      5'b01011:
        casez_tmp_145 = ldq_11_bits_uop_is_jalr;
      5'b01100:
        casez_tmp_145 = ldq_12_bits_uop_is_jalr;
      5'b01101:
        casez_tmp_145 = ldq_13_bits_uop_is_jalr;
      5'b01110:
        casez_tmp_145 = ldq_14_bits_uop_is_jalr;
      5'b01111:
        casez_tmp_145 = ldq_15_bits_uop_is_jalr;
      5'b10000:
        casez_tmp_145 = ldq_16_bits_uop_is_jalr;
      5'b10001:
        casez_tmp_145 = ldq_17_bits_uop_is_jalr;
      5'b10010:
        casez_tmp_145 = ldq_18_bits_uop_is_jalr;
      5'b10011:
        casez_tmp_145 = ldq_19_bits_uop_is_jalr;
      5'b10100:
        casez_tmp_145 = ldq_20_bits_uop_is_jalr;
      5'b10101:
        casez_tmp_145 = ldq_21_bits_uop_is_jalr;
      5'b10110:
        casez_tmp_145 = ldq_22_bits_uop_is_jalr;
      5'b10111:
        casez_tmp_145 = ldq_23_bits_uop_is_jalr;
      5'b11000:
        casez_tmp_145 = ldq_24_bits_uop_is_jalr;
      5'b11001:
        casez_tmp_145 = ldq_25_bits_uop_is_jalr;
      5'b11010:
        casez_tmp_145 = ldq_26_bits_uop_is_jalr;
      5'b11011:
        casez_tmp_145 = ldq_27_bits_uop_is_jalr;
      5'b11100:
        casez_tmp_145 = ldq_28_bits_uop_is_jalr;
      5'b11101:
        casez_tmp_145 = ldq_29_bits_uop_is_jalr;
      5'b11110:
        casez_tmp_145 = ldq_30_bits_uop_is_jalr;
      default:
        casez_tmp_145 = ldq_31_bits_uop_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_146;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_146 = ldq_0_bits_uop_is_jal;
      5'b00001:
        casez_tmp_146 = ldq_1_bits_uop_is_jal;
      5'b00010:
        casez_tmp_146 = ldq_2_bits_uop_is_jal;
      5'b00011:
        casez_tmp_146 = ldq_3_bits_uop_is_jal;
      5'b00100:
        casez_tmp_146 = ldq_4_bits_uop_is_jal;
      5'b00101:
        casez_tmp_146 = ldq_5_bits_uop_is_jal;
      5'b00110:
        casez_tmp_146 = ldq_6_bits_uop_is_jal;
      5'b00111:
        casez_tmp_146 = ldq_7_bits_uop_is_jal;
      5'b01000:
        casez_tmp_146 = ldq_8_bits_uop_is_jal;
      5'b01001:
        casez_tmp_146 = ldq_9_bits_uop_is_jal;
      5'b01010:
        casez_tmp_146 = ldq_10_bits_uop_is_jal;
      5'b01011:
        casez_tmp_146 = ldq_11_bits_uop_is_jal;
      5'b01100:
        casez_tmp_146 = ldq_12_bits_uop_is_jal;
      5'b01101:
        casez_tmp_146 = ldq_13_bits_uop_is_jal;
      5'b01110:
        casez_tmp_146 = ldq_14_bits_uop_is_jal;
      5'b01111:
        casez_tmp_146 = ldq_15_bits_uop_is_jal;
      5'b10000:
        casez_tmp_146 = ldq_16_bits_uop_is_jal;
      5'b10001:
        casez_tmp_146 = ldq_17_bits_uop_is_jal;
      5'b10010:
        casez_tmp_146 = ldq_18_bits_uop_is_jal;
      5'b10011:
        casez_tmp_146 = ldq_19_bits_uop_is_jal;
      5'b10100:
        casez_tmp_146 = ldq_20_bits_uop_is_jal;
      5'b10101:
        casez_tmp_146 = ldq_21_bits_uop_is_jal;
      5'b10110:
        casez_tmp_146 = ldq_22_bits_uop_is_jal;
      5'b10111:
        casez_tmp_146 = ldq_23_bits_uop_is_jal;
      5'b11000:
        casez_tmp_146 = ldq_24_bits_uop_is_jal;
      5'b11001:
        casez_tmp_146 = ldq_25_bits_uop_is_jal;
      5'b11010:
        casez_tmp_146 = ldq_26_bits_uop_is_jal;
      5'b11011:
        casez_tmp_146 = ldq_27_bits_uop_is_jal;
      5'b11100:
        casez_tmp_146 = ldq_28_bits_uop_is_jal;
      5'b11101:
        casez_tmp_146 = ldq_29_bits_uop_is_jal;
      5'b11110:
        casez_tmp_146 = ldq_30_bits_uop_is_jal;
      default:
        casez_tmp_146 = ldq_31_bits_uop_is_jal;
    endcase
  end // always @(*)
  reg         casez_tmp_147;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_147 = ldq_0_bits_uop_is_sfb;
      5'b00001:
        casez_tmp_147 = ldq_1_bits_uop_is_sfb;
      5'b00010:
        casez_tmp_147 = ldq_2_bits_uop_is_sfb;
      5'b00011:
        casez_tmp_147 = ldq_3_bits_uop_is_sfb;
      5'b00100:
        casez_tmp_147 = ldq_4_bits_uop_is_sfb;
      5'b00101:
        casez_tmp_147 = ldq_5_bits_uop_is_sfb;
      5'b00110:
        casez_tmp_147 = ldq_6_bits_uop_is_sfb;
      5'b00111:
        casez_tmp_147 = ldq_7_bits_uop_is_sfb;
      5'b01000:
        casez_tmp_147 = ldq_8_bits_uop_is_sfb;
      5'b01001:
        casez_tmp_147 = ldq_9_bits_uop_is_sfb;
      5'b01010:
        casez_tmp_147 = ldq_10_bits_uop_is_sfb;
      5'b01011:
        casez_tmp_147 = ldq_11_bits_uop_is_sfb;
      5'b01100:
        casez_tmp_147 = ldq_12_bits_uop_is_sfb;
      5'b01101:
        casez_tmp_147 = ldq_13_bits_uop_is_sfb;
      5'b01110:
        casez_tmp_147 = ldq_14_bits_uop_is_sfb;
      5'b01111:
        casez_tmp_147 = ldq_15_bits_uop_is_sfb;
      5'b10000:
        casez_tmp_147 = ldq_16_bits_uop_is_sfb;
      5'b10001:
        casez_tmp_147 = ldq_17_bits_uop_is_sfb;
      5'b10010:
        casez_tmp_147 = ldq_18_bits_uop_is_sfb;
      5'b10011:
        casez_tmp_147 = ldq_19_bits_uop_is_sfb;
      5'b10100:
        casez_tmp_147 = ldq_20_bits_uop_is_sfb;
      5'b10101:
        casez_tmp_147 = ldq_21_bits_uop_is_sfb;
      5'b10110:
        casez_tmp_147 = ldq_22_bits_uop_is_sfb;
      5'b10111:
        casez_tmp_147 = ldq_23_bits_uop_is_sfb;
      5'b11000:
        casez_tmp_147 = ldq_24_bits_uop_is_sfb;
      5'b11001:
        casez_tmp_147 = ldq_25_bits_uop_is_sfb;
      5'b11010:
        casez_tmp_147 = ldq_26_bits_uop_is_sfb;
      5'b11011:
        casez_tmp_147 = ldq_27_bits_uop_is_sfb;
      5'b11100:
        casez_tmp_147 = ldq_28_bits_uop_is_sfb;
      5'b11101:
        casez_tmp_147 = ldq_29_bits_uop_is_sfb;
      5'b11110:
        casez_tmp_147 = ldq_30_bits_uop_is_sfb;
      default:
        casez_tmp_147 = ldq_31_bits_uop_is_sfb;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_148;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_148 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_148 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_148 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_148 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_148 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_148 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_148 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_148 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_148 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_148 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_148 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_148 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_148 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_148 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_148 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_148 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_148 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_148 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_148 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_148 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_148 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_148 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_148 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_148 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_148 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_148 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_148 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_148 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_148 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_148 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_148 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_148 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_149;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_149 = ldq_0_bits_uop_br_tag;
      5'b00001:
        casez_tmp_149 = ldq_1_bits_uop_br_tag;
      5'b00010:
        casez_tmp_149 = ldq_2_bits_uop_br_tag;
      5'b00011:
        casez_tmp_149 = ldq_3_bits_uop_br_tag;
      5'b00100:
        casez_tmp_149 = ldq_4_bits_uop_br_tag;
      5'b00101:
        casez_tmp_149 = ldq_5_bits_uop_br_tag;
      5'b00110:
        casez_tmp_149 = ldq_6_bits_uop_br_tag;
      5'b00111:
        casez_tmp_149 = ldq_7_bits_uop_br_tag;
      5'b01000:
        casez_tmp_149 = ldq_8_bits_uop_br_tag;
      5'b01001:
        casez_tmp_149 = ldq_9_bits_uop_br_tag;
      5'b01010:
        casez_tmp_149 = ldq_10_bits_uop_br_tag;
      5'b01011:
        casez_tmp_149 = ldq_11_bits_uop_br_tag;
      5'b01100:
        casez_tmp_149 = ldq_12_bits_uop_br_tag;
      5'b01101:
        casez_tmp_149 = ldq_13_bits_uop_br_tag;
      5'b01110:
        casez_tmp_149 = ldq_14_bits_uop_br_tag;
      5'b01111:
        casez_tmp_149 = ldq_15_bits_uop_br_tag;
      5'b10000:
        casez_tmp_149 = ldq_16_bits_uop_br_tag;
      5'b10001:
        casez_tmp_149 = ldq_17_bits_uop_br_tag;
      5'b10010:
        casez_tmp_149 = ldq_18_bits_uop_br_tag;
      5'b10011:
        casez_tmp_149 = ldq_19_bits_uop_br_tag;
      5'b10100:
        casez_tmp_149 = ldq_20_bits_uop_br_tag;
      5'b10101:
        casez_tmp_149 = ldq_21_bits_uop_br_tag;
      5'b10110:
        casez_tmp_149 = ldq_22_bits_uop_br_tag;
      5'b10111:
        casez_tmp_149 = ldq_23_bits_uop_br_tag;
      5'b11000:
        casez_tmp_149 = ldq_24_bits_uop_br_tag;
      5'b11001:
        casez_tmp_149 = ldq_25_bits_uop_br_tag;
      5'b11010:
        casez_tmp_149 = ldq_26_bits_uop_br_tag;
      5'b11011:
        casez_tmp_149 = ldq_27_bits_uop_br_tag;
      5'b11100:
        casez_tmp_149 = ldq_28_bits_uop_br_tag;
      5'b11101:
        casez_tmp_149 = ldq_29_bits_uop_br_tag;
      5'b11110:
        casez_tmp_149 = ldq_30_bits_uop_br_tag;
      default:
        casez_tmp_149 = ldq_31_bits_uop_br_tag;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_150;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_150 = ldq_0_bits_uop_ftq_idx;
      5'b00001:
        casez_tmp_150 = ldq_1_bits_uop_ftq_idx;
      5'b00010:
        casez_tmp_150 = ldq_2_bits_uop_ftq_idx;
      5'b00011:
        casez_tmp_150 = ldq_3_bits_uop_ftq_idx;
      5'b00100:
        casez_tmp_150 = ldq_4_bits_uop_ftq_idx;
      5'b00101:
        casez_tmp_150 = ldq_5_bits_uop_ftq_idx;
      5'b00110:
        casez_tmp_150 = ldq_6_bits_uop_ftq_idx;
      5'b00111:
        casez_tmp_150 = ldq_7_bits_uop_ftq_idx;
      5'b01000:
        casez_tmp_150 = ldq_8_bits_uop_ftq_idx;
      5'b01001:
        casez_tmp_150 = ldq_9_bits_uop_ftq_idx;
      5'b01010:
        casez_tmp_150 = ldq_10_bits_uop_ftq_idx;
      5'b01011:
        casez_tmp_150 = ldq_11_bits_uop_ftq_idx;
      5'b01100:
        casez_tmp_150 = ldq_12_bits_uop_ftq_idx;
      5'b01101:
        casez_tmp_150 = ldq_13_bits_uop_ftq_idx;
      5'b01110:
        casez_tmp_150 = ldq_14_bits_uop_ftq_idx;
      5'b01111:
        casez_tmp_150 = ldq_15_bits_uop_ftq_idx;
      5'b10000:
        casez_tmp_150 = ldq_16_bits_uop_ftq_idx;
      5'b10001:
        casez_tmp_150 = ldq_17_bits_uop_ftq_idx;
      5'b10010:
        casez_tmp_150 = ldq_18_bits_uop_ftq_idx;
      5'b10011:
        casez_tmp_150 = ldq_19_bits_uop_ftq_idx;
      5'b10100:
        casez_tmp_150 = ldq_20_bits_uop_ftq_idx;
      5'b10101:
        casez_tmp_150 = ldq_21_bits_uop_ftq_idx;
      5'b10110:
        casez_tmp_150 = ldq_22_bits_uop_ftq_idx;
      5'b10111:
        casez_tmp_150 = ldq_23_bits_uop_ftq_idx;
      5'b11000:
        casez_tmp_150 = ldq_24_bits_uop_ftq_idx;
      5'b11001:
        casez_tmp_150 = ldq_25_bits_uop_ftq_idx;
      5'b11010:
        casez_tmp_150 = ldq_26_bits_uop_ftq_idx;
      5'b11011:
        casez_tmp_150 = ldq_27_bits_uop_ftq_idx;
      5'b11100:
        casez_tmp_150 = ldq_28_bits_uop_ftq_idx;
      5'b11101:
        casez_tmp_150 = ldq_29_bits_uop_ftq_idx;
      5'b11110:
        casez_tmp_150 = ldq_30_bits_uop_ftq_idx;
      default:
        casez_tmp_150 = ldq_31_bits_uop_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_151;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_151 = ldq_0_bits_uop_edge_inst;
      5'b00001:
        casez_tmp_151 = ldq_1_bits_uop_edge_inst;
      5'b00010:
        casez_tmp_151 = ldq_2_bits_uop_edge_inst;
      5'b00011:
        casez_tmp_151 = ldq_3_bits_uop_edge_inst;
      5'b00100:
        casez_tmp_151 = ldq_4_bits_uop_edge_inst;
      5'b00101:
        casez_tmp_151 = ldq_5_bits_uop_edge_inst;
      5'b00110:
        casez_tmp_151 = ldq_6_bits_uop_edge_inst;
      5'b00111:
        casez_tmp_151 = ldq_7_bits_uop_edge_inst;
      5'b01000:
        casez_tmp_151 = ldq_8_bits_uop_edge_inst;
      5'b01001:
        casez_tmp_151 = ldq_9_bits_uop_edge_inst;
      5'b01010:
        casez_tmp_151 = ldq_10_bits_uop_edge_inst;
      5'b01011:
        casez_tmp_151 = ldq_11_bits_uop_edge_inst;
      5'b01100:
        casez_tmp_151 = ldq_12_bits_uop_edge_inst;
      5'b01101:
        casez_tmp_151 = ldq_13_bits_uop_edge_inst;
      5'b01110:
        casez_tmp_151 = ldq_14_bits_uop_edge_inst;
      5'b01111:
        casez_tmp_151 = ldq_15_bits_uop_edge_inst;
      5'b10000:
        casez_tmp_151 = ldq_16_bits_uop_edge_inst;
      5'b10001:
        casez_tmp_151 = ldq_17_bits_uop_edge_inst;
      5'b10010:
        casez_tmp_151 = ldq_18_bits_uop_edge_inst;
      5'b10011:
        casez_tmp_151 = ldq_19_bits_uop_edge_inst;
      5'b10100:
        casez_tmp_151 = ldq_20_bits_uop_edge_inst;
      5'b10101:
        casez_tmp_151 = ldq_21_bits_uop_edge_inst;
      5'b10110:
        casez_tmp_151 = ldq_22_bits_uop_edge_inst;
      5'b10111:
        casez_tmp_151 = ldq_23_bits_uop_edge_inst;
      5'b11000:
        casez_tmp_151 = ldq_24_bits_uop_edge_inst;
      5'b11001:
        casez_tmp_151 = ldq_25_bits_uop_edge_inst;
      5'b11010:
        casez_tmp_151 = ldq_26_bits_uop_edge_inst;
      5'b11011:
        casez_tmp_151 = ldq_27_bits_uop_edge_inst;
      5'b11100:
        casez_tmp_151 = ldq_28_bits_uop_edge_inst;
      5'b11101:
        casez_tmp_151 = ldq_29_bits_uop_edge_inst;
      5'b11110:
        casez_tmp_151 = ldq_30_bits_uop_edge_inst;
      default:
        casez_tmp_151 = ldq_31_bits_uop_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_152;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_152 = ldq_0_bits_uop_pc_lob;
      5'b00001:
        casez_tmp_152 = ldq_1_bits_uop_pc_lob;
      5'b00010:
        casez_tmp_152 = ldq_2_bits_uop_pc_lob;
      5'b00011:
        casez_tmp_152 = ldq_3_bits_uop_pc_lob;
      5'b00100:
        casez_tmp_152 = ldq_4_bits_uop_pc_lob;
      5'b00101:
        casez_tmp_152 = ldq_5_bits_uop_pc_lob;
      5'b00110:
        casez_tmp_152 = ldq_6_bits_uop_pc_lob;
      5'b00111:
        casez_tmp_152 = ldq_7_bits_uop_pc_lob;
      5'b01000:
        casez_tmp_152 = ldq_8_bits_uop_pc_lob;
      5'b01001:
        casez_tmp_152 = ldq_9_bits_uop_pc_lob;
      5'b01010:
        casez_tmp_152 = ldq_10_bits_uop_pc_lob;
      5'b01011:
        casez_tmp_152 = ldq_11_bits_uop_pc_lob;
      5'b01100:
        casez_tmp_152 = ldq_12_bits_uop_pc_lob;
      5'b01101:
        casez_tmp_152 = ldq_13_bits_uop_pc_lob;
      5'b01110:
        casez_tmp_152 = ldq_14_bits_uop_pc_lob;
      5'b01111:
        casez_tmp_152 = ldq_15_bits_uop_pc_lob;
      5'b10000:
        casez_tmp_152 = ldq_16_bits_uop_pc_lob;
      5'b10001:
        casez_tmp_152 = ldq_17_bits_uop_pc_lob;
      5'b10010:
        casez_tmp_152 = ldq_18_bits_uop_pc_lob;
      5'b10011:
        casez_tmp_152 = ldq_19_bits_uop_pc_lob;
      5'b10100:
        casez_tmp_152 = ldq_20_bits_uop_pc_lob;
      5'b10101:
        casez_tmp_152 = ldq_21_bits_uop_pc_lob;
      5'b10110:
        casez_tmp_152 = ldq_22_bits_uop_pc_lob;
      5'b10111:
        casez_tmp_152 = ldq_23_bits_uop_pc_lob;
      5'b11000:
        casez_tmp_152 = ldq_24_bits_uop_pc_lob;
      5'b11001:
        casez_tmp_152 = ldq_25_bits_uop_pc_lob;
      5'b11010:
        casez_tmp_152 = ldq_26_bits_uop_pc_lob;
      5'b11011:
        casez_tmp_152 = ldq_27_bits_uop_pc_lob;
      5'b11100:
        casez_tmp_152 = ldq_28_bits_uop_pc_lob;
      5'b11101:
        casez_tmp_152 = ldq_29_bits_uop_pc_lob;
      5'b11110:
        casez_tmp_152 = ldq_30_bits_uop_pc_lob;
      default:
        casez_tmp_152 = ldq_31_bits_uop_pc_lob;
    endcase
  end // always @(*)
  reg         casez_tmp_153;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_153 = ldq_0_bits_uop_taken;
      5'b00001:
        casez_tmp_153 = ldq_1_bits_uop_taken;
      5'b00010:
        casez_tmp_153 = ldq_2_bits_uop_taken;
      5'b00011:
        casez_tmp_153 = ldq_3_bits_uop_taken;
      5'b00100:
        casez_tmp_153 = ldq_4_bits_uop_taken;
      5'b00101:
        casez_tmp_153 = ldq_5_bits_uop_taken;
      5'b00110:
        casez_tmp_153 = ldq_6_bits_uop_taken;
      5'b00111:
        casez_tmp_153 = ldq_7_bits_uop_taken;
      5'b01000:
        casez_tmp_153 = ldq_8_bits_uop_taken;
      5'b01001:
        casez_tmp_153 = ldq_9_bits_uop_taken;
      5'b01010:
        casez_tmp_153 = ldq_10_bits_uop_taken;
      5'b01011:
        casez_tmp_153 = ldq_11_bits_uop_taken;
      5'b01100:
        casez_tmp_153 = ldq_12_bits_uop_taken;
      5'b01101:
        casez_tmp_153 = ldq_13_bits_uop_taken;
      5'b01110:
        casez_tmp_153 = ldq_14_bits_uop_taken;
      5'b01111:
        casez_tmp_153 = ldq_15_bits_uop_taken;
      5'b10000:
        casez_tmp_153 = ldq_16_bits_uop_taken;
      5'b10001:
        casez_tmp_153 = ldq_17_bits_uop_taken;
      5'b10010:
        casez_tmp_153 = ldq_18_bits_uop_taken;
      5'b10011:
        casez_tmp_153 = ldq_19_bits_uop_taken;
      5'b10100:
        casez_tmp_153 = ldq_20_bits_uop_taken;
      5'b10101:
        casez_tmp_153 = ldq_21_bits_uop_taken;
      5'b10110:
        casez_tmp_153 = ldq_22_bits_uop_taken;
      5'b10111:
        casez_tmp_153 = ldq_23_bits_uop_taken;
      5'b11000:
        casez_tmp_153 = ldq_24_bits_uop_taken;
      5'b11001:
        casez_tmp_153 = ldq_25_bits_uop_taken;
      5'b11010:
        casez_tmp_153 = ldq_26_bits_uop_taken;
      5'b11011:
        casez_tmp_153 = ldq_27_bits_uop_taken;
      5'b11100:
        casez_tmp_153 = ldq_28_bits_uop_taken;
      5'b11101:
        casez_tmp_153 = ldq_29_bits_uop_taken;
      5'b11110:
        casez_tmp_153 = ldq_30_bits_uop_taken;
      default:
        casez_tmp_153 = ldq_31_bits_uop_taken;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_154;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_154 = ldq_0_bits_uop_imm_packed;
      5'b00001:
        casez_tmp_154 = ldq_1_bits_uop_imm_packed;
      5'b00010:
        casez_tmp_154 = ldq_2_bits_uop_imm_packed;
      5'b00011:
        casez_tmp_154 = ldq_3_bits_uop_imm_packed;
      5'b00100:
        casez_tmp_154 = ldq_4_bits_uop_imm_packed;
      5'b00101:
        casez_tmp_154 = ldq_5_bits_uop_imm_packed;
      5'b00110:
        casez_tmp_154 = ldq_6_bits_uop_imm_packed;
      5'b00111:
        casez_tmp_154 = ldq_7_bits_uop_imm_packed;
      5'b01000:
        casez_tmp_154 = ldq_8_bits_uop_imm_packed;
      5'b01001:
        casez_tmp_154 = ldq_9_bits_uop_imm_packed;
      5'b01010:
        casez_tmp_154 = ldq_10_bits_uop_imm_packed;
      5'b01011:
        casez_tmp_154 = ldq_11_bits_uop_imm_packed;
      5'b01100:
        casez_tmp_154 = ldq_12_bits_uop_imm_packed;
      5'b01101:
        casez_tmp_154 = ldq_13_bits_uop_imm_packed;
      5'b01110:
        casez_tmp_154 = ldq_14_bits_uop_imm_packed;
      5'b01111:
        casez_tmp_154 = ldq_15_bits_uop_imm_packed;
      5'b10000:
        casez_tmp_154 = ldq_16_bits_uop_imm_packed;
      5'b10001:
        casez_tmp_154 = ldq_17_bits_uop_imm_packed;
      5'b10010:
        casez_tmp_154 = ldq_18_bits_uop_imm_packed;
      5'b10011:
        casez_tmp_154 = ldq_19_bits_uop_imm_packed;
      5'b10100:
        casez_tmp_154 = ldq_20_bits_uop_imm_packed;
      5'b10101:
        casez_tmp_154 = ldq_21_bits_uop_imm_packed;
      5'b10110:
        casez_tmp_154 = ldq_22_bits_uop_imm_packed;
      5'b10111:
        casez_tmp_154 = ldq_23_bits_uop_imm_packed;
      5'b11000:
        casez_tmp_154 = ldq_24_bits_uop_imm_packed;
      5'b11001:
        casez_tmp_154 = ldq_25_bits_uop_imm_packed;
      5'b11010:
        casez_tmp_154 = ldq_26_bits_uop_imm_packed;
      5'b11011:
        casez_tmp_154 = ldq_27_bits_uop_imm_packed;
      5'b11100:
        casez_tmp_154 = ldq_28_bits_uop_imm_packed;
      5'b11101:
        casez_tmp_154 = ldq_29_bits_uop_imm_packed;
      5'b11110:
        casez_tmp_154 = ldq_30_bits_uop_imm_packed;
      default:
        casez_tmp_154 = ldq_31_bits_uop_imm_packed;
    endcase
  end // always @(*)
  reg  [11:0] casez_tmp_155;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_155 = ldq_0_bits_uop_csr_addr;
      5'b00001:
        casez_tmp_155 = ldq_1_bits_uop_csr_addr;
      5'b00010:
        casez_tmp_155 = ldq_2_bits_uop_csr_addr;
      5'b00011:
        casez_tmp_155 = ldq_3_bits_uop_csr_addr;
      5'b00100:
        casez_tmp_155 = ldq_4_bits_uop_csr_addr;
      5'b00101:
        casez_tmp_155 = ldq_5_bits_uop_csr_addr;
      5'b00110:
        casez_tmp_155 = ldq_6_bits_uop_csr_addr;
      5'b00111:
        casez_tmp_155 = ldq_7_bits_uop_csr_addr;
      5'b01000:
        casez_tmp_155 = ldq_8_bits_uop_csr_addr;
      5'b01001:
        casez_tmp_155 = ldq_9_bits_uop_csr_addr;
      5'b01010:
        casez_tmp_155 = ldq_10_bits_uop_csr_addr;
      5'b01011:
        casez_tmp_155 = ldq_11_bits_uop_csr_addr;
      5'b01100:
        casez_tmp_155 = ldq_12_bits_uop_csr_addr;
      5'b01101:
        casez_tmp_155 = ldq_13_bits_uop_csr_addr;
      5'b01110:
        casez_tmp_155 = ldq_14_bits_uop_csr_addr;
      5'b01111:
        casez_tmp_155 = ldq_15_bits_uop_csr_addr;
      5'b10000:
        casez_tmp_155 = ldq_16_bits_uop_csr_addr;
      5'b10001:
        casez_tmp_155 = ldq_17_bits_uop_csr_addr;
      5'b10010:
        casez_tmp_155 = ldq_18_bits_uop_csr_addr;
      5'b10011:
        casez_tmp_155 = ldq_19_bits_uop_csr_addr;
      5'b10100:
        casez_tmp_155 = ldq_20_bits_uop_csr_addr;
      5'b10101:
        casez_tmp_155 = ldq_21_bits_uop_csr_addr;
      5'b10110:
        casez_tmp_155 = ldq_22_bits_uop_csr_addr;
      5'b10111:
        casez_tmp_155 = ldq_23_bits_uop_csr_addr;
      5'b11000:
        casez_tmp_155 = ldq_24_bits_uop_csr_addr;
      5'b11001:
        casez_tmp_155 = ldq_25_bits_uop_csr_addr;
      5'b11010:
        casez_tmp_155 = ldq_26_bits_uop_csr_addr;
      5'b11011:
        casez_tmp_155 = ldq_27_bits_uop_csr_addr;
      5'b11100:
        casez_tmp_155 = ldq_28_bits_uop_csr_addr;
      5'b11101:
        casez_tmp_155 = ldq_29_bits_uop_csr_addr;
      5'b11110:
        casez_tmp_155 = ldq_30_bits_uop_csr_addr;
      default:
        casez_tmp_155 = ldq_31_bits_uop_csr_addr;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_156;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_156 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_156 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_156 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_156 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_156 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_156 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_156 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_156 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_156 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_156 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_156 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_156 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_156 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_156 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_156 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_156 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_156 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_156 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_156 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_156 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_156 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_156 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_156 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_156 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_156 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_156 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_156 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_156 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_156 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_156 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_156 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_156 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_157;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_157 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_157 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_157 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_157 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_157 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_157 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_157 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_157 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_157 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_157 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_157 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_157 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_157 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_157 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_157 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_157 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_157 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_157 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_157 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_157 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_157 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_157 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_157 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_157 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_157 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_157 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_157 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_157 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_157 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_157 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_157 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_157 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_158;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_158 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_158 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_158 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_158 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_158 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_158 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_158 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_158 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_158 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_158 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_158 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_158 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_158 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_158 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_158 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_158 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_158 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_158 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_158 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_158 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_158 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_158 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_158 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_158 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_158 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_158 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_158 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_158 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_158 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_158 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_158 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_158 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_159;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_159 = ldq_0_bits_uop_rxq_idx;
      5'b00001:
        casez_tmp_159 = ldq_1_bits_uop_rxq_idx;
      5'b00010:
        casez_tmp_159 = ldq_2_bits_uop_rxq_idx;
      5'b00011:
        casez_tmp_159 = ldq_3_bits_uop_rxq_idx;
      5'b00100:
        casez_tmp_159 = ldq_4_bits_uop_rxq_idx;
      5'b00101:
        casez_tmp_159 = ldq_5_bits_uop_rxq_idx;
      5'b00110:
        casez_tmp_159 = ldq_6_bits_uop_rxq_idx;
      5'b00111:
        casez_tmp_159 = ldq_7_bits_uop_rxq_idx;
      5'b01000:
        casez_tmp_159 = ldq_8_bits_uop_rxq_idx;
      5'b01001:
        casez_tmp_159 = ldq_9_bits_uop_rxq_idx;
      5'b01010:
        casez_tmp_159 = ldq_10_bits_uop_rxq_idx;
      5'b01011:
        casez_tmp_159 = ldq_11_bits_uop_rxq_idx;
      5'b01100:
        casez_tmp_159 = ldq_12_bits_uop_rxq_idx;
      5'b01101:
        casez_tmp_159 = ldq_13_bits_uop_rxq_idx;
      5'b01110:
        casez_tmp_159 = ldq_14_bits_uop_rxq_idx;
      5'b01111:
        casez_tmp_159 = ldq_15_bits_uop_rxq_idx;
      5'b10000:
        casez_tmp_159 = ldq_16_bits_uop_rxq_idx;
      5'b10001:
        casez_tmp_159 = ldq_17_bits_uop_rxq_idx;
      5'b10010:
        casez_tmp_159 = ldq_18_bits_uop_rxq_idx;
      5'b10011:
        casez_tmp_159 = ldq_19_bits_uop_rxq_idx;
      5'b10100:
        casez_tmp_159 = ldq_20_bits_uop_rxq_idx;
      5'b10101:
        casez_tmp_159 = ldq_21_bits_uop_rxq_idx;
      5'b10110:
        casez_tmp_159 = ldq_22_bits_uop_rxq_idx;
      5'b10111:
        casez_tmp_159 = ldq_23_bits_uop_rxq_idx;
      5'b11000:
        casez_tmp_159 = ldq_24_bits_uop_rxq_idx;
      5'b11001:
        casez_tmp_159 = ldq_25_bits_uop_rxq_idx;
      5'b11010:
        casez_tmp_159 = ldq_26_bits_uop_rxq_idx;
      5'b11011:
        casez_tmp_159 = ldq_27_bits_uop_rxq_idx;
      5'b11100:
        casez_tmp_159 = ldq_28_bits_uop_rxq_idx;
      5'b11101:
        casez_tmp_159 = ldq_29_bits_uop_rxq_idx;
      5'b11110:
        casez_tmp_159 = ldq_30_bits_uop_rxq_idx;
      default:
        casez_tmp_159 = ldq_31_bits_uop_rxq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_160;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_160 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_160 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_160 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_160 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_160 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_160 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_160 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_160 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_160 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_160 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_160 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_160 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_160 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_160 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_160 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_160 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_160 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_160 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_160 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_160 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_160 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_160 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_160 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_160 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_160 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_160 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_160 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_160 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_160 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_160 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_160 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_160 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_161;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_161 = ldq_0_bits_uop_prs1;
      5'b00001:
        casez_tmp_161 = ldq_1_bits_uop_prs1;
      5'b00010:
        casez_tmp_161 = ldq_2_bits_uop_prs1;
      5'b00011:
        casez_tmp_161 = ldq_3_bits_uop_prs1;
      5'b00100:
        casez_tmp_161 = ldq_4_bits_uop_prs1;
      5'b00101:
        casez_tmp_161 = ldq_5_bits_uop_prs1;
      5'b00110:
        casez_tmp_161 = ldq_6_bits_uop_prs1;
      5'b00111:
        casez_tmp_161 = ldq_7_bits_uop_prs1;
      5'b01000:
        casez_tmp_161 = ldq_8_bits_uop_prs1;
      5'b01001:
        casez_tmp_161 = ldq_9_bits_uop_prs1;
      5'b01010:
        casez_tmp_161 = ldq_10_bits_uop_prs1;
      5'b01011:
        casez_tmp_161 = ldq_11_bits_uop_prs1;
      5'b01100:
        casez_tmp_161 = ldq_12_bits_uop_prs1;
      5'b01101:
        casez_tmp_161 = ldq_13_bits_uop_prs1;
      5'b01110:
        casez_tmp_161 = ldq_14_bits_uop_prs1;
      5'b01111:
        casez_tmp_161 = ldq_15_bits_uop_prs1;
      5'b10000:
        casez_tmp_161 = ldq_16_bits_uop_prs1;
      5'b10001:
        casez_tmp_161 = ldq_17_bits_uop_prs1;
      5'b10010:
        casez_tmp_161 = ldq_18_bits_uop_prs1;
      5'b10011:
        casez_tmp_161 = ldq_19_bits_uop_prs1;
      5'b10100:
        casez_tmp_161 = ldq_20_bits_uop_prs1;
      5'b10101:
        casez_tmp_161 = ldq_21_bits_uop_prs1;
      5'b10110:
        casez_tmp_161 = ldq_22_bits_uop_prs1;
      5'b10111:
        casez_tmp_161 = ldq_23_bits_uop_prs1;
      5'b11000:
        casez_tmp_161 = ldq_24_bits_uop_prs1;
      5'b11001:
        casez_tmp_161 = ldq_25_bits_uop_prs1;
      5'b11010:
        casez_tmp_161 = ldq_26_bits_uop_prs1;
      5'b11011:
        casez_tmp_161 = ldq_27_bits_uop_prs1;
      5'b11100:
        casez_tmp_161 = ldq_28_bits_uop_prs1;
      5'b11101:
        casez_tmp_161 = ldq_29_bits_uop_prs1;
      5'b11110:
        casez_tmp_161 = ldq_30_bits_uop_prs1;
      default:
        casez_tmp_161 = ldq_31_bits_uop_prs1;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_162;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_162 = ldq_0_bits_uop_prs2;
      5'b00001:
        casez_tmp_162 = ldq_1_bits_uop_prs2;
      5'b00010:
        casez_tmp_162 = ldq_2_bits_uop_prs2;
      5'b00011:
        casez_tmp_162 = ldq_3_bits_uop_prs2;
      5'b00100:
        casez_tmp_162 = ldq_4_bits_uop_prs2;
      5'b00101:
        casez_tmp_162 = ldq_5_bits_uop_prs2;
      5'b00110:
        casez_tmp_162 = ldq_6_bits_uop_prs2;
      5'b00111:
        casez_tmp_162 = ldq_7_bits_uop_prs2;
      5'b01000:
        casez_tmp_162 = ldq_8_bits_uop_prs2;
      5'b01001:
        casez_tmp_162 = ldq_9_bits_uop_prs2;
      5'b01010:
        casez_tmp_162 = ldq_10_bits_uop_prs2;
      5'b01011:
        casez_tmp_162 = ldq_11_bits_uop_prs2;
      5'b01100:
        casez_tmp_162 = ldq_12_bits_uop_prs2;
      5'b01101:
        casez_tmp_162 = ldq_13_bits_uop_prs2;
      5'b01110:
        casez_tmp_162 = ldq_14_bits_uop_prs2;
      5'b01111:
        casez_tmp_162 = ldq_15_bits_uop_prs2;
      5'b10000:
        casez_tmp_162 = ldq_16_bits_uop_prs2;
      5'b10001:
        casez_tmp_162 = ldq_17_bits_uop_prs2;
      5'b10010:
        casez_tmp_162 = ldq_18_bits_uop_prs2;
      5'b10011:
        casez_tmp_162 = ldq_19_bits_uop_prs2;
      5'b10100:
        casez_tmp_162 = ldq_20_bits_uop_prs2;
      5'b10101:
        casez_tmp_162 = ldq_21_bits_uop_prs2;
      5'b10110:
        casez_tmp_162 = ldq_22_bits_uop_prs2;
      5'b10111:
        casez_tmp_162 = ldq_23_bits_uop_prs2;
      5'b11000:
        casez_tmp_162 = ldq_24_bits_uop_prs2;
      5'b11001:
        casez_tmp_162 = ldq_25_bits_uop_prs2;
      5'b11010:
        casez_tmp_162 = ldq_26_bits_uop_prs2;
      5'b11011:
        casez_tmp_162 = ldq_27_bits_uop_prs2;
      5'b11100:
        casez_tmp_162 = ldq_28_bits_uop_prs2;
      5'b11101:
        casez_tmp_162 = ldq_29_bits_uop_prs2;
      5'b11110:
        casez_tmp_162 = ldq_30_bits_uop_prs2;
      default:
        casez_tmp_162 = ldq_31_bits_uop_prs2;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_163;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_163 = ldq_0_bits_uop_prs3;
      5'b00001:
        casez_tmp_163 = ldq_1_bits_uop_prs3;
      5'b00010:
        casez_tmp_163 = ldq_2_bits_uop_prs3;
      5'b00011:
        casez_tmp_163 = ldq_3_bits_uop_prs3;
      5'b00100:
        casez_tmp_163 = ldq_4_bits_uop_prs3;
      5'b00101:
        casez_tmp_163 = ldq_5_bits_uop_prs3;
      5'b00110:
        casez_tmp_163 = ldq_6_bits_uop_prs3;
      5'b00111:
        casez_tmp_163 = ldq_7_bits_uop_prs3;
      5'b01000:
        casez_tmp_163 = ldq_8_bits_uop_prs3;
      5'b01001:
        casez_tmp_163 = ldq_9_bits_uop_prs3;
      5'b01010:
        casez_tmp_163 = ldq_10_bits_uop_prs3;
      5'b01011:
        casez_tmp_163 = ldq_11_bits_uop_prs3;
      5'b01100:
        casez_tmp_163 = ldq_12_bits_uop_prs3;
      5'b01101:
        casez_tmp_163 = ldq_13_bits_uop_prs3;
      5'b01110:
        casez_tmp_163 = ldq_14_bits_uop_prs3;
      5'b01111:
        casez_tmp_163 = ldq_15_bits_uop_prs3;
      5'b10000:
        casez_tmp_163 = ldq_16_bits_uop_prs3;
      5'b10001:
        casez_tmp_163 = ldq_17_bits_uop_prs3;
      5'b10010:
        casez_tmp_163 = ldq_18_bits_uop_prs3;
      5'b10011:
        casez_tmp_163 = ldq_19_bits_uop_prs3;
      5'b10100:
        casez_tmp_163 = ldq_20_bits_uop_prs3;
      5'b10101:
        casez_tmp_163 = ldq_21_bits_uop_prs3;
      5'b10110:
        casez_tmp_163 = ldq_22_bits_uop_prs3;
      5'b10111:
        casez_tmp_163 = ldq_23_bits_uop_prs3;
      5'b11000:
        casez_tmp_163 = ldq_24_bits_uop_prs3;
      5'b11001:
        casez_tmp_163 = ldq_25_bits_uop_prs3;
      5'b11010:
        casez_tmp_163 = ldq_26_bits_uop_prs3;
      5'b11011:
        casez_tmp_163 = ldq_27_bits_uop_prs3;
      5'b11100:
        casez_tmp_163 = ldq_28_bits_uop_prs3;
      5'b11101:
        casez_tmp_163 = ldq_29_bits_uop_prs3;
      5'b11110:
        casez_tmp_163 = ldq_30_bits_uop_prs3;
      default:
        casez_tmp_163 = ldq_31_bits_uop_prs3;
    endcase
  end // always @(*)
  reg         casez_tmp_164;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_164 = ldq_0_bits_uop_prs1_busy;
      5'b00001:
        casez_tmp_164 = ldq_1_bits_uop_prs1_busy;
      5'b00010:
        casez_tmp_164 = ldq_2_bits_uop_prs1_busy;
      5'b00011:
        casez_tmp_164 = ldq_3_bits_uop_prs1_busy;
      5'b00100:
        casez_tmp_164 = ldq_4_bits_uop_prs1_busy;
      5'b00101:
        casez_tmp_164 = ldq_5_bits_uop_prs1_busy;
      5'b00110:
        casez_tmp_164 = ldq_6_bits_uop_prs1_busy;
      5'b00111:
        casez_tmp_164 = ldq_7_bits_uop_prs1_busy;
      5'b01000:
        casez_tmp_164 = ldq_8_bits_uop_prs1_busy;
      5'b01001:
        casez_tmp_164 = ldq_9_bits_uop_prs1_busy;
      5'b01010:
        casez_tmp_164 = ldq_10_bits_uop_prs1_busy;
      5'b01011:
        casez_tmp_164 = ldq_11_bits_uop_prs1_busy;
      5'b01100:
        casez_tmp_164 = ldq_12_bits_uop_prs1_busy;
      5'b01101:
        casez_tmp_164 = ldq_13_bits_uop_prs1_busy;
      5'b01110:
        casez_tmp_164 = ldq_14_bits_uop_prs1_busy;
      5'b01111:
        casez_tmp_164 = ldq_15_bits_uop_prs1_busy;
      5'b10000:
        casez_tmp_164 = ldq_16_bits_uop_prs1_busy;
      5'b10001:
        casez_tmp_164 = ldq_17_bits_uop_prs1_busy;
      5'b10010:
        casez_tmp_164 = ldq_18_bits_uop_prs1_busy;
      5'b10011:
        casez_tmp_164 = ldq_19_bits_uop_prs1_busy;
      5'b10100:
        casez_tmp_164 = ldq_20_bits_uop_prs1_busy;
      5'b10101:
        casez_tmp_164 = ldq_21_bits_uop_prs1_busy;
      5'b10110:
        casez_tmp_164 = ldq_22_bits_uop_prs1_busy;
      5'b10111:
        casez_tmp_164 = ldq_23_bits_uop_prs1_busy;
      5'b11000:
        casez_tmp_164 = ldq_24_bits_uop_prs1_busy;
      5'b11001:
        casez_tmp_164 = ldq_25_bits_uop_prs1_busy;
      5'b11010:
        casez_tmp_164 = ldq_26_bits_uop_prs1_busy;
      5'b11011:
        casez_tmp_164 = ldq_27_bits_uop_prs1_busy;
      5'b11100:
        casez_tmp_164 = ldq_28_bits_uop_prs1_busy;
      5'b11101:
        casez_tmp_164 = ldq_29_bits_uop_prs1_busy;
      5'b11110:
        casez_tmp_164 = ldq_30_bits_uop_prs1_busy;
      default:
        casez_tmp_164 = ldq_31_bits_uop_prs1_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_165;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_165 = ldq_0_bits_uop_prs2_busy;
      5'b00001:
        casez_tmp_165 = ldq_1_bits_uop_prs2_busy;
      5'b00010:
        casez_tmp_165 = ldq_2_bits_uop_prs2_busy;
      5'b00011:
        casez_tmp_165 = ldq_3_bits_uop_prs2_busy;
      5'b00100:
        casez_tmp_165 = ldq_4_bits_uop_prs2_busy;
      5'b00101:
        casez_tmp_165 = ldq_5_bits_uop_prs2_busy;
      5'b00110:
        casez_tmp_165 = ldq_6_bits_uop_prs2_busy;
      5'b00111:
        casez_tmp_165 = ldq_7_bits_uop_prs2_busy;
      5'b01000:
        casez_tmp_165 = ldq_8_bits_uop_prs2_busy;
      5'b01001:
        casez_tmp_165 = ldq_9_bits_uop_prs2_busy;
      5'b01010:
        casez_tmp_165 = ldq_10_bits_uop_prs2_busy;
      5'b01011:
        casez_tmp_165 = ldq_11_bits_uop_prs2_busy;
      5'b01100:
        casez_tmp_165 = ldq_12_bits_uop_prs2_busy;
      5'b01101:
        casez_tmp_165 = ldq_13_bits_uop_prs2_busy;
      5'b01110:
        casez_tmp_165 = ldq_14_bits_uop_prs2_busy;
      5'b01111:
        casez_tmp_165 = ldq_15_bits_uop_prs2_busy;
      5'b10000:
        casez_tmp_165 = ldq_16_bits_uop_prs2_busy;
      5'b10001:
        casez_tmp_165 = ldq_17_bits_uop_prs2_busy;
      5'b10010:
        casez_tmp_165 = ldq_18_bits_uop_prs2_busy;
      5'b10011:
        casez_tmp_165 = ldq_19_bits_uop_prs2_busy;
      5'b10100:
        casez_tmp_165 = ldq_20_bits_uop_prs2_busy;
      5'b10101:
        casez_tmp_165 = ldq_21_bits_uop_prs2_busy;
      5'b10110:
        casez_tmp_165 = ldq_22_bits_uop_prs2_busy;
      5'b10111:
        casez_tmp_165 = ldq_23_bits_uop_prs2_busy;
      5'b11000:
        casez_tmp_165 = ldq_24_bits_uop_prs2_busy;
      5'b11001:
        casez_tmp_165 = ldq_25_bits_uop_prs2_busy;
      5'b11010:
        casez_tmp_165 = ldq_26_bits_uop_prs2_busy;
      5'b11011:
        casez_tmp_165 = ldq_27_bits_uop_prs2_busy;
      5'b11100:
        casez_tmp_165 = ldq_28_bits_uop_prs2_busy;
      5'b11101:
        casez_tmp_165 = ldq_29_bits_uop_prs2_busy;
      5'b11110:
        casez_tmp_165 = ldq_30_bits_uop_prs2_busy;
      default:
        casez_tmp_165 = ldq_31_bits_uop_prs2_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_166;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_166 = ldq_0_bits_uop_prs3_busy;
      5'b00001:
        casez_tmp_166 = ldq_1_bits_uop_prs3_busy;
      5'b00010:
        casez_tmp_166 = ldq_2_bits_uop_prs3_busy;
      5'b00011:
        casez_tmp_166 = ldq_3_bits_uop_prs3_busy;
      5'b00100:
        casez_tmp_166 = ldq_4_bits_uop_prs3_busy;
      5'b00101:
        casez_tmp_166 = ldq_5_bits_uop_prs3_busy;
      5'b00110:
        casez_tmp_166 = ldq_6_bits_uop_prs3_busy;
      5'b00111:
        casez_tmp_166 = ldq_7_bits_uop_prs3_busy;
      5'b01000:
        casez_tmp_166 = ldq_8_bits_uop_prs3_busy;
      5'b01001:
        casez_tmp_166 = ldq_9_bits_uop_prs3_busy;
      5'b01010:
        casez_tmp_166 = ldq_10_bits_uop_prs3_busy;
      5'b01011:
        casez_tmp_166 = ldq_11_bits_uop_prs3_busy;
      5'b01100:
        casez_tmp_166 = ldq_12_bits_uop_prs3_busy;
      5'b01101:
        casez_tmp_166 = ldq_13_bits_uop_prs3_busy;
      5'b01110:
        casez_tmp_166 = ldq_14_bits_uop_prs3_busy;
      5'b01111:
        casez_tmp_166 = ldq_15_bits_uop_prs3_busy;
      5'b10000:
        casez_tmp_166 = ldq_16_bits_uop_prs3_busy;
      5'b10001:
        casez_tmp_166 = ldq_17_bits_uop_prs3_busy;
      5'b10010:
        casez_tmp_166 = ldq_18_bits_uop_prs3_busy;
      5'b10011:
        casez_tmp_166 = ldq_19_bits_uop_prs3_busy;
      5'b10100:
        casez_tmp_166 = ldq_20_bits_uop_prs3_busy;
      5'b10101:
        casez_tmp_166 = ldq_21_bits_uop_prs3_busy;
      5'b10110:
        casez_tmp_166 = ldq_22_bits_uop_prs3_busy;
      5'b10111:
        casez_tmp_166 = ldq_23_bits_uop_prs3_busy;
      5'b11000:
        casez_tmp_166 = ldq_24_bits_uop_prs3_busy;
      5'b11001:
        casez_tmp_166 = ldq_25_bits_uop_prs3_busy;
      5'b11010:
        casez_tmp_166 = ldq_26_bits_uop_prs3_busy;
      5'b11011:
        casez_tmp_166 = ldq_27_bits_uop_prs3_busy;
      5'b11100:
        casez_tmp_166 = ldq_28_bits_uop_prs3_busy;
      5'b11101:
        casez_tmp_166 = ldq_29_bits_uop_prs3_busy;
      5'b11110:
        casez_tmp_166 = ldq_30_bits_uop_prs3_busy;
      default:
        casez_tmp_166 = ldq_31_bits_uop_prs3_busy;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_167;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_167 = ldq_0_bits_uop_stale_pdst;
      5'b00001:
        casez_tmp_167 = ldq_1_bits_uop_stale_pdst;
      5'b00010:
        casez_tmp_167 = ldq_2_bits_uop_stale_pdst;
      5'b00011:
        casez_tmp_167 = ldq_3_bits_uop_stale_pdst;
      5'b00100:
        casez_tmp_167 = ldq_4_bits_uop_stale_pdst;
      5'b00101:
        casez_tmp_167 = ldq_5_bits_uop_stale_pdst;
      5'b00110:
        casez_tmp_167 = ldq_6_bits_uop_stale_pdst;
      5'b00111:
        casez_tmp_167 = ldq_7_bits_uop_stale_pdst;
      5'b01000:
        casez_tmp_167 = ldq_8_bits_uop_stale_pdst;
      5'b01001:
        casez_tmp_167 = ldq_9_bits_uop_stale_pdst;
      5'b01010:
        casez_tmp_167 = ldq_10_bits_uop_stale_pdst;
      5'b01011:
        casez_tmp_167 = ldq_11_bits_uop_stale_pdst;
      5'b01100:
        casez_tmp_167 = ldq_12_bits_uop_stale_pdst;
      5'b01101:
        casez_tmp_167 = ldq_13_bits_uop_stale_pdst;
      5'b01110:
        casez_tmp_167 = ldq_14_bits_uop_stale_pdst;
      5'b01111:
        casez_tmp_167 = ldq_15_bits_uop_stale_pdst;
      5'b10000:
        casez_tmp_167 = ldq_16_bits_uop_stale_pdst;
      5'b10001:
        casez_tmp_167 = ldq_17_bits_uop_stale_pdst;
      5'b10010:
        casez_tmp_167 = ldq_18_bits_uop_stale_pdst;
      5'b10011:
        casez_tmp_167 = ldq_19_bits_uop_stale_pdst;
      5'b10100:
        casez_tmp_167 = ldq_20_bits_uop_stale_pdst;
      5'b10101:
        casez_tmp_167 = ldq_21_bits_uop_stale_pdst;
      5'b10110:
        casez_tmp_167 = ldq_22_bits_uop_stale_pdst;
      5'b10111:
        casez_tmp_167 = ldq_23_bits_uop_stale_pdst;
      5'b11000:
        casez_tmp_167 = ldq_24_bits_uop_stale_pdst;
      5'b11001:
        casez_tmp_167 = ldq_25_bits_uop_stale_pdst;
      5'b11010:
        casez_tmp_167 = ldq_26_bits_uop_stale_pdst;
      5'b11011:
        casez_tmp_167 = ldq_27_bits_uop_stale_pdst;
      5'b11100:
        casez_tmp_167 = ldq_28_bits_uop_stale_pdst;
      5'b11101:
        casez_tmp_167 = ldq_29_bits_uop_stale_pdst;
      5'b11110:
        casez_tmp_167 = ldq_30_bits_uop_stale_pdst;
      default:
        casez_tmp_167 = ldq_31_bits_uop_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_168;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_168 = ldq_0_bits_uop_exception;
      5'b00001:
        casez_tmp_168 = ldq_1_bits_uop_exception;
      5'b00010:
        casez_tmp_168 = ldq_2_bits_uop_exception;
      5'b00011:
        casez_tmp_168 = ldq_3_bits_uop_exception;
      5'b00100:
        casez_tmp_168 = ldq_4_bits_uop_exception;
      5'b00101:
        casez_tmp_168 = ldq_5_bits_uop_exception;
      5'b00110:
        casez_tmp_168 = ldq_6_bits_uop_exception;
      5'b00111:
        casez_tmp_168 = ldq_7_bits_uop_exception;
      5'b01000:
        casez_tmp_168 = ldq_8_bits_uop_exception;
      5'b01001:
        casez_tmp_168 = ldq_9_bits_uop_exception;
      5'b01010:
        casez_tmp_168 = ldq_10_bits_uop_exception;
      5'b01011:
        casez_tmp_168 = ldq_11_bits_uop_exception;
      5'b01100:
        casez_tmp_168 = ldq_12_bits_uop_exception;
      5'b01101:
        casez_tmp_168 = ldq_13_bits_uop_exception;
      5'b01110:
        casez_tmp_168 = ldq_14_bits_uop_exception;
      5'b01111:
        casez_tmp_168 = ldq_15_bits_uop_exception;
      5'b10000:
        casez_tmp_168 = ldq_16_bits_uop_exception;
      5'b10001:
        casez_tmp_168 = ldq_17_bits_uop_exception;
      5'b10010:
        casez_tmp_168 = ldq_18_bits_uop_exception;
      5'b10011:
        casez_tmp_168 = ldq_19_bits_uop_exception;
      5'b10100:
        casez_tmp_168 = ldq_20_bits_uop_exception;
      5'b10101:
        casez_tmp_168 = ldq_21_bits_uop_exception;
      5'b10110:
        casez_tmp_168 = ldq_22_bits_uop_exception;
      5'b10111:
        casez_tmp_168 = ldq_23_bits_uop_exception;
      5'b11000:
        casez_tmp_168 = ldq_24_bits_uop_exception;
      5'b11001:
        casez_tmp_168 = ldq_25_bits_uop_exception;
      5'b11010:
        casez_tmp_168 = ldq_26_bits_uop_exception;
      5'b11011:
        casez_tmp_168 = ldq_27_bits_uop_exception;
      5'b11100:
        casez_tmp_168 = ldq_28_bits_uop_exception;
      5'b11101:
        casez_tmp_168 = ldq_29_bits_uop_exception;
      5'b11110:
        casez_tmp_168 = ldq_30_bits_uop_exception;
      default:
        casez_tmp_168 = ldq_31_bits_uop_exception;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_169;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_169 = ldq_0_bits_uop_exc_cause;
      5'b00001:
        casez_tmp_169 = ldq_1_bits_uop_exc_cause;
      5'b00010:
        casez_tmp_169 = ldq_2_bits_uop_exc_cause;
      5'b00011:
        casez_tmp_169 = ldq_3_bits_uop_exc_cause;
      5'b00100:
        casez_tmp_169 = ldq_4_bits_uop_exc_cause;
      5'b00101:
        casez_tmp_169 = ldq_5_bits_uop_exc_cause;
      5'b00110:
        casez_tmp_169 = ldq_6_bits_uop_exc_cause;
      5'b00111:
        casez_tmp_169 = ldq_7_bits_uop_exc_cause;
      5'b01000:
        casez_tmp_169 = ldq_8_bits_uop_exc_cause;
      5'b01001:
        casez_tmp_169 = ldq_9_bits_uop_exc_cause;
      5'b01010:
        casez_tmp_169 = ldq_10_bits_uop_exc_cause;
      5'b01011:
        casez_tmp_169 = ldq_11_bits_uop_exc_cause;
      5'b01100:
        casez_tmp_169 = ldq_12_bits_uop_exc_cause;
      5'b01101:
        casez_tmp_169 = ldq_13_bits_uop_exc_cause;
      5'b01110:
        casez_tmp_169 = ldq_14_bits_uop_exc_cause;
      5'b01111:
        casez_tmp_169 = ldq_15_bits_uop_exc_cause;
      5'b10000:
        casez_tmp_169 = ldq_16_bits_uop_exc_cause;
      5'b10001:
        casez_tmp_169 = ldq_17_bits_uop_exc_cause;
      5'b10010:
        casez_tmp_169 = ldq_18_bits_uop_exc_cause;
      5'b10011:
        casez_tmp_169 = ldq_19_bits_uop_exc_cause;
      5'b10100:
        casez_tmp_169 = ldq_20_bits_uop_exc_cause;
      5'b10101:
        casez_tmp_169 = ldq_21_bits_uop_exc_cause;
      5'b10110:
        casez_tmp_169 = ldq_22_bits_uop_exc_cause;
      5'b10111:
        casez_tmp_169 = ldq_23_bits_uop_exc_cause;
      5'b11000:
        casez_tmp_169 = ldq_24_bits_uop_exc_cause;
      5'b11001:
        casez_tmp_169 = ldq_25_bits_uop_exc_cause;
      5'b11010:
        casez_tmp_169 = ldq_26_bits_uop_exc_cause;
      5'b11011:
        casez_tmp_169 = ldq_27_bits_uop_exc_cause;
      5'b11100:
        casez_tmp_169 = ldq_28_bits_uop_exc_cause;
      5'b11101:
        casez_tmp_169 = ldq_29_bits_uop_exc_cause;
      5'b11110:
        casez_tmp_169 = ldq_30_bits_uop_exc_cause;
      default:
        casez_tmp_169 = ldq_31_bits_uop_exc_cause;
    endcase
  end // always @(*)
  reg         casez_tmp_170;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_170 = ldq_0_bits_uop_bypassable;
      5'b00001:
        casez_tmp_170 = ldq_1_bits_uop_bypassable;
      5'b00010:
        casez_tmp_170 = ldq_2_bits_uop_bypassable;
      5'b00011:
        casez_tmp_170 = ldq_3_bits_uop_bypassable;
      5'b00100:
        casez_tmp_170 = ldq_4_bits_uop_bypassable;
      5'b00101:
        casez_tmp_170 = ldq_5_bits_uop_bypassable;
      5'b00110:
        casez_tmp_170 = ldq_6_bits_uop_bypassable;
      5'b00111:
        casez_tmp_170 = ldq_7_bits_uop_bypassable;
      5'b01000:
        casez_tmp_170 = ldq_8_bits_uop_bypassable;
      5'b01001:
        casez_tmp_170 = ldq_9_bits_uop_bypassable;
      5'b01010:
        casez_tmp_170 = ldq_10_bits_uop_bypassable;
      5'b01011:
        casez_tmp_170 = ldq_11_bits_uop_bypassable;
      5'b01100:
        casez_tmp_170 = ldq_12_bits_uop_bypassable;
      5'b01101:
        casez_tmp_170 = ldq_13_bits_uop_bypassable;
      5'b01110:
        casez_tmp_170 = ldq_14_bits_uop_bypassable;
      5'b01111:
        casez_tmp_170 = ldq_15_bits_uop_bypassable;
      5'b10000:
        casez_tmp_170 = ldq_16_bits_uop_bypassable;
      5'b10001:
        casez_tmp_170 = ldq_17_bits_uop_bypassable;
      5'b10010:
        casez_tmp_170 = ldq_18_bits_uop_bypassable;
      5'b10011:
        casez_tmp_170 = ldq_19_bits_uop_bypassable;
      5'b10100:
        casez_tmp_170 = ldq_20_bits_uop_bypassable;
      5'b10101:
        casez_tmp_170 = ldq_21_bits_uop_bypassable;
      5'b10110:
        casez_tmp_170 = ldq_22_bits_uop_bypassable;
      5'b10111:
        casez_tmp_170 = ldq_23_bits_uop_bypassable;
      5'b11000:
        casez_tmp_170 = ldq_24_bits_uop_bypassable;
      5'b11001:
        casez_tmp_170 = ldq_25_bits_uop_bypassable;
      5'b11010:
        casez_tmp_170 = ldq_26_bits_uop_bypassable;
      5'b11011:
        casez_tmp_170 = ldq_27_bits_uop_bypassable;
      5'b11100:
        casez_tmp_170 = ldq_28_bits_uop_bypassable;
      5'b11101:
        casez_tmp_170 = ldq_29_bits_uop_bypassable;
      5'b11110:
        casez_tmp_170 = ldq_30_bits_uop_bypassable;
      default:
        casez_tmp_170 = ldq_31_bits_uop_bypassable;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_171;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_171 = ldq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_171 = ldq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_171 = ldq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_171 = ldq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_171 = ldq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_171 = ldq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_171 = ldq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_171 = ldq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_171 = ldq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_171 = ldq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_171 = ldq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_171 = ldq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_171 = ldq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_171 = ldq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_171 = ldq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_171 = ldq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_171 = ldq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_171 = ldq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_171 = ldq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_171 = ldq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_171 = ldq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_171 = ldq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_171 = ldq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_171 = ldq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_171 = ldq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_171 = ldq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_171 = ldq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_171 = ldq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_171 = ldq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_171 = ldq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_171 = ldq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_171 = ldq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_172;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_172 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_172 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_172 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_172 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_172 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_172 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_172 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_172 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_172 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_172 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_172 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_172 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_172 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_172 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_172 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_172 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_172 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_172 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_172 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_172 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_172 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_172 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_172 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_172 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_172 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_172 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_172 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_172 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_172 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_172 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_172 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_172 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_173;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_173 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_173 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_173 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_173 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_173 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_173 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_173 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_173 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_173 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_173 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_173 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_173 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_173 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_173 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_173 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_173 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_173 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_173 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_173 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_173 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_173 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_173 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_173 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_173 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_173 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_173 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_173 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_173 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_173 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_173 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_173 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_173 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  reg         casez_tmp_174;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_174 = ldq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_174 = ldq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_174 = ldq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_174 = ldq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_174 = ldq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_174 = ldq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_174 = ldq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_174 = ldq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_174 = ldq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_174 = ldq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_174 = ldq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_174 = ldq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_174 = ldq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_174 = ldq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_174 = ldq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_174 = ldq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_174 = ldq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_174 = ldq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_174 = ldq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_174 = ldq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_174 = ldq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_174 = ldq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_174 = ldq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_174 = ldq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_174 = ldq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_174 = ldq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_174 = ldq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_174 = ldq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_174 = ldq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_174 = ldq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_174 = ldq_30_bits_uop_is_fence;
      default:
        casez_tmp_174 = ldq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  reg         casez_tmp_175;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_175 = ldq_0_bits_uop_is_fencei;
      5'b00001:
        casez_tmp_175 = ldq_1_bits_uop_is_fencei;
      5'b00010:
        casez_tmp_175 = ldq_2_bits_uop_is_fencei;
      5'b00011:
        casez_tmp_175 = ldq_3_bits_uop_is_fencei;
      5'b00100:
        casez_tmp_175 = ldq_4_bits_uop_is_fencei;
      5'b00101:
        casez_tmp_175 = ldq_5_bits_uop_is_fencei;
      5'b00110:
        casez_tmp_175 = ldq_6_bits_uop_is_fencei;
      5'b00111:
        casez_tmp_175 = ldq_7_bits_uop_is_fencei;
      5'b01000:
        casez_tmp_175 = ldq_8_bits_uop_is_fencei;
      5'b01001:
        casez_tmp_175 = ldq_9_bits_uop_is_fencei;
      5'b01010:
        casez_tmp_175 = ldq_10_bits_uop_is_fencei;
      5'b01011:
        casez_tmp_175 = ldq_11_bits_uop_is_fencei;
      5'b01100:
        casez_tmp_175 = ldq_12_bits_uop_is_fencei;
      5'b01101:
        casez_tmp_175 = ldq_13_bits_uop_is_fencei;
      5'b01110:
        casez_tmp_175 = ldq_14_bits_uop_is_fencei;
      5'b01111:
        casez_tmp_175 = ldq_15_bits_uop_is_fencei;
      5'b10000:
        casez_tmp_175 = ldq_16_bits_uop_is_fencei;
      5'b10001:
        casez_tmp_175 = ldq_17_bits_uop_is_fencei;
      5'b10010:
        casez_tmp_175 = ldq_18_bits_uop_is_fencei;
      5'b10011:
        casez_tmp_175 = ldq_19_bits_uop_is_fencei;
      5'b10100:
        casez_tmp_175 = ldq_20_bits_uop_is_fencei;
      5'b10101:
        casez_tmp_175 = ldq_21_bits_uop_is_fencei;
      5'b10110:
        casez_tmp_175 = ldq_22_bits_uop_is_fencei;
      5'b10111:
        casez_tmp_175 = ldq_23_bits_uop_is_fencei;
      5'b11000:
        casez_tmp_175 = ldq_24_bits_uop_is_fencei;
      5'b11001:
        casez_tmp_175 = ldq_25_bits_uop_is_fencei;
      5'b11010:
        casez_tmp_175 = ldq_26_bits_uop_is_fencei;
      5'b11011:
        casez_tmp_175 = ldq_27_bits_uop_is_fencei;
      5'b11100:
        casez_tmp_175 = ldq_28_bits_uop_is_fencei;
      5'b11101:
        casez_tmp_175 = ldq_29_bits_uop_is_fencei;
      5'b11110:
        casez_tmp_175 = ldq_30_bits_uop_is_fencei;
      default:
        casez_tmp_175 = ldq_31_bits_uop_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_176;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_176 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_176 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_176 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_176 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_176 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_176 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_176 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_176 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_176 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_176 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_176 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_176 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_176 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_176 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_176 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_176 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_176 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_176 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_176 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_176 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_176 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_176 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_176 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_176 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_176 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_176 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_176 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_176 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_176 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_176 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_176 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_176 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_177;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_177 = ldq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_177 = ldq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_177 = ldq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_177 = ldq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_177 = ldq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_177 = ldq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_177 = ldq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_177 = ldq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_177 = ldq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_177 = ldq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_177 = ldq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_177 = ldq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_177 = ldq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_177 = ldq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_177 = ldq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_177 = ldq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_177 = ldq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_177 = ldq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_177 = ldq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_177 = ldq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_177 = ldq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_177 = ldq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_177 = ldq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_177 = ldq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_177 = ldq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_177 = ldq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_177 = ldq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_177 = ldq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_177 = ldq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_177 = ldq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_177 = ldq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_177 = ldq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_178;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_178 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_178 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_178 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_178 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_178 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_178 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_178 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_178 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_178 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_178 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_178 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_178 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_178 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_178 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_178 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_178 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_178 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_178 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_178 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_178 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_178 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_178 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_178 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_178 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_178 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_178 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_178 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_178 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_178 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_178 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_178 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_178 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_179;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_179 = ldq_0_bits_uop_is_sys_pc2epc;
      5'b00001:
        casez_tmp_179 = ldq_1_bits_uop_is_sys_pc2epc;
      5'b00010:
        casez_tmp_179 = ldq_2_bits_uop_is_sys_pc2epc;
      5'b00011:
        casez_tmp_179 = ldq_3_bits_uop_is_sys_pc2epc;
      5'b00100:
        casez_tmp_179 = ldq_4_bits_uop_is_sys_pc2epc;
      5'b00101:
        casez_tmp_179 = ldq_5_bits_uop_is_sys_pc2epc;
      5'b00110:
        casez_tmp_179 = ldq_6_bits_uop_is_sys_pc2epc;
      5'b00111:
        casez_tmp_179 = ldq_7_bits_uop_is_sys_pc2epc;
      5'b01000:
        casez_tmp_179 = ldq_8_bits_uop_is_sys_pc2epc;
      5'b01001:
        casez_tmp_179 = ldq_9_bits_uop_is_sys_pc2epc;
      5'b01010:
        casez_tmp_179 = ldq_10_bits_uop_is_sys_pc2epc;
      5'b01011:
        casez_tmp_179 = ldq_11_bits_uop_is_sys_pc2epc;
      5'b01100:
        casez_tmp_179 = ldq_12_bits_uop_is_sys_pc2epc;
      5'b01101:
        casez_tmp_179 = ldq_13_bits_uop_is_sys_pc2epc;
      5'b01110:
        casez_tmp_179 = ldq_14_bits_uop_is_sys_pc2epc;
      5'b01111:
        casez_tmp_179 = ldq_15_bits_uop_is_sys_pc2epc;
      5'b10000:
        casez_tmp_179 = ldq_16_bits_uop_is_sys_pc2epc;
      5'b10001:
        casez_tmp_179 = ldq_17_bits_uop_is_sys_pc2epc;
      5'b10010:
        casez_tmp_179 = ldq_18_bits_uop_is_sys_pc2epc;
      5'b10011:
        casez_tmp_179 = ldq_19_bits_uop_is_sys_pc2epc;
      5'b10100:
        casez_tmp_179 = ldq_20_bits_uop_is_sys_pc2epc;
      5'b10101:
        casez_tmp_179 = ldq_21_bits_uop_is_sys_pc2epc;
      5'b10110:
        casez_tmp_179 = ldq_22_bits_uop_is_sys_pc2epc;
      5'b10111:
        casez_tmp_179 = ldq_23_bits_uop_is_sys_pc2epc;
      5'b11000:
        casez_tmp_179 = ldq_24_bits_uop_is_sys_pc2epc;
      5'b11001:
        casez_tmp_179 = ldq_25_bits_uop_is_sys_pc2epc;
      5'b11010:
        casez_tmp_179 = ldq_26_bits_uop_is_sys_pc2epc;
      5'b11011:
        casez_tmp_179 = ldq_27_bits_uop_is_sys_pc2epc;
      5'b11100:
        casez_tmp_179 = ldq_28_bits_uop_is_sys_pc2epc;
      5'b11101:
        casez_tmp_179 = ldq_29_bits_uop_is_sys_pc2epc;
      5'b11110:
        casez_tmp_179 = ldq_30_bits_uop_is_sys_pc2epc;
      default:
        casez_tmp_179 = ldq_31_bits_uop_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_180;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_180 = ldq_0_bits_uop_is_unique;
      5'b00001:
        casez_tmp_180 = ldq_1_bits_uop_is_unique;
      5'b00010:
        casez_tmp_180 = ldq_2_bits_uop_is_unique;
      5'b00011:
        casez_tmp_180 = ldq_3_bits_uop_is_unique;
      5'b00100:
        casez_tmp_180 = ldq_4_bits_uop_is_unique;
      5'b00101:
        casez_tmp_180 = ldq_5_bits_uop_is_unique;
      5'b00110:
        casez_tmp_180 = ldq_6_bits_uop_is_unique;
      5'b00111:
        casez_tmp_180 = ldq_7_bits_uop_is_unique;
      5'b01000:
        casez_tmp_180 = ldq_8_bits_uop_is_unique;
      5'b01001:
        casez_tmp_180 = ldq_9_bits_uop_is_unique;
      5'b01010:
        casez_tmp_180 = ldq_10_bits_uop_is_unique;
      5'b01011:
        casez_tmp_180 = ldq_11_bits_uop_is_unique;
      5'b01100:
        casez_tmp_180 = ldq_12_bits_uop_is_unique;
      5'b01101:
        casez_tmp_180 = ldq_13_bits_uop_is_unique;
      5'b01110:
        casez_tmp_180 = ldq_14_bits_uop_is_unique;
      5'b01111:
        casez_tmp_180 = ldq_15_bits_uop_is_unique;
      5'b10000:
        casez_tmp_180 = ldq_16_bits_uop_is_unique;
      5'b10001:
        casez_tmp_180 = ldq_17_bits_uop_is_unique;
      5'b10010:
        casez_tmp_180 = ldq_18_bits_uop_is_unique;
      5'b10011:
        casez_tmp_180 = ldq_19_bits_uop_is_unique;
      5'b10100:
        casez_tmp_180 = ldq_20_bits_uop_is_unique;
      5'b10101:
        casez_tmp_180 = ldq_21_bits_uop_is_unique;
      5'b10110:
        casez_tmp_180 = ldq_22_bits_uop_is_unique;
      5'b10111:
        casez_tmp_180 = ldq_23_bits_uop_is_unique;
      5'b11000:
        casez_tmp_180 = ldq_24_bits_uop_is_unique;
      5'b11001:
        casez_tmp_180 = ldq_25_bits_uop_is_unique;
      5'b11010:
        casez_tmp_180 = ldq_26_bits_uop_is_unique;
      5'b11011:
        casez_tmp_180 = ldq_27_bits_uop_is_unique;
      5'b11100:
        casez_tmp_180 = ldq_28_bits_uop_is_unique;
      5'b11101:
        casez_tmp_180 = ldq_29_bits_uop_is_unique;
      5'b11110:
        casez_tmp_180 = ldq_30_bits_uop_is_unique;
      default:
        casez_tmp_180 = ldq_31_bits_uop_is_unique;
    endcase
  end // always @(*)
  reg         casez_tmp_181;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_181 = ldq_0_bits_uop_flush_on_commit;
      5'b00001:
        casez_tmp_181 = ldq_1_bits_uop_flush_on_commit;
      5'b00010:
        casez_tmp_181 = ldq_2_bits_uop_flush_on_commit;
      5'b00011:
        casez_tmp_181 = ldq_3_bits_uop_flush_on_commit;
      5'b00100:
        casez_tmp_181 = ldq_4_bits_uop_flush_on_commit;
      5'b00101:
        casez_tmp_181 = ldq_5_bits_uop_flush_on_commit;
      5'b00110:
        casez_tmp_181 = ldq_6_bits_uop_flush_on_commit;
      5'b00111:
        casez_tmp_181 = ldq_7_bits_uop_flush_on_commit;
      5'b01000:
        casez_tmp_181 = ldq_8_bits_uop_flush_on_commit;
      5'b01001:
        casez_tmp_181 = ldq_9_bits_uop_flush_on_commit;
      5'b01010:
        casez_tmp_181 = ldq_10_bits_uop_flush_on_commit;
      5'b01011:
        casez_tmp_181 = ldq_11_bits_uop_flush_on_commit;
      5'b01100:
        casez_tmp_181 = ldq_12_bits_uop_flush_on_commit;
      5'b01101:
        casez_tmp_181 = ldq_13_bits_uop_flush_on_commit;
      5'b01110:
        casez_tmp_181 = ldq_14_bits_uop_flush_on_commit;
      5'b01111:
        casez_tmp_181 = ldq_15_bits_uop_flush_on_commit;
      5'b10000:
        casez_tmp_181 = ldq_16_bits_uop_flush_on_commit;
      5'b10001:
        casez_tmp_181 = ldq_17_bits_uop_flush_on_commit;
      5'b10010:
        casez_tmp_181 = ldq_18_bits_uop_flush_on_commit;
      5'b10011:
        casez_tmp_181 = ldq_19_bits_uop_flush_on_commit;
      5'b10100:
        casez_tmp_181 = ldq_20_bits_uop_flush_on_commit;
      5'b10101:
        casez_tmp_181 = ldq_21_bits_uop_flush_on_commit;
      5'b10110:
        casez_tmp_181 = ldq_22_bits_uop_flush_on_commit;
      5'b10111:
        casez_tmp_181 = ldq_23_bits_uop_flush_on_commit;
      5'b11000:
        casez_tmp_181 = ldq_24_bits_uop_flush_on_commit;
      5'b11001:
        casez_tmp_181 = ldq_25_bits_uop_flush_on_commit;
      5'b11010:
        casez_tmp_181 = ldq_26_bits_uop_flush_on_commit;
      5'b11011:
        casez_tmp_181 = ldq_27_bits_uop_flush_on_commit;
      5'b11100:
        casez_tmp_181 = ldq_28_bits_uop_flush_on_commit;
      5'b11101:
        casez_tmp_181 = ldq_29_bits_uop_flush_on_commit;
      5'b11110:
        casez_tmp_181 = ldq_30_bits_uop_flush_on_commit;
      default:
        casez_tmp_181 = ldq_31_bits_uop_flush_on_commit;
    endcase
  end // always @(*)
  reg         casez_tmp_182;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_182 = ldq_0_bits_uop_ldst_is_rs1;
      5'b00001:
        casez_tmp_182 = ldq_1_bits_uop_ldst_is_rs1;
      5'b00010:
        casez_tmp_182 = ldq_2_bits_uop_ldst_is_rs1;
      5'b00011:
        casez_tmp_182 = ldq_3_bits_uop_ldst_is_rs1;
      5'b00100:
        casez_tmp_182 = ldq_4_bits_uop_ldst_is_rs1;
      5'b00101:
        casez_tmp_182 = ldq_5_bits_uop_ldst_is_rs1;
      5'b00110:
        casez_tmp_182 = ldq_6_bits_uop_ldst_is_rs1;
      5'b00111:
        casez_tmp_182 = ldq_7_bits_uop_ldst_is_rs1;
      5'b01000:
        casez_tmp_182 = ldq_8_bits_uop_ldst_is_rs1;
      5'b01001:
        casez_tmp_182 = ldq_9_bits_uop_ldst_is_rs1;
      5'b01010:
        casez_tmp_182 = ldq_10_bits_uop_ldst_is_rs1;
      5'b01011:
        casez_tmp_182 = ldq_11_bits_uop_ldst_is_rs1;
      5'b01100:
        casez_tmp_182 = ldq_12_bits_uop_ldst_is_rs1;
      5'b01101:
        casez_tmp_182 = ldq_13_bits_uop_ldst_is_rs1;
      5'b01110:
        casez_tmp_182 = ldq_14_bits_uop_ldst_is_rs1;
      5'b01111:
        casez_tmp_182 = ldq_15_bits_uop_ldst_is_rs1;
      5'b10000:
        casez_tmp_182 = ldq_16_bits_uop_ldst_is_rs1;
      5'b10001:
        casez_tmp_182 = ldq_17_bits_uop_ldst_is_rs1;
      5'b10010:
        casez_tmp_182 = ldq_18_bits_uop_ldst_is_rs1;
      5'b10011:
        casez_tmp_182 = ldq_19_bits_uop_ldst_is_rs1;
      5'b10100:
        casez_tmp_182 = ldq_20_bits_uop_ldst_is_rs1;
      5'b10101:
        casez_tmp_182 = ldq_21_bits_uop_ldst_is_rs1;
      5'b10110:
        casez_tmp_182 = ldq_22_bits_uop_ldst_is_rs1;
      5'b10111:
        casez_tmp_182 = ldq_23_bits_uop_ldst_is_rs1;
      5'b11000:
        casez_tmp_182 = ldq_24_bits_uop_ldst_is_rs1;
      5'b11001:
        casez_tmp_182 = ldq_25_bits_uop_ldst_is_rs1;
      5'b11010:
        casez_tmp_182 = ldq_26_bits_uop_ldst_is_rs1;
      5'b11011:
        casez_tmp_182 = ldq_27_bits_uop_ldst_is_rs1;
      5'b11100:
        casez_tmp_182 = ldq_28_bits_uop_ldst_is_rs1;
      5'b11101:
        casez_tmp_182 = ldq_29_bits_uop_ldst_is_rs1;
      5'b11110:
        casez_tmp_182 = ldq_30_bits_uop_ldst_is_rs1;
      default:
        casez_tmp_182 = ldq_31_bits_uop_ldst_is_rs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_183;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_183 = ldq_0_bits_uop_ldst;
      5'b00001:
        casez_tmp_183 = ldq_1_bits_uop_ldst;
      5'b00010:
        casez_tmp_183 = ldq_2_bits_uop_ldst;
      5'b00011:
        casez_tmp_183 = ldq_3_bits_uop_ldst;
      5'b00100:
        casez_tmp_183 = ldq_4_bits_uop_ldst;
      5'b00101:
        casez_tmp_183 = ldq_5_bits_uop_ldst;
      5'b00110:
        casez_tmp_183 = ldq_6_bits_uop_ldst;
      5'b00111:
        casez_tmp_183 = ldq_7_bits_uop_ldst;
      5'b01000:
        casez_tmp_183 = ldq_8_bits_uop_ldst;
      5'b01001:
        casez_tmp_183 = ldq_9_bits_uop_ldst;
      5'b01010:
        casez_tmp_183 = ldq_10_bits_uop_ldst;
      5'b01011:
        casez_tmp_183 = ldq_11_bits_uop_ldst;
      5'b01100:
        casez_tmp_183 = ldq_12_bits_uop_ldst;
      5'b01101:
        casez_tmp_183 = ldq_13_bits_uop_ldst;
      5'b01110:
        casez_tmp_183 = ldq_14_bits_uop_ldst;
      5'b01111:
        casez_tmp_183 = ldq_15_bits_uop_ldst;
      5'b10000:
        casez_tmp_183 = ldq_16_bits_uop_ldst;
      5'b10001:
        casez_tmp_183 = ldq_17_bits_uop_ldst;
      5'b10010:
        casez_tmp_183 = ldq_18_bits_uop_ldst;
      5'b10011:
        casez_tmp_183 = ldq_19_bits_uop_ldst;
      5'b10100:
        casez_tmp_183 = ldq_20_bits_uop_ldst;
      5'b10101:
        casez_tmp_183 = ldq_21_bits_uop_ldst;
      5'b10110:
        casez_tmp_183 = ldq_22_bits_uop_ldst;
      5'b10111:
        casez_tmp_183 = ldq_23_bits_uop_ldst;
      5'b11000:
        casez_tmp_183 = ldq_24_bits_uop_ldst;
      5'b11001:
        casez_tmp_183 = ldq_25_bits_uop_ldst;
      5'b11010:
        casez_tmp_183 = ldq_26_bits_uop_ldst;
      5'b11011:
        casez_tmp_183 = ldq_27_bits_uop_ldst;
      5'b11100:
        casez_tmp_183 = ldq_28_bits_uop_ldst;
      5'b11101:
        casez_tmp_183 = ldq_29_bits_uop_ldst;
      5'b11110:
        casez_tmp_183 = ldq_30_bits_uop_ldst;
      default:
        casez_tmp_183 = ldq_31_bits_uop_ldst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_184;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_184 = ldq_0_bits_uop_lrs1;
      5'b00001:
        casez_tmp_184 = ldq_1_bits_uop_lrs1;
      5'b00010:
        casez_tmp_184 = ldq_2_bits_uop_lrs1;
      5'b00011:
        casez_tmp_184 = ldq_3_bits_uop_lrs1;
      5'b00100:
        casez_tmp_184 = ldq_4_bits_uop_lrs1;
      5'b00101:
        casez_tmp_184 = ldq_5_bits_uop_lrs1;
      5'b00110:
        casez_tmp_184 = ldq_6_bits_uop_lrs1;
      5'b00111:
        casez_tmp_184 = ldq_7_bits_uop_lrs1;
      5'b01000:
        casez_tmp_184 = ldq_8_bits_uop_lrs1;
      5'b01001:
        casez_tmp_184 = ldq_9_bits_uop_lrs1;
      5'b01010:
        casez_tmp_184 = ldq_10_bits_uop_lrs1;
      5'b01011:
        casez_tmp_184 = ldq_11_bits_uop_lrs1;
      5'b01100:
        casez_tmp_184 = ldq_12_bits_uop_lrs1;
      5'b01101:
        casez_tmp_184 = ldq_13_bits_uop_lrs1;
      5'b01110:
        casez_tmp_184 = ldq_14_bits_uop_lrs1;
      5'b01111:
        casez_tmp_184 = ldq_15_bits_uop_lrs1;
      5'b10000:
        casez_tmp_184 = ldq_16_bits_uop_lrs1;
      5'b10001:
        casez_tmp_184 = ldq_17_bits_uop_lrs1;
      5'b10010:
        casez_tmp_184 = ldq_18_bits_uop_lrs1;
      5'b10011:
        casez_tmp_184 = ldq_19_bits_uop_lrs1;
      5'b10100:
        casez_tmp_184 = ldq_20_bits_uop_lrs1;
      5'b10101:
        casez_tmp_184 = ldq_21_bits_uop_lrs1;
      5'b10110:
        casez_tmp_184 = ldq_22_bits_uop_lrs1;
      5'b10111:
        casez_tmp_184 = ldq_23_bits_uop_lrs1;
      5'b11000:
        casez_tmp_184 = ldq_24_bits_uop_lrs1;
      5'b11001:
        casez_tmp_184 = ldq_25_bits_uop_lrs1;
      5'b11010:
        casez_tmp_184 = ldq_26_bits_uop_lrs1;
      5'b11011:
        casez_tmp_184 = ldq_27_bits_uop_lrs1;
      5'b11100:
        casez_tmp_184 = ldq_28_bits_uop_lrs1;
      5'b11101:
        casez_tmp_184 = ldq_29_bits_uop_lrs1;
      5'b11110:
        casez_tmp_184 = ldq_30_bits_uop_lrs1;
      default:
        casez_tmp_184 = ldq_31_bits_uop_lrs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_185;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_185 = ldq_0_bits_uop_lrs2;
      5'b00001:
        casez_tmp_185 = ldq_1_bits_uop_lrs2;
      5'b00010:
        casez_tmp_185 = ldq_2_bits_uop_lrs2;
      5'b00011:
        casez_tmp_185 = ldq_3_bits_uop_lrs2;
      5'b00100:
        casez_tmp_185 = ldq_4_bits_uop_lrs2;
      5'b00101:
        casez_tmp_185 = ldq_5_bits_uop_lrs2;
      5'b00110:
        casez_tmp_185 = ldq_6_bits_uop_lrs2;
      5'b00111:
        casez_tmp_185 = ldq_7_bits_uop_lrs2;
      5'b01000:
        casez_tmp_185 = ldq_8_bits_uop_lrs2;
      5'b01001:
        casez_tmp_185 = ldq_9_bits_uop_lrs2;
      5'b01010:
        casez_tmp_185 = ldq_10_bits_uop_lrs2;
      5'b01011:
        casez_tmp_185 = ldq_11_bits_uop_lrs2;
      5'b01100:
        casez_tmp_185 = ldq_12_bits_uop_lrs2;
      5'b01101:
        casez_tmp_185 = ldq_13_bits_uop_lrs2;
      5'b01110:
        casez_tmp_185 = ldq_14_bits_uop_lrs2;
      5'b01111:
        casez_tmp_185 = ldq_15_bits_uop_lrs2;
      5'b10000:
        casez_tmp_185 = ldq_16_bits_uop_lrs2;
      5'b10001:
        casez_tmp_185 = ldq_17_bits_uop_lrs2;
      5'b10010:
        casez_tmp_185 = ldq_18_bits_uop_lrs2;
      5'b10011:
        casez_tmp_185 = ldq_19_bits_uop_lrs2;
      5'b10100:
        casez_tmp_185 = ldq_20_bits_uop_lrs2;
      5'b10101:
        casez_tmp_185 = ldq_21_bits_uop_lrs2;
      5'b10110:
        casez_tmp_185 = ldq_22_bits_uop_lrs2;
      5'b10111:
        casez_tmp_185 = ldq_23_bits_uop_lrs2;
      5'b11000:
        casez_tmp_185 = ldq_24_bits_uop_lrs2;
      5'b11001:
        casez_tmp_185 = ldq_25_bits_uop_lrs2;
      5'b11010:
        casez_tmp_185 = ldq_26_bits_uop_lrs2;
      5'b11011:
        casez_tmp_185 = ldq_27_bits_uop_lrs2;
      5'b11100:
        casez_tmp_185 = ldq_28_bits_uop_lrs2;
      5'b11101:
        casez_tmp_185 = ldq_29_bits_uop_lrs2;
      5'b11110:
        casez_tmp_185 = ldq_30_bits_uop_lrs2;
      default:
        casez_tmp_185 = ldq_31_bits_uop_lrs2;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_186;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_186 = ldq_0_bits_uop_lrs3;
      5'b00001:
        casez_tmp_186 = ldq_1_bits_uop_lrs3;
      5'b00010:
        casez_tmp_186 = ldq_2_bits_uop_lrs3;
      5'b00011:
        casez_tmp_186 = ldq_3_bits_uop_lrs3;
      5'b00100:
        casez_tmp_186 = ldq_4_bits_uop_lrs3;
      5'b00101:
        casez_tmp_186 = ldq_5_bits_uop_lrs3;
      5'b00110:
        casez_tmp_186 = ldq_6_bits_uop_lrs3;
      5'b00111:
        casez_tmp_186 = ldq_7_bits_uop_lrs3;
      5'b01000:
        casez_tmp_186 = ldq_8_bits_uop_lrs3;
      5'b01001:
        casez_tmp_186 = ldq_9_bits_uop_lrs3;
      5'b01010:
        casez_tmp_186 = ldq_10_bits_uop_lrs3;
      5'b01011:
        casez_tmp_186 = ldq_11_bits_uop_lrs3;
      5'b01100:
        casez_tmp_186 = ldq_12_bits_uop_lrs3;
      5'b01101:
        casez_tmp_186 = ldq_13_bits_uop_lrs3;
      5'b01110:
        casez_tmp_186 = ldq_14_bits_uop_lrs3;
      5'b01111:
        casez_tmp_186 = ldq_15_bits_uop_lrs3;
      5'b10000:
        casez_tmp_186 = ldq_16_bits_uop_lrs3;
      5'b10001:
        casez_tmp_186 = ldq_17_bits_uop_lrs3;
      5'b10010:
        casez_tmp_186 = ldq_18_bits_uop_lrs3;
      5'b10011:
        casez_tmp_186 = ldq_19_bits_uop_lrs3;
      5'b10100:
        casez_tmp_186 = ldq_20_bits_uop_lrs3;
      5'b10101:
        casez_tmp_186 = ldq_21_bits_uop_lrs3;
      5'b10110:
        casez_tmp_186 = ldq_22_bits_uop_lrs3;
      5'b10111:
        casez_tmp_186 = ldq_23_bits_uop_lrs3;
      5'b11000:
        casez_tmp_186 = ldq_24_bits_uop_lrs3;
      5'b11001:
        casez_tmp_186 = ldq_25_bits_uop_lrs3;
      5'b11010:
        casez_tmp_186 = ldq_26_bits_uop_lrs3;
      5'b11011:
        casez_tmp_186 = ldq_27_bits_uop_lrs3;
      5'b11100:
        casez_tmp_186 = ldq_28_bits_uop_lrs3;
      5'b11101:
        casez_tmp_186 = ldq_29_bits_uop_lrs3;
      5'b11110:
        casez_tmp_186 = ldq_30_bits_uop_lrs3;
      default:
        casez_tmp_186 = ldq_31_bits_uop_lrs3;
    endcase
  end // always @(*)
  reg         casez_tmp_187;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_187 = ldq_0_bits_uop_ldst_val;
      5'b00001:
        casez_tmp_187 = ldq_1_bits_uop_ldst_val;
      5'b00010:
        casez_tmp_187 = ldq_2_bits_uop_ldst_val;
      5'b00011:
        casez_tmp_187 = ldq_3_bits_uop_ldst_val;
      5'b00100:
        casez_tmp_187 = ldq_4_bits_uop_ldst_val;
      5'b00101:
        casez_tmp_187 = ldq_5_bits_uop_ldst_val;
      5'b00110:
        casez_tmp_187 = ldq_6_bits_uop_ldst_val;
      5'b00111:
        casez_tmp_187 = ldq_7_bits_uop_ldst_val;
      5'b01000:
        casez_tmp_187 = ldq_8_bits_uop_ldst_val;
      5'b01001:
        casez_tmp_187 = ldq_9_bits_uop_ldst_val;
      5'b01010:
        casez_tmp_187 = ldq_10_bits_uop_ldst_val;
      5'b01011:
        casez_tmp_187 = ldq_11_bits_uop_ldst_val;
      5'b01100:
        casez_tmp_187 = ldq_12_bits_uop_ldst_val;
      5'b01101:
        casez_tmp_187 = ldq_13_bits_uop_ldst_val;
      5'b01110:
        casez_tmp_187 = ldq_14_bits_uop_ldst_val;
      5'b01111:
        casez_tmp_187 = ldq_15_bits_uop_ldst_val;
      5'b10000:
        casez_tmp_187 = ldq_16_bits_uop_ldst_val;
      5'b10001:
        casez_tmp_187 = ldq_17_bits_uop_ldst_val;
      5'b10010:
        casez_tmp_187 = ldq_18_bits_uop_ldst_val;
      5'b10011:
        casez_tmp_187 = ldq_19_bits_uop_ldst_val;
      5'b10100:
        casez_tmp_187 = ldq_20_bits_uop_ldst_val;
      5'b10101:
        casez_tmp_187 = ldq_21_bits_uop_ldst_val;
      5'b10110:
        casez_tmp_187 = ldq_22_bits_uop_ldst_val;
      5'b10111:
        casez_tmp_187 = ldq_23_bits_uop_ldst_val;
      5'b11000:
        casez_tmp_187 = ldq_24_bits_uop_ldst_val;
      5'b11001:
        casez_tmp_187 = ldq_25_bits_uop_ldst_val;
      5'b11010:
        casez_tmp_187 = ldq_26_bits_uop_ldst_val;
      5'b11011:
        casez_tmp_187 = ldq_27_bits_uop_ldst_val;
      5'b11100:
        casez_tmp_187 = ldq_28_bits_uop_ldst_val;
      5'b11101:
        casez_tmp_187 = ldq_29_bits_uop_ldst_val;
      5'b11110:
        casez_tmp_187 = ldq_30_bits_uop_ldst_val;
      default:
        casez_tmp_187 = ldq_31_bits_uop_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_188;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_188 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_188 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_188 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_188 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_188 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_188 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_188 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_188 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_188 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_188 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_188 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_188 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_188 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_188 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_188 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_188 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_188 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_188 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_188 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_188 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_188 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_188 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_188 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_188 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_188 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_188 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_188 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_188 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_188 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_188 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_188 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_188 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_189;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_189 = ldq_0_bits_uop_lrs1_rtype;
      5'b00001:
        casez_tmp_189 = ldq_1_bits_uop_lrs1_rtype;
      5'b00010:
        casez_tmp_189 = ldq_2_bits_uop_lrs1_rtype;
      5'b00011:
        casez_tmp_189 = ldq_3_bits_uop_lrs1_rtype;
      5'b00100:
        casez_tmp_189 = ldq_4_bits_uop_lrs1_rtype;
      5'b00101:
        casez_tmp_189 = ldq_5_bits_uop_lrs1_rtype;
      5'b00110:
        casez_tmp_189 = ldq_6_bits_uop_lrs1_rtype;
      5'b00111:
        casez_tmp_189 = ldq_7_bits_uop_lrs1_rtype;
      5'b01000:
        casez_tmp_189 = ldq_8_bits_uop_lrs1_rtype;
      5'b01001:
        casez_tmp_189 = ldq_9_bits_uop_lrs1_rtype;
      5'b01010:
        casez_tmp_189 = ldq_10_bits_uop_lrs1_rtype;
      5'b01011:
        casez_tmp_189 = ldq_11_bits_uop_lrs1_rtype;
      5'b01100:
        casez_tmp_189 = ldq_12_bits_uop_lrs1_rtype;
      5'b01101:
        casez_tmp_189 = ldq_13_bits_uop_lrs1_rtype;
      5'b01110:
        casez_tmp_189 = ldq_14_bits_uop_lrs1_rtype;
      5'b01111:
        casez_tmp_189 = ldq_15_bits_uop_lrs1_rtype;
      5'b10000:
        casez_tmp_189 = ldq_16_bits_uop_lrs1_rtype;
      5'b10001:
        casez_tmp_189 = ldq_17_bits_uop_lrs1_rtype;
      5'b10010:
        casez_tmp_189 = ldq_18_bits_uop_lrs1_rtype;
      5'b10011:
        casez_tmp_189 = ldq_19_bits_uop_lrs1_rtype;
      5'b10100:
        casez_tmp_189 = ldq_20_bits_uop_lrs1_rtype;
      5'b10101:
        casez_tmp_189 = ldq_21_bits_uop_lrs1_rtype;
      5'b10110:
        casez_tmp_189 = ldq_22_bits_uop_lrs1_rtype;
      5'b10111:
        casez_tmp_189 = ldq_23_bits_uop_lrs1_rtype;
      5'b11000:
        casez_tmp_189 = ldq_24_bits_uop_lrs1_rtype;
      5'b11001:
        casez_tmp_189 = ldq_25_bits_uop_lrs1_rtype;
      5'b11010:
        casez_tmp_189 = ldq_26_bits_uop_lrs1_rtype;
      5'b11011:
        casez_tmp_189 = ldq_27_bits_uop_lrs1_rtype;
      5'b11100:
        casez_tmp_189 = ldq_28_bits_uop_lrs1_rtype;
      5'b11101:
        casez_tmp_189 = ldq_29_bits_uop_lrs1_rtype;
      5'b11110:
        casez_tmp_189 = ldq_30_bits_uop_lrs1_rtype;
      default:
        casez_tmp_189 = ldq_31_bits_uop_lrs1_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_190;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_190 = ldq_0_bits_uop_lrs2_rtype;
      5'b00001:
        casez_tmp_190 = ldq_1_bits_uop_lrs2_rtype;
      5'b00010:
        casez_tmp_190 = ldq_2_bits_uop_lrs2_rtype;
      5'b00011:
        casez_tmp_190 = ldq_3_bits_uop_lrs2_rtype;
      5'b00100:
        casez_tmp_190 = ldq_4_bits_uop_lrs2_rtype;
      5'b00101:
        casez_tmp_190 = ldq_5_bits_uop_lrs2_rtype;
      5'b00110:
        casez_tmp_190 = ldq_6_bits_uop_lrs2_rtype;
      5'b00111:
        casez_tmp_190 = ldq_7_bits_uop_lrs2_rtype;
      5'b01000:
        casez_tmp_190 = ldq_8_bits_uop_lrs2_rtype;
      5'b01001:
        casez_tmp_190 = ldq_9_bits_uop_lrs2_rtype;
      5'b01010:
        casez_tmp_190 = ldq_10_bits_uop_lrs2_rtype;
      5'b01011:
        casez_tmp_190 = ldq_11_bits_uop_lrs2_rtype;
      5'b01100:
        casez_tmp_190 = ldq_12_bits_uop_lrs2_rtype;
      5'b01101:
        casez_tmp_190 = ldq_13_bits_uop_lrs2_rtype;
      5'b01110:
        casez_tmp_190 = ldq_14_bits_uop_lrs2_rtype;
      5'b01111:
        casez_tmp_190 = ldq_15_bits_uop_lrs2_rtype;
      5'b10000:
        casez_tmp_190 = ldq_16_bits_uop_lrs2_rtype;
      5'b10001:
        casez_tmp_190 = ldq_17_bits_uop_lrs2_rtype;
      5'b10010:
        casez_tmp_190 = ldq_18_bits_uop_lrs2_rtype;
      5'b10011:
        casez_tmp_190 = ldq_19_bits_uop_lrs2_rtype;
      5'b10100:
        casez_tmp_190 = ldq_20_bits_uop_lrs2_rtype;
      5'b10101:
        casez_tmp_190 = ldq_21_bits_uop_lrs2_rtype;
      5'b10110:
        casez_tmp_190 = ldq_22_bits_uop_lrs2_rtype;
      5'b10111:
        casez_tmp_190 = ldq_23_bits_uop_lrs2_rtype;
      5'b11000:
        casez_tmp_190 = ldq_24_bits_uop_lrs2_rtype;
      5'b11001:
        casez_tmp_190 = ldq_25_bits_uop_lrs2_rtype;
      5'b11010:
        casez_tmp_190 = ldq_26_bits_uop_lrs2_rtype;
      5'b11011:
        casez_tmp_190 = ldq_27_bits_uop_lrs2_rtype;
      5'b11100:
        casez_tmp_190 = ldq_28_bits_uop_lrs2_rtype;
      5'b11101:
        casez_tmp_190 = ldq_29_bits_uop_lrs2_rtype;
      5'b11110:
        casez_tmp_190 = ldq_30_bits_uop_lrs2_rtype;
      default:
        casez_tmp_190 = ldq_31_bits_uop_lrs2_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_191;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_191 = ldq_0_bits_uop_frs3_en;
      5'b00001:
        casez_tmp_191 = ldq_1_bits_uop_frs3_en;
      5'b00010:
        casez_tmp_191 = ldq_2_bits_uop_frs3_en;
      5'b00011:
        casez_tmp_191 = ldq_3_bits_uop_frs3_en;
      5'b00100:
        casez_tmp_191 = ldq_4_bits_uop_frs3_en;
      5'b00101:
        casez_tmp_191 = ldq_5_bits_uop_frs3_en;
      5'b00110:
        casez_tmp_191 = ldq_6_bits_uop_frs3_en;
      5'b00111:
        casez_tmp_191 = ldq_7_bits_uop_frs3_en;
      5'b01000:
        casez_tmp_191 = ldq_8_bits_uop_frs3_en;
      5'b01001:
        casez_tmp_191 = ldq_9_bits_uop_frs3_en;
      5'b01010:
        casez_tmp_191 = ldq_10_bits_uop_frs3_en;
      5'b01011:
        casez_tmp_191 = ldq_11_bits_uop_frs3_en;
      5'b01100:
        casez_tmp_191 = ldq_12_bits_uop_frs3_en;
      5'b01101:
        casez_tmp_191 = ldq_13_bits_uop_frs3_en;
      5'b01110:
        casez_tmp_191 = ldq_14_bits_uop_frs3_en;
      5'b01111:
        casez_tmp_191 = ldq_15_bits_uop_frs3_en;
      5'b10000:
        casez_tmp_191 = ldq_16_bits_uop_frs3_en;
      5'b10001:
        casez_tmp_191 = ldq_17_bits_uop_frs3_en;
      5'b10010:
        casez_tmp_191 = ldq_18_bits_uop_frs3_en;
      5'b10011:
        casez_tmp_191 = ldq_19_bits_uop_frs3_en;
      5'b10100:
        casez_tmp_191 = ldq_20_bits_uop_frs3_en;
      5'b10101:
        casez_tmp_191 = ldq_21_bits_uop_frs3_en;
      5'b10110:
        casez_tmp_191 = ldq_22_bits_uop_frs3_en;
      5'b10111:
        casez_tmp_191 = ldq_23_bits_uop_frs3_en;
      5'b11000:
        casez_tmp_191 = ldq_24_bits_uop_frs3_en;
      5'b11001:
        casez_tmp_191 = ldq_25_bits_uop_frs3_en;
      5'b11010:
        casez_tmp_191 = ldq_26_bits_uop_frs3_en;
      5'b11011:
        casez_tmp_191 = ldq_27_bits_uop_frs3_en;
      5'b11100:
        casez_tmp_191 = ldq_28_bits_uop_frs3_en;
      5'b11101:
        casez_tmp_191 = ldq_29_bits_uop_frs3_en;
      5'b11110:
        casez_tmp_191 = ldq_30_bits_uop_frs3_en;
      default:
        casez_tmp_191 = ldq_31_bits_uop_frs3_en;
    endcase
  end // always @(*)
  reg         casez_tmp_192;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_192 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_192 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_192 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_192 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_192 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_192 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_192 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_192 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_192 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_192 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_192 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_192 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_192 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_192 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_192 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_192 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_192 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_192 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_192 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_192 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_192 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_192 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_192 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_192 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_192 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_192 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_192 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_192 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_192 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_192 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_192 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_192 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  reg         casez_tmp_193;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_193 = ldq_0_bits_uop_fp_single;
      5'b00001:
        casez_tmp_193 = ldq_1_bits_uop_fp_single;
      5'b00010:
        casez_tmp_193 = ldq_2_bits_uop_fp_single;
      5'b00011:
        casez_tmp_193 = ldq_3_bits_uop_fp_single;
      5'b00100:
        casez_tmp_193 = ldq_4_bits_uop_fp_single;
      5'b00101:
        casez_tmp_193 = ldq_5_bits_uop_fp_single;
      5'b00110:
        casez_tmp_193 = ldq_6_bits_uop_fp_single;
      5'b00111:
        casez_tmp_193 = ldq_7_bits_uop_fp_single;
      5'b01000:
        casez_tmp_193 = ldq_8_bits_uop_fp_single;
      5'b01001:
        casez_tmp_193 = ldq_9_bits_uop_fp_single;
      5'b01010:
        casez_tmp_193 = ldq_10_bits_uop_fp_single;
      5'b01011:
        casez_tmp_193 = ldq_11_bits_uop_fp_single;
      5'b01100:
        casez_tmp_193 = ldq_12_bits_uop_fp_single;
      5'b01101:
        casez_tmp_193 = ldq_13_bits_uop_fp_single;
      5'b01110:
        casez_tmp_193 = ldq_14_bits_uop_fp_single;
      5'b01111:
        casez_tmp_193 = ldq_15_bits_uop_fp_single;
      5'b10000:
        casez_tmp_193 = ldq_16_bits_uop_fp_single;
      5'b10001:
        casez_tmp_193 = ldq_17_bits_uop_fp_single;
      5'b10010:
        casez_tmp_193 = ldq_18_bits_uop_fp_single;
      5'b10011:
        casez_tmp_193 = ldq_19_bits_uop_fp_single;
      5'b10100:
        casez_tmp_193 = ldq_20_bits_uop_fp_single;
      5'b10101:
        casez_tmp_193 = ldq_21_bits_uop_fp_single;
      5'b10110:
        casez_tmp_193 = ldq_22_bits_uop_fp_single;
      5'b10111:
        casez_tmp_193 = ldq_23_bits_uop_fp_single;
      5'b11000:
        casez_tmp_193 = ldq_24_bits_uop_fp_single;
      5'b11001:
        casez_tmp_193 = ldq_25_bits_uop_fp_single;
      5'b11010:
        casez_tmp_193 = ldq_26_bits_uop_fp_single;
      5'b11011:
        casez_tmp_193 = ldq_27_bits_uop_fp_single;
      5'b11100:
        casez_tmp_193 = ldq_28_bits_uop_fp_single;
      5'b11101:
        casez_tmp_193 = ldq_29_bits_uop_fp_single;
      5'b11110:
        casez_tmp_193 = ldq_30_bits_uop_fp_single;
      default:
        casez_tmp_193 = ldq_31_bits_uop_fp_single;
    endcase
  end // always @(*)
  reg         casez_tmp_194;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_194 = ldq_0_bits_uop_xcpt_pf_if;
      5'b00001:
        casez_tmp_194 = ldq_1_bits_uop_xcpt_pf_if;
      5'b00010:
        casez_tmp_194 = ldq_2_bits_uop_xcpt_pf_if;
      5'b00011:
        casez_tmp_194 = ldq_3_bits_uop_xcpt_pf_if;
      5'b00100:
        casez_tmp_194 = ldq_4_bits_uop_xcpt_pf_if;
      5'b00101:
        casez_tmp_194 = ldq_5_bits_uop_xcpt_pf_if;
      5'b00110:
        casez_tmp_194 = ldq_6_bits_uop_xcpt_pf_if;
      5'b00111:
        casez_tmp_194 = ldq_7_bits_uop_xcpt_pf_if;
      5'b01000:
        casez_tmp_194 = ldq_8_bits_uop_xcpt_pf_if;
      5'b01001:
        casez_tmp_194 = ldq_9_bits_uop_xcpt_pf_if;
      5'b01010:
        casez_tmp_194 = ldq_10_bits_uop_xcpt_pf_if;
      5'b01011:
        casez_tmp_194 = ldq_11_bits_uop_xcpt_pf_if;
      5'b01100:
        casez_tmp_194 = ldq_12_bits_uop_xcpt_pf_if;
      5'b01101:
        casez_tmp_194 = ldq_13_bits_uop_xcpt_pf_if;
      5'b01110:
        casez_tmp_194 = ldq_14_bits_uop_xcpt_pf_if;
      5'b01111:
        casez_tmp_194 = ldq_15_bits_uop_xcpt_pf_if;
      5'b10000:
        casez_tmp_194 = ldq_16_bits_uop_xcpt_pf_if;
      5'b10001:
        casez_tmp_194 = ldq_17_bits_uop_xcpt_pf_if;
      5'b10010:
        casez_tmp_194 = ldq_18_bits_uop_xcpt_pf_if;
      5'b10011:
        casez_tmp_194 = ldq_19_bits_uop_xcpt_pf_if;
      5'b10100:
        casez_tmp_194 = ldq_20_bits_uop_xcpt_pf_if;
      5'b10101:
        casez_tmp_194 = ldq_21_bits_uop_xcpt_pf_if;
      5'b10110:
        casez_tmp_194 = ldq_22_bits_uop_xcpt_pf_if;
      5'b10111:
        casez_tmp_194 = ldq_23_bits_uop_xcpt_pf_if;
      5'b11000:
        casez_tmp_194 = ldq_24_bits_uop_xcpt_pf_if;
      5'b11001:
        casez_tmp_194 = ldq_25_bits_uop_xcpt_pf_if;
      5'b11010:
        casez_tmp_194 = ldq_26_bits_uop_xcpt_pf_if;
      5'b11011:
        casez_tmp_194 = ldq_27_bits_uop_xcpt_pf_if;
      5'b11100:
        casez_tmp_194 = ldq_28_bits_uop_xcpt_pf_if;
      5'b11101:
        casez_tmp_194 = ldq_29_bits_uop_xcpt_pf_if;
      5'b11110:
        casez_tmp_194 = ldq_30_bits_uop_xcpt_pf_if;
      default:
        casez_tmp_194 = ldq_31_bits_uop_xcpt_pf_if;
    endcase
  end // always @(*)
  reg         casez_tmp_195;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_195 = ldq_0_bits_uop_xcpt_ae_if;
      5'b00001:
        casez_tmp_195 = ldq_1_bits_uop_xcpt_ae_if;
      5'b00010:
        casez_tmp_195 = ldq_2_bits_uop_xcpt_ae_if;
      5'b00011:
        casez_tmp_195 = ldq_3_bits_uop_xcpt_ae_if;
      5'b00100:
        casez_tmp_195 = ldq_4_bits_uop_xcpt_ae_if;
      5'b00101:
        casez_tmp_195 = ldq_5_bits_uop_xcpt_ae_if;
      5'b00110:
        casez_tmp_195 = ldq_6_bits_uop_xcpt_ae_if;
      5'b00111:
        casez_tmp_195 = ldq_7_bits_uop_xcpt_ae_if;
      5'b01000:
        casez_tmp_195 = ldq_8_bits_uop_xcpt_ae_if;
      5'b01001:
        casez_tmp_195 = ldq_9_bits_uop_xcpt_ae_if;
      5'b01010:
        casez_tmp_195 = ldq_10_bits_uop_xcpt_ae_if;
      5'b01011:
        casez_tmp_195 = ldq_11_bits_uop_xcpt_ae_if;
      5'b01100:
        casez_tmp_195 = ldq_12_bits_uop_xcpt_ae_if;
      5'b01101:
        casez_tmp_195 = ldq_13_bits_uop_xcpt_ae_if;
      5'b01110:
        casez_tmp_195 = ldq_14_bits_uop_xcpt_ae_if;
      5'b01111:
        casez_tmp_195 = ldq_15_bits_uop_xcpt_ae_if;
      5'b10000:
        casez_tmp_195 = ldq_16_bits_uop_xcpt_ae_if;
      5'b10001:
        casez_tmp_195 = ldq_17_bits_uop_xcpt_ae_if;
      5'b10010:
        casez_tmp_195 = ldq_18_bits_uop_xcpt_ae_if;
      5'b10011:
        casez_tmp_195 = ldq_19_bits_uop_xcpt_ae_if;
      5'b10100:
        casez_tmp_195 = ldq_20_bits_uop_xcpt_ae_if;
      5'b10101:
        casez_tmp_195 = ldq_21_bits_uop_xcpt_ae_if;
      5'b10110:
        casez_tmp_195 = ldq_22_bits_uop_xcpt_ae_if;
      5'b10111:
        casez_tmp_195 = ldq_23_bits_uop_xcpt_ae_if;
      5'b11000:
        casez_tmp_195 = ldq_24_bits_uop_xcpt_ae_if;
      5'b11001:
        casez_tmp_195 = ldq_25_bits_uop_xcpt_ae_if;
      5'b11010:
        casez_tmp_195 = ldq_26_bits_uop_xcpt_ae_if;
      5'b11011:
        casez_tmp_195 = ldq_27_bits_uop_xcpt_ae_if;
      5'b11100:
        casez_tmp_195 = ldq_28_bits_uop_xcpt_ae_if;
      5'b11101:
        casez_tmp_195 = ldq_29_bits_uop_xcpt_ae_if;
      5'b11110:
        casez_tmp_195 = ldq_30_bits_uop_xcpt_ae_if;
      default:
        casez_tmp_195 = ldq_31_bits_uop_xcpt_ae_if;
    endcase
  end // always @(*)
  reg         casez_tmp_196;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_196 = ldq_0_bits_uop_xcpt_ma_if;
      5'b00001:
        casez_tmp_196 = ldq_1_bits_uop_xcpt_ma_if;
      5'b00010:
        casez_tmp_196 = ldq_2_bits_uop_xcpt_ma_if;
      5'b00011:
        casez_tmp_196 = ldq_3_bits_uop_xcpt_ma_if;
      5'b00100:
        casez_tmp_196 = ldq_4_bits_uop_xcpt_ma_if;
      5'b00101:
        casez_tmp_196 = ldq_5_bits_uop_xcpt_ma_if;
      5'b00110:
        casez_tmp_196 = ldq_6_bits_uop_xcpt_ma_if;
      5'b00111:
        casez_tmp_196 = ldq_7_bits_uop_xcpt_ma_if;
      5'b01000:
        casez_tmp_196 = ldq_8_bits_uop_xcpt_ma_if;
      5'b01001:
        casez_tmp_196 = ldq_9_bits_uop_xcpt_ma_if;
      5'b01010:
        casez_tmp_196 = ldq_10_bits_uop_xcpt_ma_if;
      5'b01011:
        casez_tmp_196 = ldq_11_bits_uop_xcpt_ma_if;
      5'b01100:
        casez_tmp_196 = ldq_12_bits_uop_xcpt_ma_if;
      5'b01101:
        casez_tmp_196 = ldq_13_bits_uop_xcpt_ma_if;
      5'b01110:
        casez_tmp_196 = ldq_14_bits_uop_xcpt_ma_if;
      5'b01111:
        casez_tmp_196 = ldq_15_bits_uop_xcpt_ma_if;
      5'b10000:
        casez_tmp_196 = ldq_16_bits_uop_xcpt_ma_if;
      5'b10001:
        casez_tmp_196 = ldq_17_bits_uop_xcpt_ma_if;
      5'b10010:
        casez_tmp_196 = ldq_18_bits_uop_xcpt_ma_if;
      5'b10011:
        casez_tmp_196 = ldq_19_bits_uop_xcpt_ma_if;
      5'b10100:
        casez_tmp_196 = ldq_20_bits_uop_xcpt_ma_if;
      5'b10101:
        casez_tmp_196 = ldq_21_bits_uop_xcpt_ma_if;
      5'b10110:
        casez_tmp_196 = ldq_22_bits_uop_xcpt_ma_if;
      5'b10111:
        casez_tmp_196 = ldq_23_bits_uop_xcpt_ma_if;
      5'b11000:
        casez_tmp_196 = ldq_24_bits_uop_xcpt_ma_if;
      5'b11001:
        casez_tmp_196 = ldq_25_bits_uop_xcpt_ma_if;
      5'b11010:
        casez_tmp_196 = ldq_26_bits_uop_xcpt_ma_if;
      5'b11011:
        casez_tmp_196 = ldq_27_bits_uop_xcpt_ma_if;
      5'b11100:
        casez_tmp_196 = ldq_28_bits_uop_xcpt_ma_if;
      5'b11101:
        casez_tmp_196 = ldq_29_bits_uop_xcpt_ma_if;
      5'b11110:
        casez_tmp_196 = ldq_30_bits_uop_xcpt_ma_if;
      default:
        casez_tmp_196 = ldq_31_bits_uop_xcpt_ma_if;
    endcase
  end // always @(*)
  reg         casez_tmp_197;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_197 = ldq_0_bits_uop_bp_debug_if;
      5'b00001:
        casez_tmp_197 = ldq_1_bits_uop_bp_debug_if;
      5'b00010:
        casez_tmp_197 = ldq_2_bits_uop_bp_debug_if;
      5'b00011:
        casez_tmp_197 = ldq_3_bits_uop_bp_debug_if;
      5'b00100:
        casez_tmp_197 = ldq_4_bits_uop_bp_debug_if;
      5'b00101:
        casez_tmp_197 = ldq_5_bits_uop_bp_debug_if;
      5'b00110:
        casez_tmp_197 = ldq_6_bits_uop_bp_debug_if;
      5'b00111:
        casez_tmp_197 = ldq_7_bits_uop_bp_debug_if;
      5'b01000:
        casez_tmp_197 = ldq_8_bits_uop_bp_debug_if;
      5'b01001:
        casez_tmp_197 = ldq_9_bits_uop_bp_debug_if;
      5'b01010:
        casez_tmp_197 = ldq_10_bits_uop_bp_debug_if;
      5'b01011:
        casez_tmp_197 = ldq_11_bits_uop_bp_debug_if;
      5'b01100:
        casez_tmp_197 = ldq_12_bits_uop_bp_debug_if;
      5'b01101:
        casez_tmp_197 = ldq_13_bits_uop_bp_debug_if;
      5'b01110:
        casez_tmp_197 = ldq_14_bits_uop_bp_debug_if;
      5'b01111:
        casez_tmp_197 = ldq_15_bits_uop_bp_debug_if;
      5'b10000:
        casez_tmp_197 = ldq_16_bits_uop_bp_debug_if;
      5'b10001:
        casez_tmp_197 = ldq_17_bits_uop_bp_debug_if;
      5'b10010:
        casez_tmp_197 = ldq_18_bits_uop_bp_debug_if;
      5'b10011:
        casez_tmp_197 = ldq_19_bits_uop_bp_debug_if;
      5'b10100:
        casez_tmp_197 = ldq_20_bits_uop_bp_debug_if;
      5'b10101:
        casez_tmp_197 = ldq_21_bits_uop_bp_debug_if;
      5'b10110:
        casez_tmp_197 = ldq_22_bits_uop_bp_debug_if;
      5'b10111:
        casez_tmp_197 = ldq_23_bits_uop_bp_debug_if;
      5'b11000:
        casez_tmp_197 = ldq_24_bits_uop_bp_debug_if;
      5'b11001:
        casez_tmp_197 = ldq_25_bits_uop_bp_debug_if;
      5'b11010:
        casez_tmp_197 = ldq_26_bits_uop_bp_debug_if;
      5'b11011:
        casez_tmp_197 = ldq_27_bits_uop_bp_debug_if;
      5'b11100:
        casez_tmp_197 = ldq_28_bits_uop_bp_debug_if;
      5'b11101:
        casez_tmp_197 = ldq_29_bits_uop_bp_debug_if;
      5'b11110:
        casez_tmp_197 = ldq_30_bits_uop_bp_debug_if;
      default:
        casez_tmp_197 = ldq_31_bits_uop_bp_debug_if;
    endcase
  end // always @(*)
  reg         casez_tmp_198;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_198 = ldq_0_bits_uop_bp_xcpt_if;
      5'b00001:
        casez_tmp_198 = ldq_1_bits_uop_bp_xcpt_if;
      5'b00010:
        casez_tmp_198 = ldq_2_bits_uop_bp_xcpt_if;
      5'b00011:
        casez_tmp_198 = ldq_3_bits_uop_bp_xcpt_if;
      5'b00100:
        casez_tmp_198 = ldq_4_bits_uop_bp_xcpt_if;
      5'b00101:
        casez_tmp_198 = ldq_5_bits_uop_bp_xcpt_if;
      5'b00110:
        casez_tmp_198 = ldq_6_bits_uop_bp_xcpt_if;
      5'b00111:
        casez_tmp_198 = ldq_7_bits_uop_bp_xcpt_if;
      5'b01000:
        casez_tmp_198 = ldq_8_bits_uop_bp_xcpt_if;
      5'b01001:
        casez_tmp_198 = ldq_9_bits_uop_bp_xcpt_if;
      5'b01010:
        casez_tmp_198 = ldq_10_bits_uop_bp_xcpt_if;
      5'b01011:
        casez_tmp_198 = ldq_11_bits_uop_bp_xcpt_if;
      5'b01100:
        casez_tmp_198 = ldq_12_bits_uop_bp_xcpt_if;
      5'b01101:
        casez_tmp_198 = ldq_13_bits_uop_bp_xcpt_if;
      5'b01110:
        casez_tmp_198 = ldq_14_bits_uop_bp_xcpt_if;
      5'b01111:
        casez_tmp_198 = ldq_15_bits_uop_bp_xcpt_if;
      5'b10000:
        casez_tmp_198 = ldq_16_bits_uop_bp_xcpt_if;
      5'b10001:
        casez_tmp_198 = ldq_17_bits_uop_bp_xcpt_if;
      5'b10010:
        casez_tmp_198 = ldq_18_bits_uop_bp_xcpt_if;
      5'b10011:
        casez_tmp_198 = ldq_19_bits_uop_bp_xcpt_if;
      5'b10100:
        casez_tmp_198 = ldq_20_bits_uop_bp_xcpt_if;
      5'b10101:
        casez_tmp_198 = ldq_21_bits_uop_bp_xcpt_if;
      5'b10110:
        casez_tmp_198 = ldq_22_bits_uop_bp_xcpt_if;
      5'b10111:
        casez_tmp_198 = ldq_23_bits_uop_bp_xcpt_if;
      5'b11000:
        casez_tmp_198 = ldq_24_bits_uop_bp_xcpt_if;
      5'b11001:
        casez_tmp_198 = ldq_25_bits_uop_bp_xcpt_if;
      5'b11010:
        casez_tmp_198 = ldq_26_bits_uop_bp_xcpt_if;
      5'b11011:
        casez_tmp_198 = ldq_27_bits_uop_bp_xcpt_if;
      5'b11100:
        casez_tmp_198 = ldq_28_bits_uop_bp_xcpt_if;
      5'b11101:
        casez_tmp_198 = ldq_29_bits_uop_bp_xcpt_if;
      5'b11110:
        casez_tmp_198 = ldq_30_bits_uop_bp_xcpt_if;
      default:
        casez_tmp_198 = ldq_31_bits_uop_bp_xcpt_if;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_199;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_199 = ldq_0_bits_uop_debug_fsrc;
      5'b00001:
        casez_tmp_199 = ldq_1_bits_uop_debug_fsrc;
      5'b00010:
        casez_tmp_199 = ldq_2_bits_uop_debug_fsrc;
      5'b00011:
        casez_tmp_199 = ldq_3_bits_uop_debug_fsrc;
      5'b00100:
        casez_tmp_199 = ldq_4_bits_uop_debug_fsrc;
      5'b00101:
        casez_tmp_199 = ldq_5_bits_uop_debug_fsrc;
      5'b00110:
        casez_tmp_199 = ldq_6_bits_uop_debug_fsrc;
      5'b00111:
        casez_tmp_199 = ldq_7_bits_uop_debug_fsrc;
      5'b01000:
        casez_tmp_199 = ldq_8_bits_uop_debug_fsrc;
      5'b01001:
        casez_tmp_199 = ldq_9_bits_uop_debug_fsrc;
      5'b01010:
        casez_tmp_199 = ldq_10_bits_uop_debug_fsrc;
      5'b01011:
        casez_tmp_199 = ldq_11_bits_uop_debug_fsrc;
      5'b01100:
        casez_tmp_199 = ldq_12_bits_uop_debug_fsrc;
      5'b01101:
        casez_tmp_199 = ldq_13_bits_uop_debug_fsrc;
      5'b01110:
        casez_tmp_199 = ldq_14_bits_uop_debug_fsrc;
      5'b01111:
        casez_tmp_199 = ldq_15_bits_uop_debug_fsrc;
      5'b10000:
        casez_tmp_199 = ldq_16_bits_uop_debug_fsrc;
      5'b10001:
        casez_tmp_199 = ldq_17_bits_uop_debug_fsrc;
      5'b10010:
        casez_tmp_199 = ldq_18_bits_uop_debug_fsrc;
      5'b10011:
        casez_tmp_199 = ldq_19_bits_uop_debug_fsrc;
      5'b10100:
        casez_tmp_199 = ldq_20_bits_uop_debug_fsrc;
      5'b10101:
        casez_tmp_199 = ldq_21_bits_uop_debug_fsrc;
      5'b10110:
        casez_tmp_199 = ldq_22_bits_uop_debug_fsrc;
      5'b10111:
        casez_tmp_199 = ldq_23_bits_uop_debug_fsrc;
      5'b11000:
        casez_tmp_199 = ldq_24_bits_uop_debug_fsrc;
      5'b11001:
        casez_tmp_199 = ldq_25_bits_uop_debug_fsrc;
      5'b11010:
        casez_tmp_199 = ldq_26_bits_uop_debug_fsrc;
      5'b11011:
        casez_tmp_199 = ldq_27_bits_uop_debug_fsrc;
      5'b11100:
        casez_tmp_199 = ldq_28_bits_uop_debug_fsrc;
      5'b11101:
        casez_tmp_199 = ldq_29_bits_uop_debug_fsrc;
      5'b11110:
        casez_tmp_199 = ldq_30_bits_uop_debug_fsrc;
      default:
        casez_tmp_199 = ldq_31_bits_uop_debug_fsrc;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_200;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_200 = ldq_0_bits_uop_debug_tsrc;
      5'b00001:
        casez_tmp_200 = ldq_1_bits_uop_debug_tsrc;
      5'b00010:
        casez_tmp_200 = ldq_2_bits_uop_debug_tsrc;
      5'b00011:
        casez_tmp_200 = ldq_3_bits_uop_debug_tsrc;
      5'b00100:
        casez_tmp_200 = ldq_4_bits_uop_debug_tsrc;
      5'b00101:
        casez_tmp_200 = ldq_5_bits_uop_debug_tsrc;
      5'b00110:
        casez_tmp_200 = ldq_6_bits_uop_debug_tsrc;
      5'b00111:
        casez_tmp_200 = ldq_7_bits_uop_debug_tsrc;
      5'b01000:
        casez_tmp_200 = ldq_8_bits_uop_debug_tsrc;
      5'b01001:
        casez_tmp_200 = ldq_9_bits_uop_debug_tsrc;
      5'b01010:
        casez_tmp_200 = ldq_10_bits_uop_debug_tsrc;
      5'b01011:
        casez_tmp_200 = ldq_11_bits_uop_debug_tsrc;
      5'b01100:
        casez_tmp_200 = ldq_12_bits_uop_debug_tsrc;
      5'b01101:
        casez_tmp_200 = ldq_13_bits_uop_debug_tsrc;
      5'b01110:
        casez_tmp_200 = ldq_14_bits_uop_debug_tsrc;
      5'b01111:
        casez_tmp_200 = ldq_15_bits_uop_debug_tsrc;
      5'b10000:
        casez_tmp_200 = ldq_16_bits_uop_debug_tsrc;
      5'b10001:
        casez_tmp_200 = ldq_17_bits_uop_debug_tsrc;
      5'b10010:
        casez_tmp_200 = ldq_18_bits_uop_debug_tsrc;
      5'b10011:
        casez_tmp_200 = ldq_19_bits_uop_debug_tsrc;
      5'b10100:
        casez_tmp_200 = ldq_20_bits_uop_debug_tsrc;
      5'b10101:
        casez_tmp_200 = ldq_21_bits_uop_debug_tsrc;
      5'b10110:
        casez_tmp_200 = ldq_22_bits_uop_debug_tsrc;
      5'b10111:
        casez_tmp_200 = ldq_23_bits_uop_debug_tsrc;
      5'b11000:
        casez_tmp_200 = ldq_24_bits_uop_debug_tsrc;
      5'b11001:
        casez_tmp_200 = ldq_25_bits_uop_debug_tsrc;
      5'b11010:
        casez_tmp_200 = ldq_26_bits_uop_debug_tsrc;
      5'b11011:
        casez_tmp_200 = ldq_27_bits_uop_debug_tsrc;
      5'b11100:
        casez_tmp_200 = ldq_28_bits_uop_debug_tsrc;
      5'b11101:
        casez_tmp_200 = ldq_29_bits_uop_debug_tsrc;
      5'b11110:
        casez_tmp_200 = ldq_30_bits_uop_debug_tsrc;
      default:
        casez_tmp_200 = ldq_31_bits_uop_debug_tsrc;
    endcase
  end // always @(*)
  reg         casez_tmp_201;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_201 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_201 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_201 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_201 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_201 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_201 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_201 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_201 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_201 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_201 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_201 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_201 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_201 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_201 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_201 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_201 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_201 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_201 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_201 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_201 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_201 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_201 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_201 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_201 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_201 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_201 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_201 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_201 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_201 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_201 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_201 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_201 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_202;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_202 = ldq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_202 = ldq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_202 = ldq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_202 = ldq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_202 = ldq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_202 = ldq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_202 = ldq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_202 = ldq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_202 = ldq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_202 = ldq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_202 = ldq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_202 = ldq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_202 = ldq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_202 = ldq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_202 = ldq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_202 = ldq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_202 = ldq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_202 = ldq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_202 = ldq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_202 = ldq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_202 = ldq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_202 = ldq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_202 = ldq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_202 = ldq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_202 = ldq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_202 = ldq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_202 = ldq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_202 = ldq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_202 = ldq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_202 = ldq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_202 = ldq_30_bits_addr_bits;
      default:
        casez_tmp_202 = ldq_31_bits_addr_bits;
    endcase
  end // always @(*)
  reg         casez_tmp_203;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_203 = ldq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_203 = ldq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_203 = ldq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_203 = ldq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_203 = ldq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_203 = ldq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_203 = ldq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_203 = ldq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_203 = ldq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_203 = ldq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_203 = ldq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_203 = ldq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_203 = ldq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_203 = ldq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_203 = ldq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_203 = ldq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_203 = ldq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_203 = ldq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_203 = ldq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_203 = ldq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_203 = ldq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_203 = ldq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_203 = ldq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_203 = ldq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_203 = ldq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_203 = ldq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_203 = ldq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_203 = ldq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_203 = ldq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_203 = ldq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_203 = ldq_30_bits_addr_is_virtual;
      default:
        casez_tmp_203 = ldq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         casez_tmp_204;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_204 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_204 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_204 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_204 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_204 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_204 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_204 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_204 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_204 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_204 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_204 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_204 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_204 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_204 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_204 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_204 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_204 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_204 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_204 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_204 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_204 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_204 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_204 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_204 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_204 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_204 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_204 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_204 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_204 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_204 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_204 = ldq_30_bits_executed;
      default:
        casez_tmp_204 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg         casez_tmp_205;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_205 = ldq_0_bits_order_fail;
      5'b00001:
        casez_tmp_205 = ldq_1_bits_order_fail;
      5'b00010:
        casez_tmp_205 = ldq_2_bits_order_fail;
      5'b00011:
        casez_tmp_205 = ldq_3_bits_order_fail;
      5'b00100:
        casez_tmp_205 = ldq_4_bits_order_fail;
      5'b00101:
        casez_tmp_205 = ldq_5_bits_order_fail;
      5'b00110:
        casez_tmp_205 = ldq_6_bits_order_fail;
      5'b00111:
        casez_tmp_205 = ldq_7_bits_order_fail;
      5'b01000:
        casez_tmp_205 = ldq_8_bits_order_fail;
      5'b01001:
        casez_tmp_205 = ldq_9_bits_order_fail;
      5'b01010:
        casez_tmp_205 = ldq_10_bits_order_fail;
      5'b01011:
        casez_tmp_205 = ldq_11_bits_order_fail;
      5'b01100:
        casez_tmp_205 = ldq_12_bits_order_fail;
      5'b01101:
        casez_tmp_205 = ldq_13_bits_order_fail;
      5'b01110:
        casez_tmp_205 = ldq_14_bits_order_fail;
      5'b01111:
        casez_tmp_205 = ldq_15_bits_order_fail;
      5'b10000:
        casez_tmp_205 = ldq_16_bits_order_fail;
      5'b10001:
        casez_tmp_205 = ldq_17_bits_order_fail;
      5'b10010:
        casez_tmp_205 = ldq_18_bits_order_fail;
      5'b10011:
        casez_tmp_205 = ldq_19_bits_order_fail;
      5'b10100:
        casez_tmp_205 = ldq_20_bits_order_fail;
      5'b10101:
        casez_tmp_205 = ldq_21_bits_order_fail;
      5'b10110:
        casez_tmp_205 = ldq_22_bits_order_fail;
      5'b10111:
        casez_tmp_205 = ldq_23_bits_order_fail;
      5'b11000:
        casez_tmp_205 = ldq_24_bits_order_fail;
      5'b11001:
        casez_tmp_205 = ldq_25_bits_order_fail;
      5'b11010:
        casez_tmp_205 = ldq_26_bits_order_fail;
      5'b11011:
        casez_tmp_205 = ldq_27_bits_order_fail;
      5'b11100:
        casez_tmp_205 = ldq_28_bits_order_fail;
      5'b11101:
        casez_tmp_205 = ldq_29_bits_order_fail;
      5'b11110:
        casez_tmp_205 = ldq_30_bits_order_fail;
      default:
        casez_tmp_205 = ldq_31_bits_order_fail;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_206;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_206 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_206 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_206 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_206 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_206 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_206 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_206 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_206 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_206 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_206 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_206 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_206 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_206 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_206 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_206 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_206 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_206 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_206 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_206 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_206 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_206 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_206 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_206 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_206 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_206 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_206 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_206 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_206 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_206 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_206 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_206 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_206 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  reg         casez_tmp_207;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_207 = p1_block_load_mask_0;
      5'b00001:
        casez_tmp_207 = p1_block_load_mask_1;
      5'b00010:
        casez_tmp_207 = p1_block_load_mask_2;
      5'b00011:
        casez_tmp_207 = p1_block_load_mask_3;
      5'b00100:
        casez_tmp_207 = p1_block_load_mask_4;
      5'b00101:
        casez_tmp_207 = p1_block_load_mask_5;
      5'b00110:
        casez_tmp_207 = p1_block_load_mask_6;
      5'b00111:
        casez_tmp_207 = p1_block_load_mask_7;
      5'b01000:
        casez_tmp_207 = p1_block_load_mask_8;
      5'b01001:
        casez_tmp_207 = p1_block_load_mask_9;
      5'b01010:
        casez_tmp_207 = p1_block_load_mask_10;
      5'b01011:
        casez_tmp_207 = p1_block_load_mask_11;
      5'b01100:
        casez_tmp_207 = p1_block_load_mask_12;
      5'b01101:
        casez_tmp_207 = p1_block_load_mask_13;
      5'b01110:
        casez_tmp_207 = p1_block_load_mask_14;
      5'b01111:
        casez_tmp_207 = p1_block_load_mask_15;
      5'b10000:
        casez_tmp_207 = p1_block_load_mask_16;
      5'b10001:
        casez_tmp_207 = p1_block_load_mask_17;
      5'b10010:
        casez_tmp_207 = p1_block_load_mask_18;
      5'b10011:
        casez_tmp_207 = p1_block_load_mask_19;
      5'b10100:
        casez_tmp_207 = p1_block_load_mask_20;
      5'b10101:
        casez_tmp_207 = p1_block_load_mask_21;
      5'b10110:
        casez_tmp_207 = p1_block_load_mask_22;
      5'b10111:
        casez_tmp_207 = p1_block_load_mask_23;
      5'b11000:
        casez_tmp_207 = p1_block_load_mask_24;
      5'b11001:
        casez_tmp_207 = p1_block_load_mask_25;
      5'b11010:
        casez_tmp_207 = p1_block_load_mask_26;
      5'b11011:
        casez_tmp_207 = p1_block_load_mask_27;
      5'b11100:
        casez_tmp_207 = p1_block_load_mask_28;
      5'b11101:
        casez_tmp_207 = p1_block_load_mask_29;
      5'b11110:
        casez_tmp_207 = p1_block_load_mask_30;
      default:
        casez_tmp_207 = p1_block_load_mask_31;
    endcase
  end // always @(*)
  reg         casez_tmp_208;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_208 = p2_block_load_mask_0;
      5'b00001:
        casez_tmp_208 = p2_block_load_mask_1;
      5'b00010:
        casez_tmp_208 = p2_block_load_mask_2;
      5'b00011:
        casez_tmp_208 = p2_block_load_mask_3;
      5'b00100:
        casez_tmp_208 = p2_block_load_mask_4;
      5'b00101:
        casez_tmp_208 = p2_block_load_mask_5;
      5'b00110:
        casez_tmp_208 = p2_block_load_mask_6;
      5'b00111:
        casez_tmp_208 = p2_block_load_mask_7;
      5'b01000:
        casez_tmp_208 = p2_block_load_mask_8;
      5'b01001:
        casez_tmp_208 = p2_block_load_mask_9;
      5'b01010:
        casez_tmp_208 = p2_block_load_mask_10;
      5'b01011:
        casez_tmp_208 = p2_block_load_mask_11;
      5'b01100:
        casez_tmp_208 = p2_block_load_mask_12;
      5'b01101:
        casez_tmp_208 = p2_block_load_mask_13;
      5'b01110:
        casez_tmp_208 = p2_block_load_mask_14;
      5'b01111:
        casez_tmp_208 = p2_block_load_mask_15;
      5'b10000:
        casez_tmp_208 = p2_block_load_mask_16;
      5'b10001:
        casez_tmp_208 = p2_block_load_mask_17;
      5'b10010:
        casez_tmp_208 = p2_block_load_mask_18;
      5'b10011:
        casez_tmp_208 = p2_block_load_mask_19;
      5'b10100:
        casez_tmp_208 = p2_block_load_mask_20;
      5'b10101:
        casez_tmp_208 = p2_block_load_mask_21;
      5'b10110:
        casez_tmp_208 = p2_block_load_mask_22;
      5'b10111:
        casez_tmp_208 = p2_block_load_mask_23;
      5'b11000:
        casez_tmp_208 = p2_block_load_mask_24;
      5'b11001:
        casez_tmp_208 = p2_block_load_mask_25;
      5'b11010:
        casez_tmp_208 = p2_block_load_mask_26;
      5'b11011:
        casez_tmp_208 = p2_block_load_mask_27;
      5'b11100:
        casez_tmp_208 = p2_block_load_mask_28;
      5'b11101:
        casez_tmp_208 = p2_block_load_mask_29;
      5'b11110:
        casez_tmp_208 = p2_block_load_mask_30;
      default:
        casez_tmp_208 = p2_block_load_mask_31;
    endcase
  end // always @(*)
  reg         can_fire_load_retry_REG_1;
  reg         casez_tmp_209;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_209 = stq_0_valid;
      5'b00001:
        casez_tmp_209 = stq_1_valid;
      5'b00010:
        casez_tmp_209 = stq_2_valid;
      5'b00011:
        casez_tmp_209 = stq_3_valid;
      5'b00100:
        casez_tmp_209 = stq_4_valid;
      5'b00101:
        casez_tmp_209 = stq_5_valid;
      5'b00110:
        casez_tmp_209 = stq_6_valid;
      5'b00111:
        casez_tmp_209 = stq_7_valid;
      5'b01000:
        casez_tmp_209 = stq_8_valid;
      5'b01001:
        casez_tmp_209 = stq_9_valid;
      5'b01010:
        casez_tmp_209 = stq_10_valid;
      5'b01011:
        casez_tmp_209 = stq_11_valid;
      5'b01100:
        casez_tmp_209 = stq_12_valid;
      5'b01101:
        casez_tmp_209 = stq_13_valid;
      5'b01110:
        casez_tmp_209 = stq_14_valid;
      5'b01111:
        casez_tmp_209 = stq_15_valid;
      5'b10000:
        casez_tmp_209 = stq_16_valid;
      5'b10001:
        casez_tmp_209 = stq_17_valid;
      5'b10010:
        casez_tmp_209 = stq_18_valid;
      5'b10011:
        casez_tmp_209 = stq_19_valid;
      5'b10100:
        casez_tmp_209 = stq_20_valid;
      5'b10101:
        casez_tmp_209 = stq_21_valid;
      5'b10110:
        casez_tmp_209 = stq_22_valid;
      5'b10111:
        casez_tmp_209 = stq_23_valid;
      5'b11000:
        casez_tmp_209 = stq_24_valid;
      5'b11001:
        casez_tmp_209 = stq_25_valid;
      5'b11010:
        casez_tmp_209 = stq_26_valid;
      5'b11011:
        casez_tmp_209 = stq_27_valid;
      5'b11100:
        casez_tmp_209 = stq_28_valid;
      5'b11101:
        casez_tmp_209 = stq_29_valid;
      5'b11110:
        casez_tmp_209 = stq_30_valid;
      default:
        casez_tmp_209 = stq_31_valid;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_210;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_210 = stq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_210 = stq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_210 = stq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_210 = stq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_210 = stq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_210 = stq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_210 = stq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_210 = stq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_210 = stq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_210 = stq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_210 = stq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_210 = stq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_210 = stq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_210 = stq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_210 = stq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_210 = stq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_210 = stq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_210 = stq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_210 = stq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_210 = stq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_210 = stq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_210 = stq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_210 = stq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_210 = stq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_210 = stq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_210 = stq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_210 = stq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_210 = stq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_210 = stq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_210 = stq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_210 = stq_30_bits_uop_uopc;
      default:
        casez_tmp_210 = stq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_211;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_211 = stq_0_bits_uop_inst;
      5'b00001:
        casez_tmp_211 = stq_1_bits_uop_inst;
      5'b00010:
        casez_tmp_211 = stq_2_bits_uop_inst;
      5'b00011:
        casez_tmp_211 = stq_3_bits_uop_inst;
      5'b00100:
        casez_tmp_211 = stq_4_bits_uop_inst;
      5'b00101:
        casez_tmp_211 = stq_5_bits_uop_inst;
      5'b00110:
        casez_tmp_211 = stq_6_bits_uop_inst;
      5'b00111:
        casez_tmp_211 = stq_7_bits_uop_inst;
      5'b01000:
        casez_tmp_211 = stq_8_bits_uop_inst;
      5'b01001:
        casez_tmp_211 = stq_9_bits_uop_inst;
      5'b01010:
        casez_tmp_211 = stq_10_bits_uop_inst;
      5'b01011:
        casez_tmp_211 = stq_11_bits_uop_inst;
      5'b01100:
        casez_tmp_211 = stq_12_bits_uop_inst;
      5'b01101:
        casez_tmp_211 = stq_13_bits_uop_inst;
      5'b01110:
        casez_tmp_211 = stq_14_bits_uop_inst;
      5'b01111:
        casez_tmp_211 = stq_15_bits_uop_inst;
      5'b10000:
        casez_tmp_211 = stq_16_bits_uop_inst;
      5'b10001:
        casez_tmp_211 = stq_17_bits_uop_inst;
      5'b10010:
        casez_tmp_211 = stq_18_bits_uop_inst;
      5'b10011:
        casez_tmp_211 = stq_19_bits_uop_inst;
      5'b10100:
        casez_tmp_211 = stq_20_bits_uop_inst;
      5'b10101:
        casez_tmp_211 = stq_21_bits_uop_inst;
      5'b10110:
        casez_tmp_211 = stq_22_bits_uop_inst;
      5'b10111:
        casez_tmp_211 = stq_23_bits_uop_inst;
      5'b11000:
        casez_tmp_211 = stq_24_bits_uop_inst;
      5'b11001:
        casez_tmp_211 = stq_25_bits_uop_inst;
      5'b11010:
        casez_tmp_211 = stq_26_bits_uop_inst;
      5'b11011:
        casez_tmp_211 = stq_27_bits_uop_inst;
      5'b11100:
        casez_tmp_211 = stq_28_bits_uop_inst;
      5'b11101:
        casez_tmp_211 = stq_29_bits_uop_inst;
      5'b11110:
        casez_tmp_211 = stq_30_bits_uop_inst;
      default:
        casez_tmp_211 = stq_31_bits_uop_inst;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_212;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_212 = stq_0_bits_uop_debug_inst;
      5'b00001:
        casez_tmp_212 = stq_1_bits_uop_debug_inst;
      5'b00010:
        casez_tmp_212 = stq_2_bits_uop_debug_inst;
      5'b00011:
        casez_tmp_212 = stq_3_bits_uop_debug_inst;
      5'b00100:
        casez_tmp_212 = stq_4_bits_uop_debug_inst;
      5'b00101:
        casez_tmp_212 = stq_5_bits_uop_debug_inst;
      5'b00110:
        casez_tmp_212 = stq_6_bits_uop_debug_inst;
      5'b00111:
        casez_tmp_212 = stq_7_bits_uop_debug_inst;
      5'b01000:
        casez_tmp_212 = stq_8_bits_uop_debug_inst;
      5'b01001:
        casez_tmp_212 = stq_9_bits_uop_debug_inst;
      5'b01010:
        casez_tmp_212 = stq_10_bits_uop_debug_inst;
      5'b01011:
        casez_tmp_212 = stq_11_bits_uop_debug_inst;
      5'b01100:
        casez_tmp_212 = stq_12_bits_uop_debug_inst;
      5'b01101:
        casez_tmp_212 = stq_13_bits_uop_debug_inst;
      5'b01110:
        casez_tmp_212 = stq_14_bits_uop_debug_inst;
      5'b01111:
        casez_tmp_212 = stq_15_bits_uop_debug_inst;
      5'b10000:
        casez_tmp_212 = stq_16_bits_uop_debug_inst;
      5'b10001:
        casez_tmp_212 = stq_17_bits_uop_debug_inst;
      5'b10010:
        casez_tmp_212 = stq_18_bits_uop_debug_inst;
      5'b10011:
        casez_tmp_212 = stq_19_bits_uop_debug_inst;
      5'b10100:
        casez_tmp_212 = stq_20_bits_uop_debug_inst;
      5'b10101:
        casez_tmp_212 = stq_21_bits_uop_debug_inst;
      5'b10110:
        casez_tmp_212 = stq_22_bits_uop_debug_inst;
      5'b10111:
        casez_tmp_212 = stq_23_bits_uop_debug_inst;
      5'b11000:
        casez_tmp_212 = stq_24_bits_uop_debug_inst;
      5'b11001:
        casez_tmp_212 = stq_25_bits_uop_debug_inst;
      5'b11010:
        casez_tmp_212 = stq_26_bits_uop_debug_inst;
      5'b11011:
        casez_tmp_212 = stq_27_bits_uop_debug_inst;
      5'b11100:
        casez_tmp_212 = stq_28_bits_uop_debug_inst;
      5'b11101:
        casez_tmp_212 = stq_29_bits_uop_debug_inst;
      5'b11110:
        casez_tmp_212 = stq_30_bits_uop_debug_inst;
      default:
        casez_tmp_212 = stq_31_bits_uop_debug_inst;
    endcase
  end // always @(*)
  reg         casez_tmp_213;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_213 = stq_0_bits_uop_is_rvc;
      5'b00001:
        casez_tmp_213 = stq_1_bits_uop_is_rvc;
      5'b00010:
        casez_tmp_213 = stq_2_bits_uop_is_rvc;
      5'b00011:
        casez_tmp_213 = stq_3_bits_uop_is_rvc;
      5'b00100:
        casez_tmp_213 = stq_4_bits_uop_is_rvc;
      5'b00101:
        casez_tmp_213 = stq_5_bits_uop_is_rvc;
      5'b00110:
        casez_tmp_213 = stq_6_bits_uop_is_rvc;
      5'b00111:
        casez_tmp_213 = stq_7_bits_uop_is_rvc;
      5'b01000:
        casez_tmp_213 = stq_8_bits_uop_is_rvc;
      5'b01001:
        casez_tmp_213 = stq_9_bits_uop_is_rvc;
      5'b01010:
        casez_tmp_213 = stq_10_bits_uop_is_rvc;
      5'b01011:
        casez_tmp_213 = stq_11_bits_uop_is_rvc;
      5'b01100:
        casez_tmp_213 = stq_12_bits_uop_is_rvc;
      5'b01101:
        casez_tmp_213 = stq_13_bits_uop_is_rvc;
      5'b01110:
        casez_tmp_213 = stq_14_bits_uop_is_rvc;
      5'b01111:
        casez_tmp_213 = stq_15_bits_uop_is_rvc;
      5'b10000:
        casez_tmp_213 = stq_16_bits_uop_is_rvc;
      5'b10001:
        casez_tmp_213 = stq_17_bits_uop_is_rvc;
      5'b10010:
        casez_tmp_213 = stq_18_bits_uop_is_rvc;
      5'b10011:
        casez_tmp_213 = stq_19_bits_uop_is_rvc;
      5'b10100:
        casez_tmp_213 = stq_20_bits_uop_is_rvc;
      5'b10101:
        casez_tmp_213 = stq_21_bits_uop_is_rvc;
      5'b10110:
        casez_tmp_213 = stq_22_bits_uop_is_rvc;
      5'b10111:
        casez_tmp_213 = stq_23_bits_uop_is_rvc;
      5'b11000:
        casez_tmp_213 = stq_24_bits_uop_is_rvc;
      5'b11001:
        casez_tmp_213 = stq_25_bits_uop_is_rvc;
      5'b11010:
        casez_tmp_213 = stq_26_bits_uop_is_rvc;
      5'b11011:
        casez_tmp_213 = stq_27_bits_uop_is_rvc;
      5'b11100:
        casez_tmp_213 = stq_28_bits_uop_is_rvc;
      5'b11101:
        casez_tmp_213 = stq_29_bits_uop_is_rvc;
      5'b11110:
        casez_tmp_213 = stq_30_bits_uop_is_rvc;
      default:
        casez_tmp_213 = stq_31_bits_uop_is_rvc;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_214;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_214 = stq_0_bits_uop_debug_pc;
      5'b00001:
        casez_tmp_214 = stq_1_bits_uop_debug_pc;
      5'b00010:
        casez_tmp_214 = stq_2_bits_uop_debug_pc;
      5'b00011:
        casez_tmp_214 = stq_3_bits_uop_debug_pc;
      5'b00100:
        casez_tmp_214 = stq_4_bits_uop_debug_pc;
      5'b00101:
        casez_tmp_214 = stq_5_bits_uop_debug_pc;
      5'b00110:
        casez_tmp_214 = stq_6_bits_uop_debug_pc;
      5'b00111:
        casez_tmp_214 = stq_7_bits_uop_debug_pc;
      5'b01000:
        casez_tmp_214 = stq_8_bits_uop_debug_pc;
      5'b01001:
        casez_tmp_214 = stq_9_bits_uop_debug_pc;
      5'b01010:
        casez_tmp_214 = stq_10_bits_uop_debug_pc;
      5'b01011:
        casez_tmp_214 = stq_11_bits_uop_debug_pc;
      5'b01100:
        casez_tmp_214 = stq_12_bits_uop_debug_pc;
      5'b01101:
        casez_tmp_214 = stq_13_bits_uop_debug_pc;
      5'b01110:
        casez_tmp_214 = stq_14_bits_uop_debug_pc;
      5'b01111:
        casez_tmp_214 = stq_15_bits_uop_debug_pc;
      5'b10000:
        casez_tmp_214 = stq_16_bits_uop_debug_pc;
      5'b10001:
        casez_tmp_214 = stq_17_bits_uop_debug_pc;
      5'b10010:
        casez_tmp_214 = stq_18_bits_uop_debug_pc;
      5'b10011:
        casez_tmp_214 = stq_19_bits_uop_debug_pc;
      5'b10100:
        casez_tmp_214 = stq_20_bits_uop_debug_pc;
      5'b10101:
        casez_tmp_214 = stq_21_bits_uop_debug_pc;
      5'b10110:
        casez_tmp_214 = stq_22_bits_uop_debug_pc;
      5'b10111:
        casez_tmp_214 = stq_23_bits_uop_debug_pc;
      5'b11000:
        casez_tmp_214 = stq_24_bits_uop_debug_pc;
      5'b11001:
        casez_tmp_214 = stq_25_bits_uop_debug_pc;
      5'b11010:
        casez_tmp_214 = stq_26_bits_uop_debug_pc;
      5'b11011:
        casez_tmp_214 = stq_27_bits_uop_debug_pc;
      5'b11100:
        casez_tmp_214 = stq_28_bits_uop_debug_pc;
      5'b11101:
        casez_tmp_214 = stq_29_bits_uop_debug_pc;
      5'b11110:
        casez_tmp_214 = stq_30_bits_uop_debug_pc;
      default:
        casez_tmp_214 = stq_31_bits_uop_debug_pc;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_215;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_215 = stq_0_bits_uop_iq_type;
      5'b00001:
        casez_tmp_215 = stq_1_bits_uop_iq_type;
      5'b00010:
        casez_tmp_215 = stq_2_bits_uop_iq_type;
      5'b00011:
        casez_tmp_215 = stq_3_bits_uop_iq_type;
      5'b00100:
        casez_tmp_215 = stq_4_bits_uop_iq_type;
      5'b00101:
        casez_tmp_215 = stq_5_bits_uop_iq_type;
      5'b00110:
        casez_tmp_215 = stq_6_bits_uop_iq_type;
      5'b00111:
        casez_tmp_215 = stq_7_bits_uop_iq_type;
      5'b01000:
        casez_tmp_215 = stq_8_bits_uop_iq_type;
      5'b01001:
        casez_tmp_215 = stq_9_bits_uop_iq_type;
      5'b01010:
        casez_tmp_215 = stq_10_bits_uop_iq_type;
      5'b01011:
        casez_tmp_215 = stq_11_bits_uop_iq_type;
      5'b01100:
        casez_tmp_215 = stq_12_bits_uop_iq_type;
      5'b01101:
        casez_tmp_215 = stq_13_bits_uop_iq_type;
      5'b01110:
        casez_tmp_215 = stq_14_bits_uop_iq_type;
      5'b01111:
        casez_tmp_215 = stq_15_bits_uop_iq_type;
      5'b10000:
        casez_tmp_215 = stq_16_bits_uop_iq_type;
      5'b10001:
        casez_tmp_215 = stq_17_bits_uop_iq_type;
      5'b10010:
        casez_tmp_215 = stq_18_bits_uop_iq_type;
      5'b10011:
        casez_tmp_215 = stq_19_bits_uop_iq_type;
      5'b10100:
        casez_tmp_215 = stq_20_bits_uop_iq_type;
      5'b10101:
        casez_tmp_215 = stq_21_bits_uop_iq_type;
      5'b10110:
        casez_tmp_215 = stq_22_bits_uop_iq_type;
      5'b10111:
        casez_tmp_215 = stq_23_bits_uop_iq_type;
      5'b11000:
        casez_tmp_215 = stq_24_bits_uop_iq_type;
      5'b11001:
        casez_tmp_215 = stq_25_bits_uop_iq_type;
      5'b11010:
        casez_tmp_215 = stq_26_bits_uop_iq_type;
      5'b11011:
        casez_tmp_215 = stq_27_bits_uop_iq_type;
      5'b11100:
        casez_tmp_215 = stq_28_bits_uop_iq_type;
      5'b11101:
        casez_tmp_215 = stq_29_bits_uop_iq_type;
      5'b11110:
        casez_tmp_215 = stq_30_bits_uop_iq_type;
      default:
        casez_tmp_215 = stq_31_bits_uop_iq_type;
    endcase
  end // always @(*)
  reg  [9:0]  casez_tmp_216;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_216 = stq_0_bits_uop_fu_code;
      5'b00001:
        casez_tmp_216 = stq_1_bits_uop_fu_code;
      5'b00010:
        casez_tmp_216 = stq_2_bits_uop_fu_code;
      5'b00011:
        casez_tmp_216 = stq_3_bits_uop_fu_code;
      5'b00100:
        casez_tmp_216 = stq_4_bits_uop_fu_code;
      5'b00101:
        casez_tmp_216 = stq_5_bits_uop_fu_code;
      5'b00110:
        casez_tmp_216 = stq_6_bits_uop_fu_code;
      5'b00111:
        casez_tmp_216 = stq_7_bits_uop_fu_code;
      5'b01000:
        casez_tmp_216 = stq_8_bits_uop_fu_code;
      5'b01001:
        casez_tmp_216 = stq_9_bits_uop_fu_code;
      5'b01010:
        casez_tmp_216 = stq_10_bits_uop_fu_code;
      5'b01011:
        casez_tmp_216 = stq_11_bits_uop_fu_code;
      5'b01100:
        casez_tmp_216 = stq_12_bits_uop_fu_code;
      5'b01101:
        casez_tmp_216 = stq_13_bits_uop_fu_code;
      5'b01110:
        casez_tmp_216 = stq_14_bits_uop_fu_code;
      5'b01111:
        casez_tmp_216 = stq_15_bits_uop_fu_code;
      5'b10000:
        casez_tmp_216 = stq_16_bits_uop_fu_code;
      5'b10001:
        casez_tmp_216 = stq_17_bits_uop_fu_code;
      5'b10010:
        casez_tmp_216 = stq_18_bits_uop_fu_code;
      5'b10011:
        casez_tmp_216 = stq_19_bits_uop_fu_code;
      5'b10100:
        casez_tmp_216 = stq_20_bits_uop_fu_code;
      5'b10101:
        casez_tmp_216 = stq_21_bits_uop_fu_code;
      5'b10110:
        casez_tmp_216 = stq_22_bits_uop_fu_code;
      5'b10111:
        casez_tmp_216 = stq_23_bits_uop_fu_code;
      5'b11000:
        casez_tmp_216 = stq_24_bits_uop_fu_code;
      5'b11001:
        casez_tmp_216 = stq_25_bits_uop_fu_code;
      5'b11010:
        casez_tmp_216 = stq_26_bits_uop_fu_code;
      5'b11011:
        casez_tmp_216 = stq_27_bits_uop_fu_code;
      5'b11100:
        casez_tmp_216 = stq_28_bits_uop_fu_code;
      5'b11101:
        casez_tmp_216 = stq_29_bits_uop_fu_code;
      5'b11110:
        casez_tmp_216 = stq_30_bits_uop_fu_code;
      default:
        casez_tmp_216 = stq_31_bits_uop_fu_code;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_217;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_217 = stq_0_bits_uop_ctrl_br_type;
      5'b00001:
        casez_tmp_217 = stq_1_bits_uop_ctrl_br_type;
      5'b00010:
        casez_tmp_217 = stq_2_bits_uop_ctrl_br_type;
      5'b00011:
        casez_tmp_217 = stq_3_bits_uop_ctrl_br_type;
      5'b00100:
        casez_tmp_217 = stq_4_bits_uop_ctrl_br_type;
      5'b00101:
        casez_tmp_217 = stq_5_bits_uop_ctrl_br_type;
      5'b00110:
        casez_tmp_217 = stq_6_bits_uop_ctrl_br_type;
      5'b00111:
        casez_tmp_217 = stq_7_bits_uop_ctrl_br_type;
      5'b01000:
        casez_tmp_217 = stq_8_bits_uop_ctrl_br_type;
      5'b01001:
        casez_tmp_217 = stq_9_bits_uop_ctrl_br_type;
      5'b01010:
        casez_tmp_217 = stq_10_bits_uop_ctrl_br_type;
      5'b01011:
        casez_tmp_217 = stq_11_bits_uop_ctrl_br_type;
      5'b01100:
        casez_tmp_217 = stq_12_bits_uop_ctrl_br_type;
      5'b01101:
        casez_tmp_217 = stq_13_bits_uop_ctrl_br_type;
      5'b01110:
        casez_tmp_217 = stq_14_bits_uop_ctrl_br_type;
      5'b01111:
        casez_tmp_217 = stq_15_bits_uop_ctrl_br_type;
      5'b10000:
        casez_tmp_217 = stq_16_bits_uop_ctrl_br_type;
      5'b10001:
        casez_tmp_217 = stq_17_bits_uop_ctrl_br_type;
      5'b10010:
        casez_tmp_217 = stq_18_bits_uop_ctrl_br_type;
      5'b10011:
        casez_tmp_217 = stq_19_bits_uop_ctrl_br_type;
      5'b10100:
        casez_tmp_217 = stq_20_bits_uop_ctrl_br_type;
      5'b10101:
        casez_tmp_217 = stq_21_bits_uop_ctrl_br_type;
      5'b10110:
        casez_tmp_217 = stq_22_bits_uop_ctrl_br_type;
      5'b10111:
        casez_tmp_217 = stq_23_bits_uop_ctrl_br_type;
      5'b11000:
        casez_tmp_217 = stq_24_bits_uop_ctrl_br_type;
      5'b11001:
        casez_tmp_217 = stq_25_bits_uop_ctrl_br_type;
      5'b11010:
        casez_tmp_217 = stq_26_bits_uop_ctrl_br_type;
      5'b11011:
        casez_tmp_217 = stq_27_bits_uop_ctrl_br_type;
      5'b11100:
        casez_tmp_217 = stq_28_bits_uop_ctrl_br_type;
      5'b11101:
        casez_tmp_217 = stq_29_bits_uop_ctrl_br_type;
      5'b11110:
        casez_tmp_217 = stq_30_bits_uop_ctrl_br_type;
      default:
        casez_tmp_217 = stq_31_bits_uop_ctrl_br_type;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_218;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_218 = stq_0_bits_uop_ctrl_op1_sel;
      5'b00001:
        casez_tmp_218 = stq_1_bits_uop_ctrl_op1_sel;
      5'b00010:
        casez_tmp_218 = stq_2_bits_uop_ctrl_op1_sel;
      5'b00011:
        casez_tmp_218 = stq_3_bits_uop_ctrl_op1_sel;
      5'b00100:
        casez_tmp_218 = stq_4_bits_uop_ctrl_op1_sel;
      5'b00101:
        casez_tmp_218 = stq_5_bits_uop_ctrl_op1_sel;
      5'b00110:
        casez_tmp_218 = stq_6_bits_uop_ctrl_op1_sel;
      5'b00111:
        casez_tmp_218 = stq_7_bits_uop_ctrl_op1_sel;
      5'b01000:
        casez_tmp_218 = stq_8_bits_uop_ctrl_op1_sel;
      5'b01001:
        casez_tmp_218 = stq_9_bits_uop_ctrl_op1_sel;
      5'b01010:
        casez_tmp_218 = stq_10_bits_uop_ctrl_op1_sel;
      5'b01011:
        casez_tmp_218 = stq_11_bits_uop_ctrl_op1_sel;
      5'b01100:
        casez_tmp_218 = stq_12_bits_uop_ctrl_op1_sel;
      5'b01101:
        casez_tmp_218 = stq_13_bits_uop_ctrl_op1_sel;
      5'b01110:
        casez_tmp_218 = stq_14_bits_uop_ctrl_op1_sel;
      5'b01111:
        casez_tmp_218 = stq_15_bits_uop_ctrl_op1_sel;
      5'b10000:
        casez_tmp_218 = stq_16_bits_uop_ctrl_op1_sel;
      5'b10001:
        casez_tmp_218 = stq_17_bits_uop_ctrl_op1_sel;
      5'b10010:
        casez_tmp_218 = stq_18_bits_uop_ctrl_op1_sel;
      5'b10011:
        casez_tmp_218 = stq_19_bits_uop_ctrl_op1_sel;
      5'b10100:
        casez_tmp_218 = stq_20_bits_uop_ctrl_op1_sel;
      5'b10101:
        casez_tmp_218 = stq_21_bits_uop_ctrl_op1_sel;
      5'b10110:
        casez_tmp_218 = stq_22_bits_uop_ctrl_op1_sel;
      5'b10111:
        casez_tmp_218 = stq_23_bits_uop_ctrl_op1_sel;
      5'b11000:
        casez_tmp_218 = stq_24_bits_uop_ctrl_op1_sel;
      5'b11001:
        casez_tmp_218 = stq_25_bits_uop_ctrl_op1_sel;
      5'b11010:
        casez_tmp_218 = stq_26_bits_uop_ctrl_op1_sel;
      5'b11011:
        casez_tmp_218 = stq_27_bits_uop_ctrl_op1_sel;
      5'b11100:
        casez_tmp_218 = stq_28_bits_uop_ctrl_op1_sel;
      5'b11101:
        casez_tmp_218 = stq_29_bits_uop_ctrl_op1_sel;
      5'b11110:
        casez_tmp_218 = stq_30_bits_uop_ctrl_op1_sel;
      default:
        casez_tmp_218 = stq_31_bits_uop_ctrl_op1_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_219;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_219 = stq_0_bits_uop_ctrl_op2_sel;
      5'b00001:
        casez_tmp_219 = stq_1_bits_uop_ctrl_op2_sel;
      5'b00010:
        casez_tmp_219 = stq_2_bits_uop_ctrl_op2_sel;
      5'b00011:
        casez_tmp_219 = stq_3_bits_uop_ctrl_op2_sel;
      5'b00100:
        casez_tmp_219 = stq_4_bits_uop_ctrl_op2_sel;
      5'b00101:
        casez_tmp_219 = stq_5_bits_uop_ctrl_op2_sel;
      5'b00110:
        casez_tmp_219 = stq_6_bits_uop_ctrl_op2_sel;
      5'b00111:
        casez_tmp_219 = stq_7_bits_uop_ctrl_op2_sel;
      5'b01000:
        casez_tmp_219 = stq_8_bits_uop_ctrl_op2_sel;
      5'b01001:
        casez_tmp_219 = stq_9_bits_uop_ctrl_op2_sel;
      5'b01010:
        casez_tmp_219 = stq_10_bits_uop_ctrl_op2_sel;
      5'b01011:
        casez_tmp_219 = stq_11_bits_uop_ctrl_op2_sel;
      5'b01100:
        casez_tmp_219 = stq_12_bits_uop_ctrl_op2_sel;
      5'b01101:
        casez_tmp_219 = stq_13_bits_uop_ctrl_op2_sel;
      5'b01110:
        casez_tmp_219 = stq_14_bits_uop_ctrl_op2_sel;
      5'b01111:
        casez_tmp_219 = stq_15_bits_uop_ctrl_op2_sel;
      5'b10000:
        casez_tmp_219 = stq_16_bits_uop_ctrl_op2_sel;
      5'b10001:
        casez_tmp_219 = stq_17_bits_uop_ctrl_op2_sel;
      5'b10010:
        casez_tmp_219 = stq_18_bits_uop_ctrl_op2_sel;
      5'b10011:
        casez_tmp_219 = stq_19_bits_uop_ctrl_op2_sel;
      5'b10100:
        casez_tmp_219 = stq_20_bits_uop_ctrl_op2_sel;
      5'b10101:
        casez_tmp_219 = stq_21_bits_uop_ctrl_op2_sel;
      5'b10110:
        casez_tmp_219 = stq_22_bits_uop_ctrl_op2_sel;
      5'b10111:
        casez_tmp_219 = stq_23_bits_uop_ctrl_op2_sel;
      5'b11000:
        casez_tmp_219 = stq_24_bits_uop_ctrl_op2_sel;
      5'b11001:
        casez_tmp_219 = stq_25_bits_uop_ctrl_op2_sel;
      5'b11010:
        casez_tmp_219 = stq_26_bits_uop_ctrl_op2_sel;
      5'b11011:
        casez_tmp_219 = stq_27_bits_uop_ctrl_op2_sel;
      5'b11100:
        casez_tmp_219 = stq_28_bits_uop_ctrl_op2_sel;
      5'b11101:
        casez_tmp_219 = stq_29_bits_uop_ctrl_op2_sel;
      5'b11110:
        casez_tmp_219 = stq_30_bits_uop_ctrl_op2_sel;
      default:
        casez_tmp_219 = stq_31_bits_uop_ctrl_op2_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_220;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_220 = stq_0_bits_uop_ctrl_imm_sel;
      5'b00001:
        casez_tmp_220 = stq_1_bits_uop_ctrl_imm_sel;
      5'b00010:
        casez_tmp_220 = stq_2_bits_uop_ctrl_imm_sel;
      5'b00011:
        casez_tmp_220 = stq_3_bits_uop_ctrl_imm_sel;
      5'b00100:
        casez_tmp_220 = stq_4_bits_uop_ctrl_imm_sel;
      5'b00101:
        casez_tmp_220 = stq_5_bits_uop_ctrl_imm_sel;
      5'b00110:
        casez_tmp_220 = stq_6_bits_uop_ctrl_imm_sel;
      5'b00111:
        casez_tmp_220 = stq_7_bits_uop_ctrl_imm_sel;
      5'b01000:
        casez_tmp_220 = stq_8_bits_uop_ctrl_imm_sel;
      5'b01001:
        casez_tmp_220 = stq_9_bits_uop_ctrl_imm_sel;
      5'b01010:
        casez_tmp_220 = stq_10_bits_uop_ctrl_imm_sel;
      5'b01011:
        casez_tmp_220 = stq_11_bits_uop_ctrl_imm_sel;
      5'b01100:
        casez_tmp_220 = stq_12_bits_uop_ctrl_imm_sel;
      5'b01101:
        casez_tmp_220 = stq_13_bits_uop_ctrl_imm_sel;
      5'b01110:
        casez_tmp_220 = stq_14_bits_uop_ctrl_imm_sel;
      5'b01111:
        casez_tmp_220 = stq_15_bits_uop_ctrl_imm_sel;
      5'b10000:
        casez_tmp_220 = stq_16_bits_uop_ctrl_imm_sel;
      5'b10001:
        casez_tmp_220 = stq_17_bits_uop_ctrl_imm_sel;
      5'b10010:
        casez_tmp_220 = stq_18_bits_uop_ctrl_imm_sel;
      5'b10011:
        casez_tmp_220 = stq_19_bits_uop_ctrl_imm_sel;
      5'b10100:
        casez_tmp_220 = stq_20_bits_uop_ctrl_imm_sel;
      5'b10101:
        casez_tmp_220 = stq_21_bits_uop_ctrl_imm_sel;
      5'b10110:
        casez_tmp_220 = stq_22_bits_uop_ctrl_imm_sel;
      5'b10111:
        casez_tmp_220 = stq_23_bits_uop_ctrl_imm_sel;
      5'b11000:
        casez_tmp_220 = stq_24_bits_uop_ctrl_imm_sel;
      5'b11001:
        casez_tmp_220 = stq_25_bits_uop_ctrl_imm_sel;
      5'b11010:
        casez_tmp_220 = stq_26_bits_uop_ctrl_imm_sel;
      5'b11011:
        casez_tmp_220 = stq_27_bits_uop_ctrl_imm_sel;
      5'b11100:
        casez_tmp_220 = stq_28_bits_uop_ctrl_imm_sel;
      5'b11101:
        casez_tmp_220 = stq_29_bits_uop_ctrl_imm_sel;
      5'b11110:
        casez_tmp_220 = stq_30_bits_uop_ctrl_imm_sel;
      default:
        casez_tmp_220 = stq_31_bits_uop_ctrl_imm_sel;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_221;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_221 = stq_0_bits_uop_ctrl_op_fcn;
      5'b00001:
        casez_tmp_221 = stq_1_bits_uop_ctrl_op_fcn;
      5'b00010:
        casez_tmp_221 = stq_2_bits_uop_ctrl_op_fcn;
      5'b00011:
        casez_tmp_221 = stq_3_bits_uop_ctrl_op_fcn;
      5'b00100:
        casez_tmp_221 = stq_4_bits_uop_ctrl_op_fcn;
      5'b00101:
        casez_tmp_221 = stq_5_bits_uop_ctrl_op_fcn;
      5'b00110:
        casez_tmp_221 = stq_6_bits_uop_ctrl_op_fcn;
      5'b00111:
        casez_tmp_221 = stq_7_bits_uop_ctrl_op_fcn;
      5'b01000:
        casez_tmp_221 = stq_8_bits_uop_ctrl_op_fcn;
      5'b01001:
        casez_tmp_221 = stq_9_bits_uop_ctrl_op_fcn;
      5'b01010:
        casez_tmp_221 = stq_10_bits_uop_ctrl_op_fcn;
      5'b01011:
        casez_tmp_221 = stq_11_bits_uop_ctrl_op_fcn;
      5'b01100:
        casez_tmp_221 = stq_12_bits_uop_ctrl_op_fcn;
      5'b01101:
        casez_tmp_221 = stq_13_bits_uop_ctrl_op_fcn;
      5'b01110:
        casez_tmp_221 = stq_14_bits_uop_ctrl_op_fcn;
      5'b01111:
        casez_tmp_221 = stq_15_bits_uop_ctrl_op_fcn;
      5'b10000:
        casez_tmp_221 = stq_16_bits_uop_ctrl_op_fcn;
      5'b10001:
        casez_tmp_221 = stq_17_bits_uop_ctrl_op_fcn;
      5'b10010:
        casez_tmp_221 = stq_18_bits_uop_ctrl_op_fcn;
      5'b10011:
        casez_tmp_221 = stq_19_bits_uop_ctrl_op_fcn;
      5'b10100:
        casez_tmp_221 = stq_20_bits_uop_ctrl_op_fcn;
      5'b10101:
        casez_tmp_221 = stq_21_bits_uop_ctrl_op_fcn;
      5'b10110:
        casez_tmp_221 = stq_22_bits_uop_ctrl_op_fcn;
      5'b10111:
        casez_tmp_221 = stq_23_bits_uop_ctrl_op_fcn;
      5'b11000:
        casez_tmp_221 = stq_24_bits_uop_ctrl_op_fcn;
      5'b11001:
        casez_tmp_221 = stq_25_bits_uop_ctrl_op_fcn;
      5'b11010:
        casez_tmp_221 = stq_26_bits_uop_ctrl_op_fcn;
      5'b11011:
        casez_tmp_221 = stq_27_bits_uop_ctrl_op_fcn;
      5'b11100:
        casez_tmp_221 = stq_28_bits_uop_ctrl_op_fcn;
      5'b11101:
        casez_tmp_221 = stq_29_bits_uop_ctrl_op_fcn;
      5'b11110:
        casez_tmp_221 = stq_30_bits_uop_ctrl_op_fcn;
      default:
        casez_tmp_221 = stq_31_bits_uop_ctrl_op_fcn;
    endcase
  end // always @(*)
  reg         casez_tmp_222;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_222 = stq_0_bits_uop_ctrl_fcn_dw;
      5'b00001:
        casez_tmp_222 = stq_1_bits_uop_ctrl_fcn_dw;
      5'b00010:
        casez_tmp_222 = stq_2_bits_uop_ctrl_fcn_dw;
      5'b00011:
        casez_tmp_222 = stq_3_bits_uop_ctrl_fcn_dw;
      5'b00100:
        casez_tmp_222 = stq_4_bits_uop_ctrl_fcn_dw;
      5'b00101:
        casez_tmp_222 = stq_5_bits_uop_ctrl_fcn_dw;
      5'b00110:
        casez_tmp_222 = stq_6_bits_uop_ctrl_fcn_dw;
      5'b00111:
        casez_tmp_222 = stq_7_bits_uop_ctrl_fcn_dw;
      5'b01000:
        casez_tmp_222 = stq_8_bits_uop_ctrl_fcn_dw;
      5'b01001:
        casez_tmp_222 = stq_9_bits_uop_ctrl_fcn_dw;
      5'b01010:
        casez_tmp_222 = stq_10_bits_uop_ctrl_fcn_dw;
      5'b01011:
        casez_tmp_222 = stq_11_bits_uop_ctrl_fcn_dw;
      5'b01100:
        casez_tmp_222 = stq_12_bits_uop_ctrl_fcn_dw;
      5'b01101:
        casez_tmp_222 = stq_13_bits_uop_ctrl_fcn_dw;
      5'b01110:
        casez_tmp_222 = stq_14_bits_uop_ctrl_fcn_dw;
      5'b01111:
        casez_tmp_222 = stq_15_bits_uop_ctrl_fcn_dw;
      5'b10000:
        casez_tmp_222 = stq_16_bits_uop_ctrl_fcn_dw;
      5'b10001:
        casez_tmp_222 = stq_17_bits_uop_ctrl_fcn_dw;
      5'b10010:
        casez_tmp_222 = stq_18_bits_uop_ctrl_fcn_dw;
      5'b10011:
        casez_tmp_222 = stq_19_bits_uop_ctrl_fcn_dw;
      5'b10100:
        casez_tmp_222 = stq_20_bits_uop_ctrl_fcn_dw;
      5'b10101:
        casez_tmp_222 = stq_21_bits_uop_ctrl_fcn_dw;
      5'b10110:
        casez_tmp_222 = stq_22_bits_uop_ctrl_fcn_dw;
      5'b10111:
        casez_tmp_222 = stq_23_bits_uop_ctrl_fcn_dw;
      5'b11000:
        casez_tmp_222 = stq_24_bits_uop_ctrl_fcn_dw;
      5'b11001:
        casez_tmp_222 = stq_25_bits_uop_ctrl_fcn_dw;
      5'b11010:
        casez_tmp_222 = stq_26_bits_uop_ctrl_fcn_dw;
      5'b11011:
        casez_tmp_222 = stq_27_bits_uop_ctrl_fcn_dw;
      5'b11100:
        casez_tmp_222 = stq_28_bits_uop_ctrl_fcn_dw;
      5'b11101:
        casez_tmp_222 = stq_29_bits_uop_ctrl_fcn_dw;
      5'b11110:
        casez_tmp_222 = stq_30_bits_uop_ctrl_fcn_dw;
      default:
        casez_tmp_222 = stq_31_bits_uop_ctrl_fcn_dw;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_223;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_223 = stq_0_bits_uop_ctrl_csr_cmd;
      5'b00001:
        casez_tmp_223 = stq_1_bits_uop_ctrl_csr_cmd;
      5'b00010:
        casez_tmp_223 = stq_2_bits_uop_ctrl_csr_cmd;
      5'b00011:
        casez_tmp_223 = stq_3_bits_uop_ctrl_csr_cmd;
      5'b00100:
        casez_tmp_223 = stq_4_bits_uop_ctrl_csr_cmd;
      5'b00101:
        casez_tmp_223 = stq_5_bits_uop_ctrl_csr_cmd;
      5'b00110:
        casez_tmp_223 = stq_6_bits_uop_ctrl_csr_cmd;
      5'b00111:
        casez_tmp_223 = stq_7_bits_uop_ctrl_csr_cmd;
      5'b01000:
        casez_tmp_223 = stq_8_bits_uop_ctrl_csr_cmd;
      5'b01001:
        casez_tmp_223 = stq_9_bits_uop_ctrl_csr_cmd;
      5'b01010:
        casez_tmp_223 = stq_10_bits_uop_ctrl_csr_cmd;
      5'b01011:
        casez_tmp_223 = stq_11_bits_uop_ctrl_csr_cmd;
      5'b01100:
        casez_tmp_223 = stq_12_bits_uop_ctrl_csr_cmd;
      5'b01101:
        casez_tmp_223 = stq_13_bits_uop_ctrl_csr_cmd;
      5'b01110:
        casez_tmp_223 = stq_14_bits_uop_ctrl_csr_cmd;
      5'b01111:
        casez_tmp_223 = stq_15_bits_uop_ctrl_csr_cmd;
      5'b10000:
        casez_tmp_223 = stq_16_bits_uop_ctrl_csr_cmd;
      5'b10001:
        casez_tmp_223 = stq_17_bits_uop_ctrl_csr_cmd;
      5'b10010:
        casez_tmp_223 = stq_18_bits_uop_ctrl_csr_cmd;
      5'b10011:
        casez_tmp_223 = stq_19_bits_uop_ctrl_csr_cmd;
      5'b10100:
        casez_tmp_223 = stq_20_bits_uop_ctrl_csr_cmd;
      5'b10101:
        casez_tmp_223 = stq_21_bits_uop_ctrl_csr_cmd;
      5'b10110:
        casez_tmp_223 = stq_22_bits_uop_ctrl_csr_cmd;
      5'b10111:
        casez_tmp_223 = stq_23_bits_uop_ctrl_csr_cmd;
      5'b11000:
        casez_tmp_223 = stq_24_bits_uop_ctrl_csr_cmd;
      5'b11001:
        casez_tmp_223 = stq_25_bits_uop_ctrl_csr_cmd;
      5'b11010:
        casez_tmp_223 = stq_26_bits_uop_ctrl_csr_cmd;
      5'b11011:
        casez_tmp_223 = stq_27_bits_uop_ctrl_csr_cmd;
      5'b11100:
        casez_tmp_223 = stq_28_bits_uop_ctrl_csr_cmd;
      5'b11101:
        casez_tmp_223 = stq_29_bits_uop_ctrl_csr_cmd;
      5'b11110:
        casez_tmp_223 = stq_30_bits_uop_ctrl_csr_cmd;
      default:
        casez_tmp_223 = stq_31_bits_uop_ctrl_csr_cmd;
    endcase
  end // always @(*)
  reg         casez_tmp_224;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_224 = stq_0_bits_uop_ctrl_is_load;
      5'b00001:
        casez_tmp_224 = stq_1_bits_uop_ctrl_is_load;
      5'b00010:
        casez_tmp_224 = stq_2_bits_uop_ctrl_is_load;
      5'b00011:
        casez_tmp_224 = stq_3_bits_uop_ctrl_is_load;
      5'b00100:
        casez_tmp_224 = stq_4_bits_uop_ctrl_is_load;
      5'b00101:
        casez_tmp_224 = stq_5_bits_uop_ctrl_is_load;
      5'b00110:
        casez_tmp_224 = stq_6_bits_uop_ctrl_is_load;
      5'b00111:
        casez_tmp_224 = stq_7_bits_uop_ctrl_is_load;
      5'b01000:
        casez_tmp_224 = stq_8_bits_uop_ctrl_is_load;
      5'b01001:
        casez_tmp_224 = stq_9_bits_uop_ctrl_is_load;
      5'b01010:
        casez_tmp_224 = stq_10_bits_uop_ctrl_is_load;
      5'b01011:
        casez_tmp_224 = stq_11_bits_uop_ctrl_is_load;
      5'b01100:
        casez_tmp_224 = stq_12_bits_uop_ctrl_is_load;
      5'b01101:
        casez_tmp_224 = stq_13_bits_uop_ctrl_is_load;
      5'b01110:
        casez_tmp_224 = stq_14_bits_uop_ctrl_is_load;
      5'b01111:
        casez_tmp_224 = stq_15_bits_uop_ctrl_is_load;
      5'b10000:
        casez_tmp_224 = stq_16_bits_uop_ctrl_is_load;
      5'b10001:
        casez_tmp_224 = stq_17_bits_uop_ctrl_is_load;
      5'b10010:
        casez_tmp_224 = stq_18_bits_uop_ctrl_is_load;
      5'b10011:
        casez_tmp_224 = stq_19_bits_uop_ctrl_is_load;
      5'b10100:
        casez_tmp_224 = stq_20_bits_uop_ctrl_is_load;
      5'b10101:
        casez_tmp_224 = stq_21_bits_uop_ctrl_is_load;
      5'b10110:
        casez_tmp_224 = stq_22_bits_uop_ctrl_is_load;
      5'b10111:
        casez_tmp_224 = stq_23_bits_uop_ctrl_is_load;
      5'b11000:
        casez_tmp_224 = stq_24_bits_uop_ctrl_is_load;
      5'b11001:
        casez_tmp_224 = stq_25_bits_uop_ctrl_is_load;
      5'b11010:
        casez_tmp_224 = stq_26_bits_uop_ctrl_is_load;
      5'b11011:
        casez_tmp_224 = stq_27_bits_uop_ctrl_is_load;
      5'b11100:
        casez_tmp_224 = stq_28_bits_uop_ctrl_is_load;
      5'b11101:
        casez_tmp_224 = stq_29_bits_uop_ctrl_is_load;
      5'b11110:
        casez_tmp_224 = stq_30_bits_uop_ctrl_is_load;
      default:
        casez_tmp_224 = stq_31_bits_uop_ctrl_is_load;
    endcase
  end // always @(*)
  reg         casez_tmp_225;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_225 = stq_0_bits_uop_ctrl_is_sta;
      5'b00001:
        casez_tmp_225 = stq_1_bits_uop_ctrl_is_sta;
      5'b00010:
        casez_tmp_225 = stq_2_bits_uop_ctrl_is_sta;
      5'b00011:
        casez_tmp_225 = stq_3_bits_uop_ctrl_is_sta;
      5'b00100:
        casez_tmp_225 = stq_4_bits_uop_ctrl_is_sta;
      5'b00101:
        casez_tmp_225 = stq_5_bits_uop_ctrl_is_sta;
      5'b00110:
        casez_tmp_225 = stq_6_bits_uop_ctrl_is_sta;
      5'b00111:
        casez_tmp_225 = stq_7_bits_uop_ctrl_is_sta;
      5'b01000:
        casez_tmp_225 = stq_8_bits_uop_ctrl_is_sta;
      5'b01001:
        casez_tmp_225 = stq_9_bits_uop_ctrl_is_sta;
      5'b01010:
        casez_tmp_225 = stq_10_bits_uop_ctrl_is_sta;
      5'b01011:
        casez_tmp_225 = stq_11_bits_uop_ctrl_is_sta;
      5'b01100:
        casez_tmp_225 = stq_12_bits_uop_ctrl_is_sta;
      5'b01101:
        casez_tmp_225 = stq_13_bits_uop_ctrl_is_sta;
      5'b01110:
        casez_tmp_225 = stq_14_bits_uop_ctrl_is_sta;
      5'b01111:
        casez_tmp_225 = stq_15_bits_uop_ctrl_is_sta;
      5'b10000:
        casez_tmp_225 = stq_16_bits_uop_ctrl_is_sta;
      5'b10001:
        casez_tmp_225 = stq_17_bits_uop_ctrl_is_sta;
      5'b10010:
        casez_tmp_225 = stq_18_bits_uop_ctrl_is_sta;
      5'b10011:
        casez_tmp_225 = stq_19_bits_uop_ctrl_is_sta;
      5'b10100:
        casez_tmp_225 = stq_20_bits_uop_ctrl_is_sta;
      5'b10101:
        casez_tmp_225 = stq_21_bits_uop_ctrl_is_sta;
      5'b10110:
        casez_tmp_225 = stq_22_bits_uop_ctrl_is_sta;
      5'b10111:
        casez_tmp_225 = stq_23_bits_uop_ctrl_is_sta;
      5'b11000:
        casez_tmp_225 = stq_24_bits_uop_ctrl_is_sta;
      5'b11001:
        casez_tmp_225 = stq_25_bits_uop_ctrl_is_sta;
      5'b11010:
        casez_tmp_225 = stq_26_bits_uop_ctrl_is_sta;
      5'b11011:
        casez_tmp_225 = stq_27_bits_uop_ctrl_is_sta;
      5'b11100:
        casez_tmp_225 = stq_28_bits_uop_ctrl_is_sta;
      5'b11101:
        casez_tmp_225 = stq_29_bits_uop_ctrl_is_sta;
      5'b11110:
        casez_tmp_225 = stq_30_bits_uop_ctrl_is_sta;
      default:
        casez_tmp_225 = stq_31_bits_uop_ctrl_is_sta;
    endcase
  end // always @(*)
  reg         casez_tmp_226;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_226 = stq_0_bits_uop_ctrl_is_std;
      5'b00001:
        casez_tmp_226 = stq_1_bits_uop_ctrl_is_std;
      5'b00010:
        casez_tmp_226 = stq_2_bits_uop_ctrl_is_std;
      5'b00011:
        casez_tmp_226 = stq_3_bits_uop_ctrl_is_std;
      5'b00100:
        casez_tmp_226 = stq_4_bits_uop_ctrl_is_std;
      5'b00101:
        casez_tmp_226 = stq_5_bits_uop_ctrl_is_std;
      5'b00110:
        casez_tmp_226 = stq_6_bits_uop_ctrl_is_std;
      5'b00111:
        casez_tmp_226 = stq_7_bits_uop_ctrl_is_std;
      5'b01000:
        casez_tmp_226 = stq_8_bits_uop_ctrl_is_std;
      5'b01001:
        casez_tmp_226 = stq_9_bits_uop_ctrl_is_std;
      5'b01010:
        casez_tmp_226 = stq_10_bits_uop_ctrl_is_std;
      5'b01011:
        casez_tmp_226 = stq_11_bits_uop_ctrl_is_std;
      5'b01100:
        casez_tmp_226 = stq_12_bits_uop_ctrl_is_std;
      5'b01101:
        casez_tmp_226 = stq_13_bits_uop_ctrl_is_std;
      5'b01110:
        casez_tmp_226 = stq_14_bits_uop_ctrl_is_std;
      5'b01111:
        casez_tmp_226 = stq_15_bits_uop_ctrl_is_std;
      5'b10000:
        casez_tmp_226 = stq_16_bits_uop_ctrl_is_std;
      5'b10001:
        casez_tmp_226 = stq_17_bits_uop_ctrl_is_std;
      5'b10010:
        casez_tmp_226 = stq_18_bits_uop_ctrl_is_std;
      5'b10011:
        casez_tmp_226 = stq_19_bits_uop_ctrl_is_std;
      5'b10100:
        casez_tmp_226 = stq_20_bits_uop_ctrl_is_std;
      5'b10101:
        casez_tmp_226 = stq_21_bits_uop_ctrl_is_std;
      5'b10110:
        casez_tmp_226 = stq_22_bits_uop_ctrl_is_std;
      5'b10111:
        casez_tmp_226 = stq_23_bits_uop_ctrl_is_std;
      5'b11000:
        casez_tmp_226 = stq_24_bits_uop_ctrl_is_std;
      5'b11001:
        casez_tmp_226 = stq_25_bits_uop_ctrl_is_std;
      5'b11010:
        casez_tmp_226 = stq_26_bits_uop_ctrl_is_std;
      5'b11011:
        casez_tmp_226 = stq_27_bits_uop_ctrl_is_std;
      5'b11100:
        casez_tmp_226 = stq_28_bits_uop_ctrl_is_std;
      5'b11101:
        casez_tmp_226 = stq_29_bits_uop_ctrl_is_std;
      5'b11110:
        casez_tmp_226 = stq_30_bits_uop_ctrl_is_std;
      default:
        casez_tmp_226 = stq_31_bits_uop_ctrl_is_std;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_227;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_227 = stq_0_bits_uop_iw_state;
      5'b00001:
        casez_tmp_227 = stq_1_bits_uop_iw_state;
      5'b00010:
        casez_tmp_227 = stq_2_bits_uop_iw_state;
      5'b00011:
        casez_tmp_227 = stq_3_bits_uop_iw_state;
      5'b00100:
        casez_tmp_227 = stq_4_bits_uop_iw_state;
      5'b00101:
        casez_tmp_227 = stq_5_bits_uop_iw_state;
      5'b00110:
        casez_tmp_227 = stq_6_bits_uop_iw_state;
      5'b00111:
        casez_tmp_227 = stq_7_bits_uop_iw_state;
      5'b01000:
        casez_tmp_227 = stq_8_bits_uop_iw_state;
      5'b01001:
        casez_tmp_227 = stq_9_bits_uop_iw_state;
      5'b01010:
        casez_tmp_227 = stq_10_bits_uop_iw_state;
      5'b01011:
        casez_tmp_227 = stq_11_bits_uop_iw_state;
      5'b01100:
        casez_tmp_227 = stq_12_bits_uop_iw_state;
      5'b01101:
        casez_tmp_227 = stq_13_bits_uop_iw_state;
      5'b01110:
        casez_tmp_227 = stq_14_bits_uop_iw_state;
      5'b01111:
        casez_tmp_227 = stq_15_bits_uop_iw_state;
      5'b10000:
        casez_tmp_227 = stq_16_bits_uop_iw_state;
      5'b10001:
        casez_tmp_227 = stq_17_bits_uop_iw_state;
      5'b10010:
        casez_tmp_227 = stq_18_bits_uop_iw_state;
      5'b10011:
        casez_tmp_227 = stq_19_bits_uop_iw_state;
      5'b10100:
        casez_tmp_227 = stq_20_bits_uop_iw_state;
      5'b10101:
        casez_tmp_227 = stq_21_bits_uop_iw_state;
      5'b10110:
        casez_tmp_227 = stq_22_bits_uop_iw_state;
      5'b10111:
        casez_tmp_227 = stq_23_bits_uop_iw_state;
      5'b11000:
        casez_tmp_227 = stq_24_bits_uop_iw_state;
      5'b11001:
        casez_tmp_227 = stq_25_bits_uop_iw_state;
      5'b11010:
        casez_tmp_227 = stq_26_bits_uop_iw_state;
      5'b11011:
        casez_tmp_227 = stq_27_bits_uop_iw_state;
      5'b11100:
        casez_tmp_227 = stq_28_bits_uop_iw_state;
      5'b11101:
        casez_tmp_227 = stq_29_bits_uop_iw_state;
      5'b11110:
        casez_tmp_227 = stq_30_bits_uop_iw_state;
      default:
        casez_tmp_227 = stq_31_bits_uop_iw_state;
    endcase
  end // always @(*)
  reg         casez_tmp_228;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_228 = stq_0_bits_uop_iw_p1_poisoned;
      5'b00001:
        casez_tmp_228 = stq_1_bits_uop_iw_p1_poisoned;
      5'b00010:
        casez_tmp_228 = stq_2_bits_uop_iw_p1_poisoned;
      5'b00011:
        casez_tmp_228 = stq_3_bits_uop_iw_p1_poisoned;
      5'b00100:
        casez_tmp_228 = stq_4_bits_uop_iw_p1_poisoned;
      5'b00101:
        casez_tmp_228 = stq_5_bits_uop_iw_p1_poisoned;
      5'b00110:
        casez_tmp_228 = stq_6_bits_uop_iw_p1_poisoned;
      5'b00111:
        casez_tmp_228 = stq_7_bits_uop_iw_p1_poisoned;
      5'b01000:
        casez_tmp_228 = stq_8_bits_uop_iw_p1_poisoned;
      5'b01001:
        casez_tmp_228 = stq_9_bits_uop_iw_p1_poisoned;
      5'b01010:
        casez_tmp_228 = stq_10_bits_uop_iw_p1_poisoned;
      5'b01011:
        casez_tmp_228 = stq_11_bits_uop_iw_p1_poisoned;
      5'b01100:
        casez_tmp_228 = stq_12_bits_uop_iw_p1_poisoned;
      5'b01101:
        casez_tmp_228 = stq_13_bits_uop_iw_p1_poisoned;
      5'b01110:
        casez_tmp_228 = stq_14_bits_uop_iw_p1_poisoned;
      5'b01111:
        casez_tmp_228 = stq_15_bits_uop_iw_p1_poisoned;
      5'b10000:
        casez_tmp_228 = stq_16_bits_uop_iw_p1_poisoned;
      5'b10001:
        casez_tmp_228 = stq_17_bits_uop_iw_p1_poisoned;
      5'b10010:
        casez_tmp_228 = stq_18_bits_uop_iw_p1_poisoned;
      5'b10011:
        casez_tmp_228 = stq_19_bits_uop_iw_p1_poisoned;
      5'b10100:
        casez_tmp_228 = stq_20_bits_uop_iw_p1_poisoned;
      5'b10101:
        casez_tmp_228 = stq_21_bits_uop_iw_p1_poisoned;
      5'b10110:
        casez_tmp_228 = stq_22_bits_uop_iw_p1_poisoned;
      5'b10111:
        casez_tmp_228 = stq_23_bits_uop_iw_p1_poisoned;
      5'b11000:
        casez_tmp_228 = stq_24_bits_uop_iw_p1_poisoned;
      5'b11001:
        casez_tmp_228 = stq_25_bits_uop_iw_p1_poisoned;
      5'b11010:
        casez_tmp_228 = stq_26_bits_uop_iw_p1_poisoned;
      5'b11011:
        casez_tmp_228 = stq_27_bits_uop_iw_p1_poisoned;
      5'b11100:
        casez_tmp_228 = stq_28_bits_uop_iw_p1_poisoned;
      5'b11101:
        casez_tmp_228 = stq_29_bits_uop_iw_p1_poisoned;
      5'b11110:
        casez_tmp_228 = stq_30_bits_uop_iw_p1_poisoned;
      default:
        casez_tmp_228 = stq_31_bits_uop_iw_p1_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_229;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_229 = stq_0_bits_uop_iw_p2_poisoned;
      5'b00001:
        casez_tmp_229 = stq_1_bits_uop_iw_p2_poisoned;
      5'b00010:
        casez_tmp_229 = stq_2_bits_uop_iw_p2_poisoned;
      5'b00011:
        casez_tmp_229 = stq_3_bits_uop_iw_p2_poisoned;
      5'b00100:
        casez_tmp_229 = stq_4_bits_uop_iw_p2_poisoned;
      5'b00101:
        casez_tmp_229 = stq_5_bits_uop_iw_p2_poisoned;
      5'b00110:
        casez_tmp_229 = stq_6_bits_uop_iw_p2_poisoned;
      5'b00111:
        casez_tmp_229 = stq_7_bits_uop_iw_p2_poisoned;
      5'b01000:
        casez_tmp_229 = stq_8_bits_uop_iw_p2_poisoned;
      5'b01001:
        casez_tmp_229 = stq_9_bits_uop_iw_p2_poisoned;
      5'b01010:
        casez_tmp_229 = stq_10_bits_uop_iw_p2_poisoned;
      5'b01011:
        casez_tmp_229 = stq_11_bits_uop_iw_p2_poisoned;
      5'b01100:
        casez_tmp_229 = stq_12_bits_uop_iw_p2_poisoned;
      5'b01101:
        casez_tmp_229 = stq_13_bits_uop_iw_p2_poisoned;
      5'b01110:
        casez_tmp_229 = stq_14_bits_uop_iw_p2_poisoned;
      5'b01111:
        casez_tmp_229 = stq_15_bits_uop_iw_p2_poisoned;
      5'b10000:
        casez_tmp_229 = stq_16_bits_uop_iw_p2_poisoned;
      5'b10001:
        casez_tmp_229 = stq_17_bits_uop_iw_p2_poisoned;
      5'b10010:
        casez_tmp_229 = stq_18_bits_uop_iw_p2_poisoned;
      5'b10011:
        casez_tmp_229 = stq_19_bits_uop_iw_p2_poisoned;
      5'b10100:
        casez_tmp_229 = stq_20_bits_uop_iw_p2_poisoned;
      5'b10101:
        casez_tmp_229 = stq_21_bits_uop_iw_p2_poisoned;
      5'b10110:
        casez_tmp_229 = stq_22_bits_uop_iw_p2_poisoned;
      5'b10111:
        casez_tmp_229 = stq_23_bits_uop_iw_p2_poisoned;
      5'b11000:
        casez_tmp_229 = stq_24_bits_uop_iw_p2_poisoned;
      5'b11001:
        casez_tmp_229 = stq_25_bits_uop_iw_p2_poisoned;
      5'b11010:
        casez_tmp_229 = stq_26_bits_uop_iw_p2_poisoned;
      5'b11011:
        casez_tmp_229 = stq_27_bits_uop_iw_p2_poisoned;
      5'b11100:
        casez_tmp_229 = stq_28_bits_uop_iw_p2_poisoned;
      5'b11101:
        casez_tmp_229 = stq_29_bits_uop_iw_p2_poisoned;
      5'b11110:
        casez_tmp_229 = stq_30_bits_uop_iw_p2_poisoned;
      default:
        casez_tmp_229 = stq_31_bits_uop_iw_p2_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_230;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_230 = stq_0_bits_uop_is_br;
      5'b00001:
        casez_tmp_230 = stq_1_bits_uop_is_br;
      5'b00010:
        casez_tmp_230 = stq_2_bits_uop_is_br;
      5'b00011:
        casez_tmp_230 = stq_3_bits_uop_is_br;
      5'b00100:
        casez_tmp_230 = stq_4_bits_uop_is_br;
      5'b00101:
        casez_tmp_230 = stq_5_bits_uop_is_br;
      5'b00110:
        casez_tmp_230 = stq_6_bits_uop_is_br;
      5'b00111:
        casez_tmp_230 = stq_7_bits_uop_is_br;
      5'b01000:
        casez_tmp_230 = stq_8_bits_uop_is_br;
      5'b01001:
        casez_tmp_230 = stq_9_bits_uop_is_br;
      5'b01010:
        casez_tmp_230 = stq_10_bits_uop_is_br;
      5'b01011:
        casez_tmp_230 = stq_11_bits_uop_is_br;
      5'b01100:
        casez_tmp_230 = stq_12_bits_uop_is_br;
      5'b01101:
        casez_tmp_230 = stq_13_bits_uop_is_br;
      5'b01110:
        casez_tmp_230 = stq_14_bits_uop_is_br;
      5'b01111:
        casez_tmp_230 = stq_15_bits_uop_is_br;
      5'b10000:
        casez_tmp_230 = stq_16_bits_uop_is_br;
      5'b10001:
        casez_tmp_230 = stq_17_bits_uop_is_br;
      5'b10010:
        casez_tmp_230 = stq_18_bits_uop_is_br;
      5'b10011:
        casez_tmp_230 = stq_19_bits_uop_is_br;
      5'b10100:
        casez_tmp_230 = stq_20_bits_uop_is_br;
      5'b10101:
        casez_tmp_230 = stq_21_bits_uop_is_br;
      5'b10110:
        casez_tmp_230 = stq_22_bits_uop_is_br;
      5'b10111:
        casez_tmp_230 = stq_23_bits_uop_is_br;
      5'b11000:
        casez_tmp_230 = stq_24_bits_uop_is_br;
      5'b11001:
        casez_tmp_230 = stq_25_bits_uop_is_br;
      5'b11010:
        casez_tmp_230 = stq_26_bits_uop_is_br;
      5'b11011:
        casez_tmp_230 = stq_27_bits_uop_is_br;
      5'b11100:
        casez_tmp_230 = stq_28_bits_uop_is_br;
      5'b11101:
        casez_tmp_230 = stq_29_bits_uop_is_br;
      5'b11110:
        casez_tmp_230 = stq_30_bits_uop_is_br;
      default:
        casez_tmp_230 = stq_31_bits_uop_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_231;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_231 = stq_0_bits_uop_is_jalr;
      5'b00001:
        casez_tmp_231 = stq_1_bits_uop_is_jalr;
      5'b00010:
        casez_tmp_231 = stq_2_bits_uop_is_jalr;
      5'b00011:
        casez_tmp_231 = stq_3_bits_uop_is_jalr;
      5'b00100:
        casez_tmp_231 = stq_4_bits_uop_is_jalr;
      5'b00101:
        casez_tmp_231 = stq_5_bits_uop_is_jalr;
      5'b00110:
        casez_tmp_231 = stq_6_bits_uop_is_jalr;
      5'b00111:
        casez_tmp_231 = stq_7_bits_uop_is_jalr;
      5'b01000:
        casez_tmp_231 = stq_8_bits_uop_is_jalr;
      5'b01001:
        casez_tmp_231 = stq_9_bits_uop_is_jalr;
      5'b01010:
        casez_tmp_231 = stq_10_bits_uop_is_jalr;
      5'b01011:
        casez_tmp_231 = stq_11_bits_uop_is_jalr;
      5'b01100:
        casez_tmp_231 = stq_12_bits_uop_is_jalr;
      5'b01101:
        casez_tmp_231 = stq_13_bits_uop_is_jalr;
      5'b01110:
        casez_tmp_231 = stq_14_bits_uop_is_jalr;
      5'b01111:
        casez_tmp_231 = stq_15_bits_uop_is_jalr;
      5'b10000:
        casez_tmp_231 = stq_16_bits_uop_is_jalr;
      5'b10001:
        casez_tmp_231 = stq_17_bits_uop_is_jalr;
      5'b10010:
        casez_tmp_231 = stq_18_bits_uop_is_jalr;
      5'b10011:
        casez_tmp_231 = stq_19_bits_uop_is_jalr;
      5'b10100:
        casez_tmp_231 = stq_20_bits_uop_is_jalr;
      5'b10101:
        casez_tmp_231 = stq_21_bits_uop_is_jalr;
      5'b10110:
        casez_tmp_231 = stq_22_bits_uop_is_jalr;
      5'b10111:
        casez_tmp_231 = stq_23_bits_uop_is_jalr;
      5'b11000:
        casez_tmp_231 = stq_24_bits_uop_is_jalr;
      5'b11001:
        casez_tmp_231 = stq_25_bits_uop_is_jalr;
      5'b11010:
        casez_tmp_231 = stq_26_bits_uop_is_jalr;
      5'b11011:
        casez_tmp_231 = stq_27_bits_uop_is_jalr;
      5'b11100:
        casez_tmp_231 = stq_28_bits_uop_is_jalr;
      5'b11101:
        casez_tmp_231 = stq_29_bits_uop_is_jalr;
      5'b11110:
        casez_tmp_231 = stq_30_bits_uop_is_jalr;
      default:
        casez_tmp_231 = stq_31_bits_uop_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_232;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_232 = stq_0_bits_uop_is_jal;
      5'b00001:
        casez_tmp_232 = stq_1_bits_uop_is_jal;
      5'b00010:
        casez_tmp_232 = stq_2_bits_uop_is_jal;
      5'b00011:
        casez_tmp_232 = stq_3_bits_uop_is_jal;
      5'b00100:
        casez_tmp_232 = stq_4_bits_uop_is_jal;
      5'b00101:
        casez_tmp_232 = stq_5_bits_uop_is_jal;
      5'b00110:
        casez_tmp_232 = stq_6_bits_uop_is_jal;
      5'b00111:
        casez_tmp_232 = stq_7_bits_uop_is_jal;
      5'b01000:
        casez_tmp_232 = stq_8_bits_uop_is_jal;
      5'b01001:
        casez_tmp_232 = stq_9_bits_uop_is_jal;
      5'b01010:
        casez_tmp_232 = stq_10_bits_uop_is_jal;
      5'b01011:
        casez_tmp_232 = stq_11_bits_uop_is_jal;
      5'b01100:
        casez_tmp_232 = stq_12_bits_uop_is_jal;
      5'b01101:
        casez_tmp_232 = stq_13_bits_uop_is_jal;
      5'b01110:
        casez_tmp_232 = stq_14_bits_uop_is_jal;
      5'b01111:
        casez_tmp_232 = stq_15_bits_uop_is_jal;
      5'b10000:
        casez_tmp_232 = stq_16_bits_uop_is_jal;
      5'b10001:
        casez_tmp_232 = stq_17_bits_uop_is_jal;
      5'b10010:
        casez_tmp_232 = stq_18_bits_uop_is_jal;
      5'b10011:
        casez_tmp_232 = stq_19_bits_uop_is_jal;
      5'b10100:
        casez_tmp_232 = stq_20_bits_uop_is_jal;
      5'b10101:
        casez_tmp_232 = stq_21_bits_uop_is_jal;
      5'b10110:
        casez_tmp_232 = stq_22_bits_uop_is_jal;
      5'b10111:
        casez_tmp_232 = stq_23_bits_uop_is_jal;
      5'b11000:
        casez_tmp_232 = stq_24_bits_uop_is_jal;
      5'b11001:
        casez_tmp_232 = stq_25_bits_uop_is_jal;
      5'b11010:
        casez_tmp_232 = stq_26_bits_uop_is_jal;
      5'b11011:
        casez_tmp_232 = stq_27_bits_uop_is_jal;
      5'b11100:
        casez_tmp_232 = stq_28_bits_uop_is_jal;
      5'b11101:
        casez_tmp_232 = stq_29_bits_uop_is_jal;
      5'b11110:
        casez_tmp_232 = stq_30_bits_uop_is_jal;
      default:
        casez_tmp_232 = stq_31_bits_uop_is_jal;
    endcase
  end // always @(*)
  reg         casez_tmp_233;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_233 = stq_0_bits_uop_is_sfb;
      5'b00001:
        casez_tmp_233 = stq_1_bits_uop_is_sfb;
      5'b00010:
        casez_tmp_233 = stq_2_bits_uop_is_sfb;
      5'b00011:
        casez_tmp_233 = stq_3_bits_uop_is_sfb;
      5'b00100:
        casez_tmp_233 = stq_4_bits_uop_is_sfb;
      5'b00101:
        casez_tmp_233 = stq_5_bits_uop_is_sfb;
      5'b00110:
        casez_tmp_233 = stq_6_bits_uop_is_sfb;
      5'b00111:
        casez_tmp_233 = stq_7_bits_uop_is_sfb;
      5'b01000:
        casez_tmp_233 = stq_8_bits_uop_is_sfb;
      5'b01001:
        casez_tmp_233 = stq_9_bits_uop_is_sfb;
      5'b01010:
        casez_tmp_233 = stq_10_bits_uop_is_sfb;
      5'b01011:
        casez_tmp_233 = stq_11_bits_uop_is_sfb;
      5'b01100:
        casez_tmp_233 = stq_12_bits_uop_is_sfb;
      5'b01101:
        casez_tmp_233 = stq_13_bits_uop_is_sfb;
      5'b01110:
        casez_tmp_233 = stq_14_bits_uop_is_sfb;
      5'b01111:
        casez_tmp_233 = stq_15_bits_uop_is_sfb;
      5'b10000:
        casez_tmp_233 = stq_16_bits_uop_is_sfb;
      5'b10001:
        casez_tmp_233 = stq_17_bits_uop_is_sfb;
      5'b10010:
        casez_tmp_233 = stq_18_bits_uop_is_sfb;
      5'b10011:
        casez_tmp_233 = stq_19_bits_uop_is_sfb;
      5'b10100:
        casez_tmp_233 = stq_20_bits_uop_is_sfb;
      5'b10101:
        casez_tmp_233 = stq_21_bits_uop_is_sfb;
      5'b10110:
        casez_tmp_233 = stq_22_bits_uop_is_sfb;
      5'b10111:
        casez_tmp_233 = stq_23_bits_uop_is_sfb;
      5'b11000:
        casez_tmp_233 = stq_24_bits_uop_is_sfb;
      5'b11001:
        casez_tmp_233 = stq_25_bits_uop_is_sfb;
      5'b11010:
        casez_tmp_233 = stq_26_bits_uop_is_sfb;
      5'b11011:
        casez_tmp_233 = stq_27_bits_uop_is_sfb;
      5'b11100:
        casez_tmp_233 = stq_28_bits_uop_is_sfb;
      5'b11101:
        casez_tmp_233 = stq_29_bits_uop_is_sfb;
      5'b11110:
        casez_tmp_233 = stq_30_bits_uop_is_sfb;
      default:
        casez_tmp_233 = stq_31_bits_uop_is_sfb;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_234;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_234 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_234 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_234 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_234 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_234 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_234 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_234 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_234 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_234 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_234 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_234 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_234 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_234 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_234 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_234 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_234 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_234 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_234 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_234 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_234 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_234 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_234 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_234 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_234 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_234 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_234 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_234 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_234 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_234 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_234 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_234 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_234 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_235;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_235 = stq_0_bits_uop_br_tag;
      5'b00001:
        casez_tmp_235 = stq_1_bits_uop_br_tag;
      5'b00010:
        casez_tmp_235 = stq_2_bits_uop_br_tag;
      5'b00011:
        casez_tmp_235 = stq_3_bits_uop_br_tag;
      5'b00100:
        casez_tmp_235 = stq_4_bits_uop_br_tag;
      5'b00101:
        casez_tmp_235 = stq_5_bits_uop_br_tag;
      5'b00110:
        casez_tmp_235 = stq_6_bits_uop_br_tag;
      5'b00111:
        casez_tmp_235 = stq_7_bits_uop_br_tag;
      5'b01000:
        casez_tmp_235 = stq_8_bits_uop_br_tag;
      5'b01001:
        casez_tmp_235 = stq_9_bits_uop_br_tag;
      5'b01010:
        casez_tmp_235 = stq_10_bits_uop_br_tag;
      5'b01011:
        casez_tmp_235 = stq_11_bits_uop_br_tag;
      5'b01100:
        casez_tmp_235 = stq_12_bits_uop_br_tag;
      5'b01101:
        casez_tmp_235 = stq_13_bits_uop_br_tag;
      5'b01110:
        casez_tmp_235 = stq_14_bits_uop_br_tag;
      5'b01111:
        casez_tmp_235 = stq_15_bits_uop_br_tag;
      5'b10000:
        casez_tmp_235 = stq_16_bits_uop_br_tag;
      5'b10001:
        casez_tmp_235 = stq_17_bits_uop_br_tag;
      5'b10010:
        casez_tmp_235 = stq_18_bits_uop_br_tag;
      5'b10011:
        casez_tmp_235 = stq_19_bits_uop_br_tag;
      5'b10100:
        casez_tmp_235 = stq_20_bits_uop_br_tag;
      5'b10101:
        casez_tmp_235 = stq_21_bits_uop_br_tag;
      5'b10110:
        casez_tmp_235 = stq_22_bits_uop_br_tag;
      5'b10111:
        casez_tmp_235 = stq_23_bits_uop_br_tag;
      5'b11000:
        casez_tmp_235 = stq_24_bits_uop_br_tag;
      5'b11001:
        casez_tmp_235 = stq_25_bits_uop_br_tag;
      5'b11010:
        casez_tmp_235 = stq_26_bits_uop_br_tag;
      5'b11011:
        casez_tmp_235 = stq_27_bits_uop_br_tag;
      5'b11100:
        casez_tmp_235 = stq_28_bits_uop_br_tag;
      5'b11101:
        casez_tmp_235 = stq_29_bits_uop_br_tag;
      5'b11110:
        casez_tmp_235 = stq_30_bits_uop_br_tag;
      default:
        casez_tmp_235 = stq_31_bits_uop_br_tag;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_236;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_236 = stq_0_bits_uop_ftq_idx;
      5'b00001:
        casez_tmp_236 = stq_1_bits_uop_ftq_idx;
      5'b00010:
        casez_tmp_236 = stq_2_bits_uop_ftq_idx;
      5'b00011:
        casez_tmp_236 = stq_3_bits_uop_ftq_idx;
      5'b00100:
        casez_tmp_236 = stq_4_bits_uop_ftq_idx;
      5'b00101:
        casez_tmp_236 = stq_5_bits_uop_ftq_idx;
      5'b00110:
        casez_tmp_236 = stq_6_bits_uop_ftq_idx;
      5'b00111:
        casez_tmp_236 = stq_7_bits_uop_ftq_idx;
      5'b01000:
        casez_tmp_236 = stq_8_bits_uop_ftq_idx;
      5'b01001:
        casez_tmp_236 = stq_9_bits_uop_ftq_idx;
      5'b01010:
        casez_tmp_236 = stq_10_bits_uop_ftq_idx;
      5'b01011:
        casez_tmp_236 = stq_11_bits_uop_ftq_idx;
      5'b01100:
        casez_tmp_236 = stq_12_bits_uop_ftq_idx;
      5'b01101:
        casez_tmp_236 = stq_13_bits_uop_ftq_idx;
      5'b01110:
        casez_tmp_236 = stq_14_bits_uop_ftq_idx;
      5'b01111:
        casez_tmp_236 = stq_15_bits_uop_ftq_idx;
      5'b10000:
        casez_tmp_236 = stq_16_bits_uop_ftq_idx;
      5'b10001:
        casez_tmp_236 = stq_17_bits_uop_ftq_idx;
      5'b10010:
        casez_tmp_236 = stq_18_bits_uop_ftq_idx;
      5'b10011:
        casez_tmp_236 = stq_19_bits_uop_ftq_idx;
      5'b10100:
        casez_tmp_236 = stq_20_bits_uop_ftq_idx;
      5'b10101:
        casez_tmp_236 = stq_21_bits_uop_ftq_idx;
      5'b10110:
        casez_tmp_236 = stq_22_bits_uop_ftq_idx;
      5'b10111:
        casez_tmp_236 = stq_23_bits_uop_ftq_idx;
      5'b11000:
        casez_tmp_236 = stq_24_bits_uop_ftq_idx;
      5'b11001:
        casez_tmp_236 = stq_25_bits_uop_ftq_idx;
      5'b11010:
        casez_tmp_236 = stq_26_bits_uop_ftq_idx;
      5'b11011:
        casez_tmp_236 = stq_27_bits_uop_ftq_idx;
      5'b11100:
        casez_tmp_236 = stq_28_bits_uop_ftq_idx;
      5'b11101:
        casez_tmp_236 = stq_29_bits_uop_ftq_idx;
      5'b11110:
        casez_tmp_236 = stq_30_bits_uop_ftq_idx;
      default:
        casez_tmp_236 = stq_31_bits_uop_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_237;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_237 = stq_0_bits_uop_edge_inst;
      5'b00001:
        casez_tmp_237 = stq_1_bits_uop_edge_inst;
      5'b00010:
        casez_tmp_237 = stq_2_bits_uop_edge_inst;
      5'b00011:
        casez_tmp_237 = stq_3_bits_uop_edge_inst;
      5'b00100:
        casez_tmp_237 = stq_4_bits_uop_edge_inst;
      5'b00101:
        casez_tmp_237 = stq_5_bits_uop_edge_inst;
      5'b00110:
        casez_tmp_237 = stq_6_bits_uop_edge_inst;
      5'b00111:
        casez_tmp_237 = stq_7_bits_uop_edge_inst;
      5'b01000:
        casez_tmp_237 = stq_8_bits_uop_edge_inst;
      5'b01001:
        casez_tmp_237 = stq_9_bits_uop_edge_inst;
      5'b01010:
        casez_tmp_237 = stq_10_bits_uop_edge_inst;
      5'b01011:
        casez_tmp_237 = stq_11_bits_uop_edge_inst;
      5'b01100:
        casez_tmp_237 = stq_12_bits_uop_edge_inst;
      5'b01101:
        casez_tmp_237 = stq_13_bits_uop_edge_inst;
      5'b01110:
        casez_tmp_237 = stq_14_bits_uop_edge_inst;
      5'b01111:
        casez_tmp_237 = stq_15_bits_uop_edge_inst;
      5'b10000:
        casez_tmp_237 = stq_16_bits_uop_edge_inst;
      5'b10001:
        casez_tmp_237 = stq_17_bits_uop_edge_inst;
      5'b10010:
        casez_tmp_237 = stq_18_bits_uop_edge_inst;
      5'b10011:
        casez_tmp_237 = stq_19_bits_uop_edge_inst;
      5'b10100:
        casez_tmp_237 = stq_20_bits_uop_edge_inst;
      5'b10101:
        casez_tmp_237 = stq_21_bits_uop_edge_inst;
      5'b10110:
        casez_tmp_237 = stq_22_bits_uop_edge_inst;
      5'b10111:
        casez_tmp_237 = stq_23_bits_uop_edge_inst;
      5'b11000:
        casez_tmp_237 = stq_24_bits_uop_edge_inst;
      5'b11001:
        casez_tmp_237 = stq_25_bits_uop_edge_inst;
      5'b11010:
        casez_tmp_237 = stq_26_bits_uop_edge_inst;
      5'b11011:
        casez_tmp_237 = stq_27_bits_uop_edge_inst;
      5'b11100:
        casez_tmp_237 = stq_28_bits_uop_edge_inst;
      5'b11101:
        casez_tmp_237 = stq_29_bits_uop_edge_inst;
      5'b11110:
        casez_tmp_237 = stq_30_bits_uop_edge_inst;
      default:
        casez_tmp_237 = stq_31_bits_uop_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_238;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_238 = stq_0_bits_uop_pc_lob;
      5'b00001:
        casez_tmp_238 = stq_1_bits_uop_pc_lob;
      5'b00010:
        casez_tmp_238 = stq_2_bits_uop_pc_lob;
      5'b00011:
        casez_tmp_238 = stq_3_bits_uop_pc_lob;
      5'b00100:
        casez_tmp_238 = stq_4_bits_uop_pc_lob;
      5'b00101:
        casez_tmp_238 = stq_5_bits_uop_pc_lob;
      5'b00110:
        casez_tmp_238 = stq_6_bits_uop_pc_lob;
      5'b00111:
        casez_tmp_238 = stq_7_bits_uop_pc_lob;
      5'b01000:
        casez_tmp_238 = stq_8_bits_uop_pc_lob;
      5'b01001:
        casez_tmp_238 = stq_9_bits_uop_pc_lob;
      5'b01010:
        casez_tmp_238 = stq_10_bits_uop_pc_lob;
      5'b01011:
        casez_tmp_238 = stq_11_bits_uop_pc_lob;
      5'b01100:
        casez_tmp_238 = stq_12_bits_uop_pc_lob;
      5'b01101:
        casez_tmp_238 = stq_13_bits_uop_pc_lob;
      5'b01110:
        casez_tmp_238 = stq_14_bits_uop_pc_lob;
      5'b01111:
        casez_tmp_238 = stq_15_bits_uop_pc_lob;
      5'b10000:
        casez_tmp_238 = stq_16_bits_uop_pc_lob;
      5'b10001:
        casez_tmp_238 = stq_17_bits_uop_pc_lob;
      5'b10010:
        casez_tmp_238 = stq_18_bits_uop_pc_lob;
      5'b10011:
        casez_tmp_238 = stq_19_bits_uop_pc_lob;
      5'b10100:
        casez_tmp_238 = stq_20_bits_uop_pc_lob;
      5'b10101:
        casez_tmp_238 = stq_21_bits_uop_pc_lob;
      5'b10110:
        casez_tmp_238 = stq_22_bits_uop_pc_lob;
      5'b10111:
        casez_tmp_238 = stq_23_bits_uop_pc_lob;
      5'b11000:
        casez_tmp_238 = stq_24_bits_uop_pc_lob;
      5'b11001:
        casez_tmp_238 = stq_25_bits_uop_pc_lob;
      5'b11010:
        casez_tmp_238 = stq_26_bits_uop_pc_lob;
      5'b11011:
        casez_tmp_238 = stq_27_bits_uop_pc_lob;
      5'b11100:
        casez_tmp_238 = stq_28_bits_uop_pc_lob;
      5'b11101:
        casez_tmp_238 = stq_29_bits_uop_pc_lob;
      5'b11110:
        casez_tmp_238 = stq_30_bits_uop_pc_lob;
      default:
        casez_tmp_238 = stq_31_bits_uop_pc_lob;
    endcase
  end // always @(*)
  reg         casez_tmp_239;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_239 = stq_0_bits_uop_taken;
      5'b00001:
        casez_tmp_239 = stq_1_bits_uop_taken;
      5'b00010:
        casez_tmp_239 = stq_2_bits_uop_taken;
      5'b00011:
        casez_tmp_239 = stq_3_bits_uop_taken;
      5'b00100:
        casez_tmp_239 = stq_4_bits_uop_taken;
      5'b00101:
        casez_tmp_239 = stq_5_bits_uop_taken;
      5'b00110:
        casez_tmp_239 = stq_6_bits_uop_taken;
      5'b00111:
        casez_tmp_239 = stq_7_bits_uop_taken;
      5'b01000:
        casez_tmp_239 = stq_8_bits_uop_taken;
      5'b01001:
        casez_tmp_239 = stq_9_bits_uop_taken;
      5'b01010:
        casez_tmp_239 = stq_10_bits_uop_taken;
      5'b01011:
        casez_tmp_239 = stq_11_bits_uop_taken;
      5'b01100:
        casez_tmp_239 = stq_12_bits_uop_taken;
      5'b01101:
        casez_tmp_239 = stq_13_bits_uop_taken;
      5'b01110:
        casez_tmp_239 = stq_14_bits_uop_taken;
      5'b01111:
        casez_tmp_239 = stq_15_bits_uop_taken;
      5'b10000:
        casez_tmp_239 = stq_16_bits_uop_taken;
      5'b10001:
        casez_tmp_239 = stq_17_bits_uop_taken;
      5'b10010:
        casez_tmp_239 = stq_18_bits_uop_taken;
      5'b10011:
        casez_tmp_239 = stq_19_bits_uop_taken;
      5'b10100:
        casez_tmp_239 = stq_20_bits_uop_taken;
      5'b10101:
        casez_tmp_239 = stq_21_bits_uop_taken;
      5'b10110:
        casez_tmp_239 = stq_22_bits_uop_taken;
      5'b10111:
        casez_tmp_239 = stq_23_bits_uop_taken;
      5'b11000:
        casez_tmp_239 = stq_24_bits_uop_taken;
      5'b11001:
        casez_tmp_239 = stq_25_bits_uop_taken;
      5'b11010:
        casez_tmp_239 = stq_26_bits_uop_taken;
      5'b11011:
        casez_tmp_239 = stq_27_bits_uop_taken;
      5'b11100:
        casez_tmp_239 = stq_28_bits_uop_taken;
      5'b11101:
        casez_tmp_239 = stq_29_bits_uop_taken;
      5'b11110:
        casez_tmp_239 = stq_30_bits_uop_taken;
      default:
        casez_tmp_239 = stq_31_bits_uop_taken;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_240;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_240 = stq_0_bits_uop_imm_packed;
      5'b00001:
        casez_tmp_240 = stq_1_bits_uop_imm_packed;
      5'b00010:
        casez_tmp_240 = stq_2_bits_uop_imm_packed;
      5'b00011:
        casez_tmp_240 = stq_3_bits_uop_imm_packed;
      5'b00100:
        casez_tmp_240 = stq_4_bits_uop_imm_packed;
      5'b00101:
        casez_tmp_240 = stq_5_bits_uop_imm_packed;
      5'b00110:
        casez_tmp_240 = stq_6_bits_uop_imm_packed;
      5'b00111:
        casez_tmp_240 = stq_7_bits_uop_imm_packed;
      5'b01000:
        casez_tmp_240 = stq_8_bits_uop_imm_packed;
      5'b01001:
        casez_tmp_240 = stq_9_bits_uop_imm_packed;
      5'b01010:
        casez_tmp_240 = stq_10_bits_uop_imm_packed;
      5'b01011:
        casez_tmp_240 = stq_11_bits_uop_imm_packed;
      5'b01100:
        casez_tmp_240 = stq_12_bits_uop_imm_packed;
      5'b01101:
        casez_tmp_240 = stq_13_bits_uop_imm_packed;
      5'b01110:
        casez_tmp_240 = stq_14_bits_uop_imm_packed;
      5'b01111:
        casez_tmp_240 = stq_15_bits_uop_imm_packed;
      5'b10000:
        casez_tmp_240 = stq_16_bits_uop_imm_packed;
      5'b10001:
        casez_tmp_240 = stq_17_bits_uop_imm_packed;
      5'b10010:
        casez_tmp_240 = stq_18_bits_uop_imm_packed;
      5'b10011:
        casez_tmp_240 = stq_19_bits_uop_imm_packed;
      5'b10100:
        casez_tmp_240 = stq_20_bits_uop_imm_packed;
      5'b10101:
        casez_tmp_240 = stq_21_bits_uop_imm_packed;
      5'b10110:
        casez_tmp_240 = stq_22_bits_uop_imm_packed;
      5'b10111:
        casez_tmp_240 = stq_23_bits_uop_imm_packed;
      5'b11000:
        casez_tmp_240 = stq_24_bits_uop_imm_packed;
      5'b11001:
        casez_tmp_240 = stq_25_bits_uop_imm_packed;
      5'b11010:
        casez_tmp_240 = stq_26_bits_uop_imm_packed;
      5'b11011:
        casez_tmp_240 = stq_27_bits_uop_imm_packed;
      5'b11100:
        casez_tmp_240 = stq_28_bits_uop_imm_packed;
      5'b11101:
        casez_tmp_240 = stq_29_bits_uop_imm_packed;
      5'b11110:
        casez_tmp_240 = stq_30_bits_uop_imm_packed;
      default:
        casez_tmp_240 = stq_31_bits_uop_imm_packed;
    endcase
  end // always @(*)
  reg  [11:0] casez_tmp_241;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_241 = stq_0_bits_uop_csr_addr;
      5'b00001:
        casez_tmp_241 = stq_1_bits_uop_csr_addr;
      5'b00010:
        casez_tmp_241 = stq_2_bits_uop_csr_addr;
      5'b00011:
        casez_tmp_241 = stq_3_bits_uop_csr_addr;
      5'b00100:
        casez_tmp_241 = stq_4_bits_uop_csr_addr;
      5'b00101:
        casez_tmp_241 = stq_5_bits_uop_csr_addr;
      5'b00110:
        casez_tmp_241 = stq_6_bits_uop_csr_addr;
      5'b00111:
        casez_tmp_241 = stq_7_bits_uop_csr_addr;
      5'b01000:
        casez_tmp_241 = stq_8_bits_uop_csr_addr;
      5'b01001:
        casez_tmp_241 = stq_9_bits_uop_csr_addr;
      5'b01010:
        casez_tmp_241 = stq_10_bits_uop_csr_addr;
      5'b01011:
        casez_tmp_241 = stq_11_bits_uop_csr_addr;
      5'b01100:
        casez_tmp_241 = stq_12_bits_uop_csr_addr;
      5'b01101:
        casez_tmp_241 = stq_13_bits_uop_csr_addr;
      5'b01110:
        casez_tmp_241 = stq_14_bits_uop_csr_addr;
      5'b01111:
        casez_tmp_241 = stq_15_bits_uop_csr_addr;
      5'b10000:
        casez_tmp_241 = stq_16_bits_uop_csr_addr;
      5'b10001:
        casez_tmp_241 = stq_17_bits_uop_csr_addr;
      5'b10010:
        casez_tmp_241 = stq_18_bits_uop_csr_addr;
      5'b10011:
        casez_tmp_241 = stq_19_bits_uop_csr_addr;
      5'b10100:
        casez_tmp_241 = stq_20_bits_uop_csr_addr;
      5'b10101:
        casez_tmp_241 = stq_21_bits_uop_csr_addr;
      5'b10110:
        casez_tmp_241 = stq_22_bits_uop_csr_addr;
      5'b10111:
        casez_tmp_241 = stq_23_bits_uop_csr_addr;
      5'b11000:
        casez_tmp_241 = stq_24_bits_uop_csr_addr;
      5'b11001:
        casez_tmp_241 = stq_25_bits_uop_csr_addr;
      5'b11010:
        casez_tmp_241 = stq_26_bits_uop_csr_addr;
      5'b11011:
        casez_tmp_241 = stq_27_bits_uop_csr_addr;
      5'b11100:
        casez_tmp_241 = stq_28_bits_uop_csr_addr;
      5'b11101:
        casez_tmp_241 = stq_29_bits_uop_csr_addr;
      5'b11110:
        casez_tmp_241 = stq_30_bits_uop_csr_addr;
      default:
        casez_tmp_241 = stq_31_bits_uop_csr_addr;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_242;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_242 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_242 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_242 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_242 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_242 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_242 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_242 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_242 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_242 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_242 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_242 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_242 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_242 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_242 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_242 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_242 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_242 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_242 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_242 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_242 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_242 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_242 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_242 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_242 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_242 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_242 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_242 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_242 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_242 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_242 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_242 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_242 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_243;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_243 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_243 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_243 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_243 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_243 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_243 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_243 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_243 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_243 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_243 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_243 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_243 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_243 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_243 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_243 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_243 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_243 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_243 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_243 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_243 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_243 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_243 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_243 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_243 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_243 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_243 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_243 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_243 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_243 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_243 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_243 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_243 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_244;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_244 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_244 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_244 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_244 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_244 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_244 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_244 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_244 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_244 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_244 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_244 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_244 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_244 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_244 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_244 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_244 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_244 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_244 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_244 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_244 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_244 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_244 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_244 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_244 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_244 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_244 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_244 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_244 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_244 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_244 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_244 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_244 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_245;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_245 = stq_0_bits_uop_rxq_idx;
      5'b00001:
        casez_tmp_245 = stq_1_bits_uop_rxq_idx;
      5'b00010:
        casez_tmp_245 = stq_2_bits_uop_rxq_idx;
      5'b00011:
        casez_tmp_245 = stq_3_bits_uop_rxq_idx;
      5'b00100:
        casez_tmp_245 = stq_4_bits_uop_rxq_idx;
      5'b00101:
        casez_tmp_245 = stq_5_bits_uop_rxq_idx;
      5'b00110:
        casez_tmp_245 = stq_6_bits_uop_rxq_idx;
      5'b00111:
        casez_tmp_245 = stq_7_bits_uop_rxq_idx;
      5'b01000:
        casez_tmp_245 = stq_8_bits_uop_rxq_idx;
      5'b01001:
        casez_tmp_245 = stq_9_bits_uop_rxq_idx;
      5'b01010:
        casez_tmp_245 = stq_10_bits_uop_rxq_idx;
      5'b01011:
        casez_tmp_245 = stq_11_bits_uop_rxq_idx;
      5'b01100:
        casez_tmp_245 = stq_12_bits_uop_rxq_idx;
      5'b01101:
        casez_tmp_245 = stq_13_bits_uop_rxq_idx;
      5'b01110:
        casez_tmp_245 = stq_14_bits_uop_rxq_idx;
      5'b01111:
        casez_tmp_245 = stq_15_bits_uop_rxq_idx;
      5'b10000:
        casez_tmp_245 = stq_16_bits_uop_rxq_idx;
      5'b10001:
        casez_tmp_245 = stq_17_bits_uop_rxq_idx;
      5'b10010:
        casez_tmp_245 = stq_18_bits_uop_rxq_idx;
      5'b10011:
        casez_tmp_245 = stq_19_bits_uop_rxq_idx;
      5'b10100:
        casez_tmp_245 = stq_20_bits_uop_rxq_idx;
      5'b10101:
        casez_tmp_245 = stq_21_bits_uop_rxq_idx;
      5'b10110:
        casez_tmp_245 = stq_22_bits_uop_rxq_idx;
      5'b10111:
        casez_tmp_245 = stq_23_bits_uop_rxq_idx;
      5'b11000:
        casez_tmp_245 = stq_24_bits_uop_rxq_idx;
      5'b11001:
        casez_tmp_245 = stq_25_bits_uop_rxq_idx;
      5'b11010:
        casez_tmp_245 = stq_26_bits_uop_rxq_idx;
      5'b11011:
        casez_tmp_245 = stq_27_bits_uop_rxq_idx;
      5'b11100:
        casez_tmp_245 = stq_28_bits_uop_rxq_idx;
      5'b11101:
        casez_tmp_245 = stq_29_bits_uop_rxq_idx;
      5'b11110:
        casez_tmp_245 = stq_30_bits_uop_rxq_idx;
      default:
        casez_tmp_245 = stq_31_bits_uop_rxq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_246;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_246 = stq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_246 = stq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_246 = stq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_246 = stq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_246 = stq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_246 = stq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_246 = stq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_246 = stq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_246 = stq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_246 = stq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_246 = stq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_246 = stq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_246 = stq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_246 = stq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_246 = stq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_246 = stq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_246 = stq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_246 = stq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_246 = stq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_246 = stq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_246 = stq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_246 = stq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_246 = stq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_246 = stq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_246 = stq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_246 = stq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_246 = stq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_246 = stq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_246 = stq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_246 = stq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_246 = stq_30_bits_uop_pdst;
      default:
        casez_tmp_246 = stq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_247;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_247 = stq_0_bits_uop_prs1;
      5'b00001:
        casez_tmp_247 = stq_1_bits_uop_prs1;
      5'b00010:
        casez_tmp_247 = stq_2_bits_uop_prs1;
      5'b00011:
        casez_tmp_247 = stq_3_bits_uop_prs1;
      5'b00100:
        casez_tmp_247 = stq_4_bits_uop_prs1;
      5'b00101:
        casez_tmp_247 = stq_5_bits_uop_prs1;
      5'b00110:
        casez_tmp_247 = stq_6_bits_uop_prs1;
      5'b00111:
        casez_tmp_247 = stq_7_bits_uop_prs1;
      5'b01000:
        casez_tmp_247 = stq_8_bits_uop_prs1;
      5'b01001:
        casez_tmp_247 = stq_9_bits_uop_prs1;
      5'b01010:
        casez_tmp_247 = stq_10_bits_uop_prs1;
      5'b01011:
        casez_tmp_247 = stq_11_bits_uop_prs1;
      5'b01100:
        casez_tmp_247 = stq_12_bits_uop_prs1;
      5'b01101:
        casez_tmp_247 = stq_13_bits_uop_prs1;
      5'b01110:
        casez_tmp_247 = stq_14_bits_uop_prs1;
      5'b01111:
        casez_tmp_247 = stq_15_bits_uop_prs1;
      5'b10000:
        casez_tmp_247 = stq_16_bits_uop_prs1;
      5'b10001:
        casez_tmp_247 = stq_17_bits_uop_prs1;
      5'b10010:
        casez_tmp_247 = stq_18_bits_uop_prs1;
      5'b10011:
        casez_tmp_247 = stq_19_bits_uop_prs1;
      5'b10100:
        casez_tmp_247 = stq_20_bits_uop_prs1;
      5'b10101:
        casez_tmp_247 = stq_21_bits_uop_prs1;
      5'b10110:
        casez_tmp_247 = stq_22_bits_uop_prs1;
      5'b10111:
        casez_tmp_247 = stq_23_bits_uop_prs1;
      5'b11000:
        casez_tmp_247 = stq_24_bits_uop_prs1;
      5'b11001:
        casez_tmp_247 = stq_25_bits_uop_prs1;
      5'b11010:
        casez_tmp_247 = stq_26_bits_uop_prs1;
      5'b11011:
        casez_tmp_247 = stq_27_bits_uop_prs1;
      5'b11100:
        casez_tmp_247 = stq_28_bits_uop_prs1;
      5'b11101:
        casez_tmp_247 = stq_29_bits_uop_prs1;
      5'b11110:
        casez_tmp_247 = stq_30_bits_uop_prs1;
      default:
        casez_tmp_247 = stq_31_bits_uop_prs1;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_248;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_248 = stq_0_bits_uop_prs2;
      5'b00001:
        casez_tmp_248 = stq_1_bits_uop_prs2;
      5'b00010:
        casez_tmp_248 = stq_2_bits_uop_prs2;
      5'b00011:
        casez_tmp_248 = stq_3_bits_uop_prs2;
      5'b00100:
        casez_tmp_248 = stq_4_bits_uop_prs2;
      5'b00101:
        casez_tmp_248 = stq_5_bits_uop_prs2;
      5'b00110:
        casez_tmp_248 = stq_6_bits_uop_prs2;
      5'b00111:
        casez_tmp_248 = stq_7_bits_uop_prs2;
      5'b01000:
        casez_tmp_248 = stq_8_bits_uop_prs2;
      5'b01001:
        casez_tmp_248 = stq_9_bits_uop_prs2;
      5'b01010:
        casez_tmp_248 = stq_10_bits_uop_prs2;
      5'b01011:
        casez_tmp_248 = stq_11_bits_uop_prs2;
      5'b01100:
        casez_tmp_248 = stq_12_bits_uop_prs2;
      5'b01101:
        casez_tmp_248 = stq_13_bits_uop_prs2;
      5'b01110:
        casez_tmp_248 = stq_14_bits_uop_prs2;
      5'b01111:
        casez_tmp_248 = stq_15_bits_uop_prs2;
      5'b10000:
        casez_tmp_248 = stq_16_bits_uop_prs2;
      5'b10001:
        casez_tmp_248 = stq_17_bits_uop_prs2;
      5'b10010:
        casez_tmp_248 = stq_18_bits_uop_prs2;
      5'b10011:
        casez_tmp_248 = stq_19_bits_uop_prs2;
      5'b10100:
        casez_tmp_248 = stq_20_bits_uop_prs2;
      5'b10101:
        casez_tmp_248 = stq_21_bits_uop_prs2;
      5'b10110:
        casez_tmp_248 = stq_22_bits_uop_prs2;
      5'b10111:
        casez_tmp_248 = stq_23_bits_uop_prs2;
      5'b11000:
        casez_tmp_248 = stq_24_bits_uop_prs2;
      5'b11001:
        casez_tmp_248 = stq_25_bits_uop_prs2;
      5'b11010:
        casez_tmp_248 = stq_26_bits_uop_prs2;
      5'b11011:
        casez_tmp_248 = stq_27_bits_uop_prs2;
      5'b11100:
        casez_tmp_248 = stq_28_bits_uop_prs2;
      5'b11101:
        casez_tmp_248 = stq_29_bits_uop_prs2;
      5'b11110:
        casez_tmp_248 = stq_30_bits_uop_prs2;
      default:
        casez_tmp_248 = stq_31_bits_uop_prs2;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_249;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_249 = stq_0_bits_uop_prs3;
      5'b00001:
        casez_tmp_249 = stq_1_bits_uop_prs3;
      5'b00010:
        casez_tmp_249 = stq_2_bits_uop_prs3;
      5'b00011:
        casez_tmp_249 = stq_3_bits_uop_prs3;
      5'b00100:
        casez_tmp_249 = stq_4_bits_uop_prs3;
      5'b00101:
        casez_tmp_249 = stq_5_bits_uop_prs3;
      5'b00110:
        casez_tmp_249 = stq_6_bits_uop_prs3;
      5'b00111:
        casez_tmp_249 = stq_7_bits_uop_prs3;
      5'b01000:
        casez_tmp_249 = stq_8_bits_uop_prs3;
      5'b01001:
        casez_tmp_249 = stq_9_bits_uop_prs3;
      5'b01010:
        casez_tmp_249 = stq_10_bits_uop_prs3;
      5'b01011:
        casez_tmp_249 = stq_11_bits_uop_prs3;
      5'b01100:
        casez_tmp_249 = stq_12_bits_uop_prs3;
      5'b01101:
        casez_tmp_249 = stq_13_bits_uop_prs3;
      5'b01110:
        casez_tmp_249 = stq_14_bits_uop_prs3;
      5'b01111:
        casez_tmp_249 = stq_15_bits_uop_prs3;
      5'b10000:
        casez_tmp_249 = stq_16_bits_uop_prs3;
      5'b10001:
        casez_tmp_249 = stq_17_bits_uop_prs3;
      5'b10010:
        casez_tmp_249 = stq_18_bits_uop_prs3;
      5'b10011:
        casez_tmp_249 = stq_19_bits_uop_prs3;
      5'b10100:
        casez_tmp_249 = stq_20_bits_uop_prs3;
      5'b10101:
        casez_tmp_249 = stq_21_bits_uop_prs3;
      5'b10110:
        casez_tmp_249 = stq_22_bits_uop_prs3;
      5'b10111:
        casez_tmp_249 = stq_23_bits_uop_prs3;
      5'b11000:
        casez_tmp_249 = stq_24_bits_uop_prs3;
      5'b11001:
        casez_tmp_249 = stq_25_bits_uop_prs3;
      5'b11010:
        casez_tmp_249 = stq_26_bits_uop_prs3;
      5'b11011:
        casez_tmp_249 = stq_27_bits_uop_prs3;
      5'b11100:
        casez_tmp_249 = stq_28_bits_uop_prs3;
      5'b11101:
        casez_tmp_249 = stq_29_bits_uop_prs3;
      5'b11110:
        casez_tmp_249 = stq_30_bits_uop_prs3;
      default:
        casez_tmp_249 = stq_31_bits_uop_prs3;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_250;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_250 = stq_0_bits_uop_ppred;
      5'b00001:
        casez_tmp_250 = stq_1_bits_uop_ppred;
      5'b00010:
        casez_tmp_250 = stq_2_bits_uop_ppred;
      5'b00011:
        casez_tmp_250 = stq_3_bits_uop_ppred;
      5'b00100:
        casez_tmp_250 = stq_4_bits_uop_ppred;
      5'b00101:
        casez_tmp_250 = stq_5_bits_uop_ppred;
      5'b00110:
        casez_tmp_250 = stq_6_bits_uop_ppred;
      5'b00111:
        casez_tmp_250 = stq_7_bits_uop_ppred;
      5'b01000:
        casez_tmp_250 = stq_8_bits_uop_ppred;
      5'b01001:
        casez_tmp_250 = stq_9_bits_uop_ppred;
      5'b01010:
        casez_tmp_250 = stq_10_bits_uop_ppred;
      5'b01011:
        casez_tmp_250 = stq_11_bits_uop_ppred;
      5'b01100:
        casez_tmp_250 = stq_12_bits_uop_ppred;
      5'b01101:
        casez_tmp_250 = stq_13_bits_uop_ppred;
      5'b01110:
        casez_tmp_250 = stq_14_bits_uop_ppred;
      5'b01111:
        casez_tmp_250 = stq_15_bits_uop_ppred;
      5'b10000:
        casez_tmp_250 = stq_16_bits_uop_ppred;
      5'b10001:
        casez_tmp_250 = stq_17_bits_uop_ppred;
      5'b10010:
        casez_tmp_250 = stq_18_bits_uop_ppred;
      5'b10011:
        casez_tmp_250 = stq_19_bits_uop_ppred;
      5'b10100:
        casez_tmp_250 = stq_20_bits_uop_ppred;
      5'b10101:
        casez_tmp_250 = stq_21_bits_uop_ppred;
      5'b10110:
        casez_tmp_250 = stq_22_bits_uop_ppred;
      5'b10111:
        casez_tmp_250 = stq_23_bits_uop_ppred;
      5'b11000:
        casez_tmp_250 = stq_24_bits_uop_ppred;
      5'b11001:
        casez_tmp_250 = stq_25_bits_uop_ppred;
      5'b11010:
        casez_tmp_250 = stq_26_bits_uop_ppred;
      5'b11011:
        casez_tmp_250 = stq_27_bits_uop_ppred;
      5'b11100:
        casez_tmp_250 = stq_28_bits_uop_ppred;
      5'b11101:
        casez_tmp_250 = stq_29_bits_uop_ppred;
      5'b11110:
        casez_tmp_250 = stq_30_bits_uop_ppred;
      default:
        casez_tmp_250 = stq_31_bits_uop_ppred;
    endcase
  end // always @(*)
  reg         casez_tmp_251;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_251 = stq_0_bits_uop_prs1_busy;
      5'b00001:
        casez_tmp_251 = stq_1_bits_uop_prs1_busy;
      5'b00010:
        casez_tmp_251 = stq_2_bits_uop_prs1_busy;
      5'b00011:
        casez_tmp_251 = stq_3_bits_uop_prs1_busy;
      5'b00100:
        casez_tmp_251 = stq_4_bits_uop_prs1_busy;
      5'b00101:
        casez_tmp_251 = stq_5_bits_uop_prs1_busy;
      5'b00110:
        casez_tmp_251 = stq_6_bits_uop_prs1_busy;
      5'b00111:
        casez_tmp_251 = stq_7_bits_uop_prs1_busy;
      5'b01000:
        casez_tmp_251 = stq_8_bits_uop_prs1_busy;
      5'b01001:
        casez_tmp_251 = stq_9_bits_uop_prs1_busy;
      5'b01010:
        casez_tmp_251 = stq_10_bits_uop_prs1_busy;
      5'b01011:
        casez_tmp_251 = stq_11_bits_uop_prs1_busy;
      5'b01100:
        casez_tmp_251 = stq_12_bits_uop_prs1_busy;
      5'b01101:
        casez_tmp_251 = stq_13_bits_uop_prs1_busy;
      5'b01110:
        casez_tmp_251 = stq_14_bits_uop_prs1_busy;
      5'b01111:
        casez_tmp_251 = stq_15_bits_uop_prs1_busy;
      5'b10000:
        casez_tmp_251 = stq_16_bits_uop_prs1_busy;
      5'b10001:
        casez_tmp_251 = stq_17_bits_uop_prs1_busy;
      5'b10010:
        casez_tmp_251 = stq_18_bits_uop_prs1_busy;
      5'b10011:
        casez_tmp_251 = stq_19_bits_uop_prs1_busy;
      5'b10100:
        casez_tmp_251 = stq_20_bits_uop_prs1_busy;
      5'b10101:
        casez_tmp_251 = stq_21_bits_uop_prs1_busy;
      5'b10110:
        casez_tmp_251 = stq_22_bits_uop_prs1_busy;
      5'b10111:
        casez_tmp_251 = stq_23_bits_uop_prs1_busy;
      5'b11000:
        casez_tmp_251 = stq_24_bits_uop_prs1_busy;
      5'b11001:
        casez_tmp_251 = stq_25_bits_uop_prs1_busy;
      5'b11010:
        casez_tmp_251 = stq_26_bits_uop_prs1_busy;
      5'b11011:
        casez_tmp_251 = stq_27_bits_uop_prs1_busy;
      5'b11100:
        casez_tmp_251 = stq_28_bits_uop_prs1_busy;
      5'b11101:
        casez_tmp_251 = stq_29_bits_uop_prs1_busy;
      5'b11110:
        casez_tmp_251 = stq_30_bits_uop_prs1_busy;
      default:
        casez_tmp_251 = stq_31_bits_uop_prs1_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_252;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_252 = stq_0_bits_uop_prs2_busy;
      5'b00001:
        casez_tmp_252 = stq_1_bits_uop_prs2_busy;
      5'b00010:
        casez_tmp_252 = stq_2_bits_uop_prs2_busy;
      5'b00011:
        casez_tmp_252 = stq_3_bits_uop_prs2_busy;
      5'b00100:
        casez_tmp_252 = stq_4_bits_uop_prs2_busy;
      5'b00101:
        casez_tmp_252 = stq_5_bits_uop_prs2_busy;
      5'b00110:
        casez_tmp_252 = stq_6_bits_uop_prs2_busy;
      5'b00111:
        casez_tmp_252 = stq_7_bits_uop_prs2_busy;
      5'b01000:
        casez_tmp_252 = stq_8_bits_uop_prs2_busy;
      5'b01001:
        casez_tmp_252 = stq_9_bits_uop_prs2_busy;
      5'b01010:
        casez_tmp_252 = stq_10_bits_uop_prs2_busy;
      5'b01011:
        casez_tmp_252 = stq_11_bits_uop_prs2_busy;
      5'b01100:
        casez_tmp_252 = stq_12_bits_uop_prs2_busy;
      5'b01101:
        casez_tmp_252 = stq_13_bits_uop_prs2_busy;
      5'b01110:
        casez_tmp_252 = stq_14_bits_uop_prs2_busy;
      5'b01111:
        casez_tmp_252 = stq_15_bits_uop_prs2_busy;
      5'b10000:
        casez_tmp_252 = stq_16_bits_uop_prs2_busy;
      5'b10001:
        casez_tmp_252 = stq_17_bits_uop_prs2_busy;
      5'b10010:
        casez_tmp_252 = stq_18_bits_uop_prs2_busy;
      5'b10011:
        casez_tmp_252 = stq_19_bits_uop_prs2_busy;
      5'b10100:
        casez_tmp_252 = stq_20_bits_uop_prs2_busy;
      5'b10101:
        casez_tmp_252 = stq_21_bits_uop_prs2_busy;
      5'b10110:
        casez_tmp_252 = stq_22_bits_uop_prs2_busy;
      5'b10111:
        casez_tmp_252 = stq_23_bits_uop_prs2_busy;
      5'b11000:
        casez_tmp_252 = stq_24_bits_uop_prs2_busy;
      5'b11001:
        casez_tmp_252 = stq_25_bits_uop_prs2_busy;
      5'b11010:
        casez_tmp_252 = stq_26_bits_uop_prs2_busy;
      5'b11011:
        casez_tmp_252 = stq_27_bits_uop_prs2_busy;
      5'b11100:
        casez_tmp_252 = stq_28_bits_uop_prs2_busy;
      5'b11101:
        casez_tmp_252 = stq_29_bits_uop_prs2_busy;
      5'b11110:
        casez_tmp_252 = stq_30_bits_uop_prs2_busy;
      default:
        casez_tmp_252 = stq_31_bits_uop_prs2_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_253;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_253 = stq_0_bits_uop_prs3_busy;
      5'b00001:
        casez_tmp_253 = stq_1_bits_uop_prs3_busy;
      5'b00010:
        casez_tmp_253 = stq_2_bits_uop_prs3_busy;
      5'b00011:
        casez_tmp_253 = stq_3_bits_uop_prs3_busy;
      5'b00100:
        casez_tmp_253 = stq_4_bits_uop_prs3_busy;
      5'b00101:
        casez_tmp_253 = stq_5_bits_uop_prs3_busy;
      5'b00110:
        casez_tmp_253 = stq_6_bits_uop_prs3_busy;
      5'b00111:
        casez_tmp_253 = stq_7_bits_uop_prs3_busy;
      5'b01000:
        casez_tmp_253 = stq_8_bits_uop_prs3_busy;
      5'b01001:
        casez_tmp_253 = stq_9_bits_uop_prs3_busy;
      5'b01010:
        casez_tmp_253 = stq_10_bits_uop_prs3_busy;
      5'b01011:
        casez_tmp_253 = stq_11_bits_uop_prs3_busy;
      5'b01100:
        casez_tmp_253 = stq_12_bits_uop_prs3_busy;
      5'b01101:
        casez_tmp_253 = stq_13_bits_uop_prs3_busy;
      5'b01110:
        casez_tmp_253 = stq_14_bits_uop_prs3_busy;
      5'b01111:
        casez_tmp_253 = stq_15_bits_uop_prs3_busy;
      5'b10000:
        casez_tmp_253 = stq_16_bits_uop_prs3_busy;
      5'b10001:
        casez_tmp_253 = stq_17_bits_uop_prs3_busy;
      5'b10010:
        casez_tmp_253 = stq_18_bits_uop_prs3_busy;
      5'b10011:
        casez_tmp_253 = stq_19_bits_uop_prs3_busy;
      5'b10100:
        casez_tmp_253 = stq_20_bits_uop_prs3_busy;
      5'b10101:
        casez_tmp_253 = stq_21_bits_uop_prs3_busy;
      5'b10110:
        casez_tmp_253 = stq_22_bits_uop_prs3_busy;
      5'b10111:
        casez_tmp_253 = stq_23_bits_uop_prs3_busy;
      5'b11000:
        casez_tmp_253 = stq_24_bits_uop_prs3_busy;
      5'b11001:
        casez_tmp_253 = stq_25_bits_uop_prs3_busy;
      5'b11010:
        casez_tmp_253 = stq_26_bits_uop_prs3_busy;
      5'b11011:
        casez_tmp_253 = stq_27_bits_uop_prs3_busy;
      5'b11100:
        casez_tmp_253 = stq_28_bits_uop_prs3_busy;
      5'b11101:
        casez_tmp_253 = stq_29_bits_uop_prs3_busy;
      5'b11110:
        casez_tmp_253 = stq_30_bits_uop_prs3_busy;
      default:
        casez_tmp_253 = stq_31_bits_uop_prs3_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_254;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_254 = stq_0_bits_uop_ppred_busy;
      5'b00001:
        casez_tmp_254 = stq_1_bits_uop_ppred_busy;
      5'b00010:
        casez_tmp_254 = stq_2_bits_uop_ppred_busy;
      5'b00011:
        casez_tmp_254 = stq_3_bits_uop_ppred_busy;
      5'b00100:
        casez_tmp_254 = stq_4_bits_uop_ppred_busy;
      5'b00101:
        casez_tmp_254 = stq_5_bits_uop_ppred_busy;
      5'b00110:
        casez_tmp_254 = stq_6_bits_uop_ppred_busy;
      5'b00111:
        casez_tmp_254 = stq_7_bits_uop_ppred_busy;
      5'b01000:
        casez_tmp_254 = stq_8_bits_uop_ppred_busy;
      5'b01001:
        casez_tmp_254 = stq_9_bits_uop_ppred_busy;
      5'b01010:
        casez_tmp_254 = stq_10_bits_uop_ppred_busy;
      5'b01011:
        casez_tmp_254 = stq_11_bits_uop_ppred_busy;
      5'b01100:
        casez_tmp_254 = stq_12_bits_uop_ppred_busy;
      5'b01101:
        casez_tmp_254 = stq_13_bits_uop_ppred_busy;
      5'b01110:
        casez_tmp_254 = stq_14_bits_uop_ppred_busy;
      5'b01111:
        casez_tmp_254 = stq_15_bits_uop_ppred_busy;
      5'b10000:
        casez_tmp_254 = stq_16_bits_uop_ppred_busy;
      5'b10001:
        casez_tmp_254 = stq_17_bits_uop_ppred_busy;
      5'b10010:
        casez_tmp_254 = stq_18_bits_uop_ppred_busy;
      5'b10011:
        casez_tmp_254 = stq_19_bits_uop_ppred_busy;
      5'b10100:
        casez_tmp_254 = stq_20_bits_uop_ppred_busy;
      5'b10101:
        casez_tmp_254 = stq_21_bits_uop_ppred_busy;
      5'b10110:
        casez_tmp_254 = stq_22_bits_uop_ppred_busy;
      5'b10111:
        casez_tmp_254 = stq_23_bits_uop_ppred_busy;
      5'b11000:
        casez_tmp_254 = stq_24_bits_uop_ppred_busy;
      5'b11001:
        casez_tmp_254 = stq_25_bits_uop_ppred_busy;
      5'b11010:
        casez_tmp_254 = stq_26_bits_uop_ppred_busy;
      5'b11011:
        casez_tmp_254 = stq_27_bits_uop_ppred_busy;
      5'b11100:
        casez_tmp_254 = stq_28_bits_uop_ppred_busy;
      5'b11101:
        casez_tmp_254 = stq_29_bits_uop_ppred_busy;
      5'b11110:
        casez_tmp_254 = stq_30_bits_uop_ppred_busy;
      default:
        casez_tmp_254 = stq_31_bits_uop_ppred_busy;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_255;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_255 = stq_0_bits_uop_stale_pdst;
      5'b00001:
        casez_tmp_255 = stq_1_bits_uop_stale_pdst;
      5'b00010:
        casez_tmp_255 = stq_2_bits_uop_stale_pdst;
      5'b00011:
        casez_tmp_255 = stq_3_bits_uop_stale_pdst;
      5'b00100:
        casez_tmp_255 = stq_4_bits_uop_stale_pdst;
      5'b00101:
        casez_tmp_255 = stq_5_bits_uop_stale_pdst;
      5'b00110:
        casez_tmp_255 = stq_6_bits_uop_stale_pdst;
      5'b00111:
        casez_tmp_255 = stq_7_bits_uop_stale_pdst;
      5'b01000:
        casez_tmp_255 = stq_8_bits_uop_stale_pdst;
      5'b01001:
        casez_tmp_255 = stq_9_bits_uop_stale_pdst;
      5'b01010:
        casez_tmp_255 = stq_10_bits_uop_stale_pdst;
      5'b01011:
        casez_tmp_255 = stq_11_bits_uop_stale_pdst;
      5'b01100:
        casez_tmp_255 = stq_12_bits_uop_stale_pdst;
      5'b01101:
        casez_tmp_255 = stq_13_bits_uop_stale_pdst;
      5'b01110:
        casez_tmp_255 = stq_14_bits_uop_stale_pdst;
      5'b01111:
        casez_tmp_255 = stq_15_bits_uop_stale_pdst;
      5'b10000:
        casez_tmp_255 = stq_16_bits_uop_stale_pdst;
      5'b10001:
        casez_tmp_255 = stq_17_bits_uop_stale_pdst;
      5'b10010:
        casez_tmp_255 = stq_18_bits_uop_stale_pdst;
      5'b10011:
        casez_tmp_255 = stq_19_bits_uop_stale_pdst;
      5'b10100:
        casez_tmp_255 = stq_20_bits_uop_stale_pdst;
      5'b10101:
        casez_tmp_255 = stq_21_bits_uop_stale_pdst;
      5'b10110:
        casez_tmp_255 = stq_22_bits_uop_stale_pdst;
      5'b10111:
        casez_tmp_255 = stq_23_bits_uop_stale_pdst;
      5'b11000:
        casez_tmp_255 = stq_24_bits_uop_stale_pdst;
      5'b11001:
        casez_tmp_255 = stq_25_bits_uop_stale_pdst;
      5'b11010:
        casez_tmp_255 = stq_26_bits_uop_stale_pdst;
      5'b11011:
        casez_tmp_255 = stq_27_bits_uop_stale_pdst;
      5'b11100:
        casez_tmp_255 = stq_28_bits_uop_stale_pdst;
      5'b11101:
        casez_tmp_255 = stq_29_bits_uop_stale_pdst;
      5'b11110:
        casez_tmp_255 = stq_30_bits_uop_stale_pdst;
      default:
        casez_tmp_255 = stq_31_bits_uop_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_256;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_256 = stq_0_bits_uop_exception;
      5'b00001:
        casez_tmp_256 = stq_1_bits_uop_exception;
      5'b00010:
        casez_tmp_256 = stq_2_bits_uop_exception;
      5'b00011:
        casez_tmp_256 = stq_3_bits_uop_exception;
      5'b00100:
        casez_tmp_256 = stq_4_bits_uop_exception;
      5'b00101:
        casez_tmp_256 = stq_5_bits_uop_exception;
      5'b00110:
        casez_tmp_256 = stq_6_bits_uop_exception;
      5'b00111:
        casez_tmp_256 = stq_7_bits_uop_exception;
      5'b01000:
        casez_tmp_256 = stq_8_bits_uop_exception;
      5'b01001:
        casez_tmp_256 = stq_9_bits_uop_exception;
      5'b01010:
        casez_tmp_256 = stq_10_bits_uop_exception;
      5'b01011:
        casez_tmp_256 = stq_11_bits_uop_exception;
      5'b01100:
        casez_tmp_256 = stq_12_bits_uop_exception;
      5'b01101:
        casez_tmp_256 = stq_13_bits_uop_exception;
      5'b01110:
        casez_tmp_256 = stq_14_bits_uop_exception;
      5'b01111:
        casez_tmp_256 = stq_15_bits_uop_exception;
      5'b10000:
        casez_tmp_256 = stq_16_bits_uop_exception;
      5'b10001:
        casez_tmp_256 = stq_17_bits_uop_exception;
      5'b10010:
        casez_tmp_256 = stq_18_bits_uop_exception;
      5'b10011:
        casez_tmp_256 = stq_19_bits_uop_exception;
      5'b10100:
        casez_tmp_256 = stq_20_bits_uop_exception;
      5'b10101:
        casez_tmp_256 = stq_21_bits_uop_exception;
      5'b10110:
        casez_tmp_256 = stq_22_bits_uop_exception;
      5'b10111:
        casez_tmp_256 = stq_23_bits_uop_exception;
      5'b11000:
        casez_tmp_256 = stq_24_bits_uop_exception;
      5'b11001:
        casez_tmp_256 = stq_25_bits_uop_exception;
      5'b11010:
        casez_tmp_256 = stq_26_bits_uop_exception;
      5'b11011:
        casez_tmp_256 = stq_27_bits_uop_exception;
      5'b11100:
        casez_tmp_256 = stq_28_bits_uop_exception;
      5'b11101:
        casez_tmp_256 = stq_29_bits_uop_exception;
      5'b11110:
        casez_tmp_256 = stq_30_bits_uop_exception;
      default:
        casez_tmp_256 = stq_31_bits_uop_exception;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_257;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_257 = stq_0_bits_uop_exc_cause;
      5'b00001:
        casez_tmp_257 = stq_1_bits_uop_exc_cause;
      5'b00010:
        casez_tmp_257 = stq_2_bits_uop_exc_cause;
      5'b00011:
        casez_tmp_257 = stq_3_bits_uop_exc_cause;
      5'b00100:
        casez_tmp_257 = stq_4_bits_uop_exc_cause;
      5'b00101:
        casez_tmp_257 = stq_5_bits_uop_exc_cause;
      5'b00110:
        casez_tmp_257 = stq_6_bits_uop_exc_cause;
      5'b00111:
        casez_tmp_257 = stq_7_bits_uop_exc_cause;
      5'b01000:
        casez_tmp_257 = stq_8_bits_uop_exc_cause;
      5'b01001:
        casez_tmp_257 = stq_9_bits_uop_exc_cause;
      5'b01010:
        casez_tmp_257 = stq_10_bits_uop_exc_cause;
      5'b01011:
        casez_tmp_257 = stq_11_bits_uop_exc_cause;
      5'b01100:
        casez_tmp_257 = stq_12_bits_uop_exc_cause;
      5'b01101:
        casez_tmp_257 = stq_13_bits_uop_exc_cause;
      5'b01110:
        casez_tmp_257 = stq_14_bits_uop_exc_cause;
      5'b01111:
        casez_tmp_257 = stq_15_bits_uop_exc_cause;
      5'b10000:
        casez_tmp_257 = stq_16_bits_uop_exc_cause;
      5'b10001:
        casez_tmp_257 = stq_17_bits_uop_exc_cause;
      5'b10010:
        casez_tmp_257 = stq_18_bits_uop_exc_cause;
      5'b10011:
        casez_tmp_257 = stq_19_bits_uop_exc_cause;
      5'b10100:
        casez_tmp_257 = stq_20_bits_uop_exc_cause;
      5'b10101:
        casez_tmp_257 = stq_21_bits_uop_exc_cause;
      5'b10110:
        casez_tmp_257 = stq_22_bits_uop_exc_cause;
      5'b10111:
        casez_tmp_257 = stq_23_bits_uop_exc_cause;
      5'b11000:
        casez_tmp_257 = stq_24_bits_uop_exc_cause;
      5'b11001:
        casez_tmp_257 = stq_25_bits_uop_exc_cause;
      5'b11010:
        casez_tmp_257 = stq_26_bits_uop_exc_cause;
      5'b11011:
        casez_tmp_257 = stq_27_bits_uop_exc_cause;
      5'b11100:
        casez_tmp_257 = stq_28_bits_uop_exc_cause;
      5'b11101:
        casez_tmp_257 = stq_29_bits_uop_exc_cause;
      5'b11110:
        casez_tmp_257 = stq_30_bits_uop_exc_cause;
      default:
        casez_tmp_257 = stq_31_bits_uop_exc_cause;
    endcase
  end // always @(*)
  reg         casez_tmp_258;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_258 = stq_0_bits_uop_bypassable;
      5'b00001:
        casez_tmp_258 = stq_1_bits_uop_bypassable;
      5'b00010:
        casez_tmp_258 = stq_2_bits_uop_bypassable;
      5'b00011:
        casez_tmp_258 = stq_3_bits_uop_bypassable;
      5'b00100:
        casez_tmp_258 = stq_4_bits_uop_bypassable;
      5'b00101:
        casez_tmp_258 = stq_5_bits_uop_bypassable;
      5'b00110:
        casez_tmp_258 = stq_6_bits_uop_bypassable;
      5'b00111:
        casez_tmp_258 = stq_7_bits_uop_bypassable;
      5'b01000:
        casez_tmp_258 = stq_8_bits_uop_bypassable;
      5'b01001:
        casez_tmp_258 = stq_9_bits_uop_bypassable;
      5'b01010:
        casez_tmp_258 = stq_10_bits_uop_bypassable;
      5'b01011:
        casez_tmp_258 = stq_11_bits_uop_bypassable;
      5'b01100:
        casez_tmp_258 = stq_12_bits_uop_bypassable;
      5'b01101:
        casez_tmp_258 = stq_13_bits_uop_bypassable;
      5'b01110:
        casez_tmp_258 = stq_14_bits_uop_bypassable;
      5'b01111:
        casez_tmp_258 = stq_15_bits_uop_bypassable;
      5'b10000:
        casez_tmp_258 = stq_16_bits_uop_bypassable;
      5'b10001:
        casez_tmp_258 = stq_17_bits_uop_bypassable;
      5'b10010:
        casez_tmp_258 = stq_18_bits_uop_bypassable;
      5'b10011:
        casez_tmp_258 = stq_19_bits_uop_bypassable;
      5'b10100:
        casez_tmp_258 = stq_20_bits_uop_bypassable;
      5'b10101:
        casez_tmp_258 = stq_21_bits_uop_bypassable;
      5'b10110:
        casez_tmp_258 = stq_22_bits_uop_bypassable;
      5'b10111:
        casez_tmp_258 = stq_23_bits_uop_bypassable;
      5'b11000:
        casez_tmp_258 = stq_24_bits_uop_bypassable;
      5'b11001:
        casez_tmp_258 = stq_25_bits_uop_bypassable;
      5'b11010:
        casez_tmp_258 = stq_26_bits_uop_bypassable;
      5'b11011:
        casez_tmp_258 = stq_27_bits_uop_bypassable;
      5'b11100:
        casez_tmp_258 = stq_28_bits_uop_bypassable;
      5'b11101:
        casez_tmp_258 = stq_29_bits_uop_bypassable;
      5'b11110:
        casez_tmp_258 = stq_30_bits_uop_bypassable;
      default:
        casez_tmp_258 = stq_31_bits_uop_bypassable;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_259;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_259 = stq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_259 = stq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_259 = stq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_259 = stq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_259 = stq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_259 = stq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_259 = stq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_259 = stq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_259 = stq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_259 = stq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_259 = stq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_259 = stq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_259 = stq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_259 = stq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_259 = stq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_259 = stq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_259 = stq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_259 = stq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_259 = stq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_259 = stq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_259 = stq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_259 = stq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_259 = stq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_259 = stq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_259 = stq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_259 = stq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_259 = stq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_259 = stq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_259 = stq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_259 = stq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_259 = stq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_259 = stq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_260;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_260 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_260 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_260 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_260 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_260 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_260 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_260 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_260 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_260 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_260 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_260 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_260 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_260 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_260 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_260 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_260 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_260 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_260 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_260 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_260 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_260 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_260 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_260 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_260 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_260 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_260 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_260 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_260 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_260 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_260 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_260 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_260 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_261;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_261 = stq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_261 = stq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_261 = stq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_261 = stq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_261 = stq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_261 = stq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_261 = stq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_261 = stq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_261 = stq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_261 = stq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_261 = stq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_261 = stq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_261 = stq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_261 = stq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_261 = stq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_261 = stq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_261 = stq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_261 = stq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_261 = stq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_261 = stq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_261 = stq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_261 = stq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_261 = stq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_261 = stq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_261 = stq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_261 = stq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_261 = stq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_261 = stq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_261 = stq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_261 = stq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_261 = stq_30_bits_uop_mem_signed;
      default:
        casez_tmp_261 = stq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  reg         casez_tmp_262;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_262 = stq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_262 = stq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_262 = stq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_262 = stq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_262 = stq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_262 = stq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_262 = stq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_262 = stq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_262 = stq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_262 = stq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_262 = stq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_262 = stq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_262 = stq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_262 = stq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_262 = stq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_262 = stq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_262 = stq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_262 = stq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_262 = stq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_262 = stq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_262 = stq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_262 = stq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_262 = stq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_262 = stq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_262 = stq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_262 = stq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_262 = stq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_262 = stq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_262 = stq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_262 = stq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_262 = stq_30_bits_uop_is_fence;
      default:
        casez_tmp_262 = stq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  reg         casez_tmp_263;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_263 = stq_0_bits_uop_is_fencei;
      5'b00001:
        casez_tmp_263 = stq_1_bits_uop_is_fencei;
      5'b00010:
        casez_tmp_263 = stq_2_bits_uop_is_fencei;
      5'b00011:
        casez_tmp_263 = stq_3_bits_uop_is_fencei;
      5'b00100:
        casez_tmp_263 = stq_4_bits_uop_is_fencei;
      5'b00101:
        casez_tmp_263 = stq_5_bits_uop_is_fencei;
      5'b00110:
        casez_tmp_263 = stq_6_bits_uop_is_fencei;
      5'b00111:
        casez_tmp_263 = stq_7_bits_uop_is_fencei;
      5'b01000:
        casez_tmp_263 = stq_8_bits_uop_is_fencei;
      5'b01001:
        casez_tmp_263 = stq_9_bits_uop_is_fencei;
      5'b01010:
        casez_tmp_263 = stq_10_bits_uop_is_fencei;
      5'b01011:
        casez_tmp_263 = stq_11_bits_uop_is_fencei;
      5'b01100:
        casez_tmp_263 = stq_12_bits_uop_is_fencei;
      5'b01101:
        casez_tmp_263 = stq_13_bits_uop_is_fencei;
      5'b01110:
        casez_tmp_263 = stq_14_bits_uop_is_fencei;
      5'b01111:
        casez_tmp_263 = stq_15_bits_uop_is_fencei;
      5'b10000:
        casez_tmp_263 = stq_16_bits_uop_is_fencei;
      5'b10001:
        casez_tmp_263 = stq_17_bits_uop_is_fencei;
      5'b10010:
        casez_tmp_263 = stq_18_bits_uop_is_fencei;
      5'b10011:
        casez_tmp_263 = stq_19_bits_uop_is_fencei;
      5'b10100:
        casez_tmp_263 = stq_20_bits_uop_is_fencei;
      5'b10101:
        casez_tmp_263 = stq_21_bits_uop_is_fencei;
      5'b10110:
        casez_tmp_263 = stq_22_bits_uop_is_fencei;
      5'b10111:
        casez_tmp_263 = stq_23_bits_uop_is_fencei;
      5'b11000:
        casez_tmp_263 = stq_24_bits_uop_is_fencei;
      5'b11001:
        casez_tmp_263 = stq_25_bits_uop_is_fencei;
      5'b11010:
        casez_tmp_263 = stq_26_bits_uop_is_fencei;
      5'b11011:
        casez_tmp_263 = stq_27_bits_uop_is_fencei;
      5'b11100:
        casez_tmp_263 = stq_28_bits_uop_is_fencei;
      5'b11101:
        casez_tmp_263 = stq_29_bits_uop_is_fencei;
      5'b11110:
        casez_tmp_263 = stq_30_bits_uop_is_fencei;
      default:
        casez_tmp_263 = stq_31_bits_uop_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_264;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_264 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_264 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_264 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_264 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_264 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_264 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_264 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_264 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_264 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_264 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_264 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_264 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_264 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_264 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_264 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_264 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_264 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_264 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_264 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_264 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_264 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_264 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_264 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_264 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_264 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_264 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_264 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_264 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_264 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_264 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_264 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_264 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_265;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_265 = stq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_265 = stq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_265 = stq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_265 = stq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_265 = stq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_265 = stq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_265 = stq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_265 = stq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_265 = stq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_265 = stq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_265 = stq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_265 = stq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_265 = stq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_265 = stq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_265 = stq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_265 = stq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_265 = stq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_265 = stq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_265 = stq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_265 = stq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_265 = stq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_265 = stq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_265 = stq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_265 = stq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_265 = stq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_265 = stq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_265 = stq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_265 = stq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_265 = stq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_265 = stq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_265 = stq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_265 = stq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_266;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_266 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_266 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_266 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_266 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_266 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_266 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_266 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_266 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_266 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_266 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_266 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_266 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_266 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_266 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_266 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_266 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_266 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_266 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_266 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_266 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_266 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_266 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_266 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_266 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_266 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_266 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_266 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_266 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_266 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_266 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_266 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_266 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_267;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_267 = stq_0_bits_uop_is_sys_pc2epc;
      5'b00001:
        casez_tmp_267 = stq_1_bits_uop_is_sys_pc2epc;
      5'b00010:
        casez_tmp_267 = stq_2_bits_uop_is_sys_pc2epc;
      5'b00011:
        casez_tmp_267 = stq_3_bits_uop_is_sys_pc2epc;
      5'b00100:
        casez_tmp_267 = stq_4_bits_uop_is_sys_pc2epc;
      5'b00101:
        casez_tmp_267 = stq_5_bits_uop_is_sys_pc2epc;
      5'b00110:
        casez_tmp_267 = stq_6_bits_uop_is_sys_pc2epc;
      5'b00111:
        casez_tmp_267 = stq_7_bits_uop_is_sys_pc2epc;
      5'b01000:
        casez_tmp_267 = stq_8_bits_uop_is_sys_pc2epc;
      5'b01001:
        casez_tmp_267 = stq_9_bits_uop_is_sys_pc2epc;
      5'b01010:
        casez_tmp_267 = stq_10_bits_uop_is_sys_pc2epc;
      5'b01011:
        casez_tmp_267 = stq_11_bits_uop_is_sys_pc2epc;
      5'b01100:
        casez_tmp_267 = stq_12_bits_uop_is_sys_pc2epc;
      5'b01101:
        casez_tmp_267 = stq_13_bits_uop_is_sys_pc2epc;
      5'b01110:
        casez_tmp_267 = stq_14_bits_uop_is_sys_pc2epc;
      5'b01111:
        casez_tmp_267 = stq_15_bits_uop_is_sys_pc2epc;
      5'b10000:
        casez_tmp_267 = stq_16_bits_uop_is_sys_pc2epc;
      5'b10001:
        casez_tmp_267 = stq_17_bits_uop_is_sys_pc2epc;
      5'b10010:
        casez_tmp_267 = stq_18_bits_uop_is_sys_pc2epc;
      5'b10011:
        casez_tmp_267 = stq_19_bits_uop_is_sys_pc2epc;
      5'b10100:
        casez_tmp_267 = stq_20_bits_uop_is_sys_pc2epc;
      5'b10101:
        casez_tmp_267 = stq_21_bits_uop_is_sys_pc2epc;
      5'b10110:
        casez_tmp_267 = stq_22_bits_uop_is_sys_pc2epc;
      5'b10111:
        casez_tmp_267 = stq_23_bits_uop_is_sys_pc2epc;
      5'b11000:
        casez_tmp_267 = stq_24_bits_uop_is_sys_pc2epc;
      5'b11001:
        casez_tmp_267 = stq_25_bits_uop_is_sys_pc2epc;
      5'b11010:
        casez_tmp_267 = stq_26_bits_uop_is_sys_pc2epc;
      5'b11011:
        casez_tmp_267 = stq_27_bits_uop_is_sys_pc2epc;
      5'b11100:
        casez_tmp_267 = stq_28_bits_uop_is_sys_pc2epc;
      5'b11101:
        casez_tmp_267 = stq_29_bits_uop_is_sys_pc2epc;
      5'b11110:
        casez_tmp_267 = stq_30_bits_uop_is_sys_pc2epc;
      default:
        casez_tmp_267 = stq_31_bits_uop_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_268;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_268 = stq_0_bits_uop_is_unique;
      5'b00001:
        casez_tmp_268 = stq_1_bits_uop_is_unique;
      5'b00010:
        casez_tmp_268 = stq_2_bits_uop_is_unique;
      5'b00011:
        casez_tmp_268 = stq_3_bits_uop_is_unique;
      5'b00100:
        casez_tmp_268 = stq_4_bits_uop_is_unique;
      5'b00101:
        casez_tmp_268 = stq_5_bits_uop_is_unique;
      5'b00110:
        casez_tmp_268 = stq_6_bits_uop_is_unique;
      5'b00111:
        casez_tmp_268 = stq_7_bits_uop_is_unique;
      5'b01000:
        casez_tmp_268 = stq_8_bits_uop_is_unique;
      5'b01001:
        casez_tmp_268 = stq_9_bits_uop_is_unique;
      5'b01010:
        casez_tmp_268 = stq_10_bits_uop_is_unique;
      5'b01011:
        casez_tmp_268 = stq_11_bits_uop_is_unique;
      5'b01100:
        casez_tmp_268 = stq_12_bits_uop_is_unique;
      5'b01101:
        casez_tmp_268 = stq_13_bits_uop_is_unique;
      5'b01110:
        casez_tmp_268 = stq_14_bits_uop_is_unique;
      5'b01111:
        casez_tmp_268 = stq_15_bits_uop_is_unique;
      5'b10000:
        casez_tmp_268 = stq_16_bits_uop_is_unique;
      5'b10001:
        casez_tmp_268 = stq_17_bits_uop_is_unique;
      5'b10010:
        casez_tmp_268 = stq_18_bits_uop_is_unique;
      5'b10011:
        casez_tmp_268 = stq_19_bits_uop_is_unique;
      5'b10100:
        casez_tmp_268 = stq_20_bits_uop_is_unique;
      5'b10101:
        casez_tmp_268 = stq_21_bits_uop_is_unique;
      5'b10110:
        casez_tmp_268 = stq_22_bits_uop_is_unique;
      5'b10111:
        casez_tmp_268 = stq_23_bits_uop_is_unique;
      5'b11000:
        casez_tmp_268 = stq_24_bits_uop_is_unique;
      5'b11001:
        casez_tmp_268 = stq_25_bits_uop_is_unique;
      5'b11010:
        casez_tmp_268 = stq_26_bits_uop_is_unique;
      5'b11011:
        casez_tmp_268 = stq_27_bits_uop_is_unique;
      5'b11100:
        casez_tmp_268 = stq_28_bits_uop_is_unique;
      5'b11101:
        casez_tmp_268 = stq_29_bits_uop_is_unique;
      5'b11110:
        casez_tmp_268 = stq_30_bits_uop_is_unique;
      default:
        casez_tmp_268 = stq_31_bits_uop_is_unique;
    endcase
  end // always @(*)
  reg         casez_tmp_269;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_269 = stq_0_bits_uop_flush_on_commit;
      5'b00001:
        casez_tmp_269 = stq_1_bits_uop_flush_on_commit;
      5'b00010:
        casez_tmp_269 = stq_2_bits_uop_flush_on_commit;
      5'b00011:
        casez_tmp_269 = stq_3_bits_uop_flush_on_commit;
      5'b00100:
        casez_tmp_269 = stq_4_bits_uop_flush_on_commit;
      5'b00101:
        casez_tmp_269 = stq_5_bits_uop_flush_on_commit;
      5'b00110:
        casez_tmp_269 = stq_6_bits_uop_flush_on_commit;
      5'b00111:
        casez_tmp_269 = stq_7_bits_uop_flush_on_commit;
      5'b01000:
        casez_tmp_269 = stq_8_bits_uop_flush_on_commit;
      5'b01001:
        casez_tmp_269 = stq_9_bits_uop_flush_on_commit;
      5'b01010:
        casez_tmp_269 = stq_10_bits_uop_flush_on_commit;
      5'b01011:
        casez_tmp_269 = stq_11_bits_uop_flush_on_commit;
      5'b01100:
        casez_tmp_269 = stq_12_bits_uop_flush_on_commit;
      5'b01101:
        casez_tmp_269 = stq_13_bits_uop_flush_on_commit;
      5'b01110:
        casez_tmp_269 = stq_14_bits_uop_flush_on_commit;
      5'b01111:
        casez_tmp_269 = stq_15_bits_uop_flush_on_commit;
      5'b10000:
        casez_tmp_269 = stq_16_bits_uop_flush_on_commit;
      5'b10001:
        casez_tmp_269 = stq_17_bits_uop_flush_on_commit;
      5'b10010:
        casez_tmp_269 = stq_18_bits_uop_flush_on_commit;
      5'b10011:
        casez_tmp_269 = stq_19_bits_uop_flush_on_commit;
      5'b10100:
        casez_tmp_269 = stq_20_bits_uop_flush_on_commit;
      5'b10101:
        casez_tmp_269 = stq_21_bits_uop_flush_on_commit;
      5'b10110:
        casez_tmp_269 = stq_22_bits_uop_flush_on_commit;
      5'b10111:
        casez_tmp_269 = stq_23_bits_uop_flush_on_commit;
      5'b11000:
        casez_tmp_269 = stq_24_bits_uop_flush_on_commit;
      5'b11001:
        casez_tmp_269 = stq_25_bits_uop_flush_on_commit;
      5'b11010:
        casez_tmp_269 = stq_26_bits_uop_flush_on_commit;
      5'b11011:
        casez_tmp_269 = stq_27_bits_uop_flush_on_commit;
      5'b11100:
        casez_tmp_269 = stq_28_bits_uop_flush_on_commit;
      5'b11101:
        casez_tmp_269 = stq_29_bits_uop_flush_on_commit;
      5'b11110:
        casez_tmp_269 = stq_30_bits_uop_flush_on_commit;
      default:
        casez_tmp_269 = stq_31_bits_uop_flush_on_commit;
    endcase
  end // always @(*)
  reg         casez_tmp_270;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_270 = stq_0_bits_uop_ldst_is_rs1;
      5'b00001:
        casez_tmp_270 = stq_1_bits_uop_ldst_is_rs1;
      5'b00010:
        casez_tmp_270 = stq_2_bits_uop_ldst_is_rs1;
      5'b00011:
        casez_tmp_270 = stq_3_bits_uop_ldst_is_rs1;
      5'b00100:
        casez_tmp_270 = stq_4_bits_uop_ldst_is_rs1;
      5'b00101:
        casez_tmp_270 = stq_5_bits_uop_ldst_is_rs1;
      5'b00110:
        casez_tmp_270 = stq_6_bits_uop_ldst_is_rs1;
      5'b00111:
        casez_tmp_270 = stq_7_bits_uop_ldst_is_rs1;
      5'b01000:
        casez_tmp_270 = stq_8_bits_uop_ldst_is_rs1;
      5'b01001:
        casez_tmp_270 = stq_9_bits_uop_ldst_is_rs1;
      5'b01010:
        casez_tmp_270 = stq_10_bits_uop_ldst_is_rs1;
      5'b01011:
        casez_tmp_270 = stq_11_bits_uop_ldst_is_rs1;
      5'b01100:
        casez_tmp_270 = stq_12_bits_uop_ldst_is_rs1;
      5'b01101:
        casez_tmp_270 = stq_13_bits_uop_ldst_is_rs1;
      5'b01110:
        casez_tmp_270 = stq_14_bits_uop_ldst_is_rs1;
      5'b01111:
        casez_tmp_270 = stq_15_bits_uop_ldst_is_rs1;
      5'b10000:
        casez_tmp_270 = stq_16_bits_uop_ldst_is_rs1;
      5'b10001:
        casez_tmp_270 = stq_17_bits_uop_ldst_is_rs1;
      5'b10010:
        casez_tmp_270 = stq_18_bits_uop_ldst_is_rs1;
      5'b10011:
        casez_tmp_270 = stq_19_bits_uop_ldst_is_rs1;
      5'b10100:
        casez_tmp_270 = stq_20_bits_uop_ldst_is_rs1;
      5'b10101:
        casez_tmp_270 = stq_21_bits_uop_ldst_is_rs1;
      5'b10110:
        casez_tmp_270 = stq_22_bits_uop_ldst_is_rs1;
      5'b10111:
        casez_tmp_270 = stq_23_bits_uop_ldst_is_rs1;
      5'b11000:
        casez_tmp_270 = stq_24_bits_uop_ldst_is_rs1;
      5'b11001:
        casez_tmp_270 = stq_25_bits_uop_ldst_is_rs1;
      5'b11010:
        casez_tmp_270 = stq_26_bits_uop_ldst_is_rs1;
      5'b11011:
        casez_tmp_270 = stq_27_bits_uop_ldst_is_rs1;
      5'b11100:
        casez_tmp_270 = stq_28_bits_uop_ldst_is_rs1;
      5'b11101:
        casez_tmp_270 = stq_29_bits_uop_ldst_is_rs1;
      5'b11110:
        casez_tmp_270 = stq_30_bits_uop_ldst_is_rs1;
      default:
        casez_tmp_270 = stq_31_bits_uop_ldst_is_rs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_271;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_271 = stq_0_bits_uop_ldst;
      5'b00001:
        casez_tmp_271 = stq_1_bits_uop_ldst;
      5'b00010:
        casez_tmp_271 = stq_2_bits_uop_ldst;
      5'b00011:
        casez_tmp_271 = stq_3_bits_uop_ldst;
      5'b00100:
        casez_tmp_271 = stq_4_bits_uop_ldst;
      5'b00101:
        casez_tmp_271 = stq_5_bits_uop_ldst;
      5'b00110:
        casez_tmp_271 = stq_6_bits_uop_ldst;
      5'b00111:
        casez_tmp_271 = stq_7_bits_uop_ldst;
      5'b01000:
        casez_tmp_271 = stq_8_bits_uop_ldst;
      5'b01001:
        casez_tmp_271 = stq_9_bits_uop_ldst;
      5'b01010:
        casez_tmp_271 = stq_10_bits_uop_ldst;
      5'b01011:
        casez_tmp_271 = stq_11_bits_uop_ldst;
      5'b01100:
        casez_tmp_271 = stq_12_bits_uop_ldst;
      5'b01101:
        casez_tmp_271 = stq_13_bits_uop_ldst;
      5'b01110:
        casez_tmp_271 = stq_14_bits_uop_ldst;
      5'b01111:
        casez_tmp_271 = stq_15_bits_uop_ldst;
      5'b10000:
        casez_tmp_271 = stq_16_bits_uop_ldst;
      5'b10001:
        casez_tmp_271 = stq_17_bits_uop_ldst;
      5'b10010:
        casez_tmp_271 = stq_18_bits_uop_ldst;
      5'b10011:
        casez_tmp_271 = stq_19_bits_uop_ldst;
      5'b10100:
        casez_tmp_271 = stq_20_bits_uop_ldst;
      5'b10101:
        casez_tmp_271 = stq_21_bits_uop_ldst;
      5'b10110:
        casez_tmp_271 = stq_22_bits_uop_ldst;
      5'b10111:
        casez_tmp_271 = stq_23_bits_uop_ldst;
      5'b11000:
        casez_tmp_271 = stq_24_bits_uop_ldst;
      5'b11001:
        casez_tmp_271 = stq_25_bits_uop_ldst;
      5'b11010:
        casez_tmp_271 = stq_26_bits_uop_ldst;
      5'b11011:
        casez_tmp_271 = stq_27_bits_uop_ldst;
      5'b11100:
        casez_tmp_271 = stq_28_bits_uop_ldst;
      5'b11101:
        casez_tmp_271 = stq_29_bits_uop_ldst;
      5'b11110:
        casez_tmp_271 = stq_30_bits_uop_ldst;
      default:
        casez_tmp_271 = stq_31_bits_uop_ldst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_272;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_272 = stq_0_bits_uop_lrs1;
      5'b00001:
        casez_tmp_272 = stq_1_bits_uop_lrs1;
      5'b00010:
        casez_tmp_272 = stq_2_bits_uop_lrs1;
      5'b00011:
        casez_tmp_272 = stq_3_bits_uop_lrs1;
      5'b00100:
        casez_tmp_272 = stq_4_bits_uop_lrs1;
      5'b00101:
        casez_tmp_272 = stq_5_bits_uop_lrs1;
      5'b00110:
        casez_tmp_272 = stq_6_bits_uop_lrs1;
      5'b00111:
        casez_tmp_272 = stq_7_bits_uop_lrs1;
      5'b01000:
        casez_tmp_272 = stq_8_bits_uop_lrs1;
      5'b01001:
        casez_tmp_272 = stq_9_bits_uop_lrs1;
      5'b01010:
        casez_tmp_272 = stq_10_bits_uop_lrs1;
      5'b01011:
        casez_tmp_272 = stq_11_bits_uop_lrs1;
      5'b01100:
        casez_tmp_272 = stq_12_bits_uop_lrs1;
      5'b01101:
        casez_tmp_272 = stq_13_bits_uop_lrs1;
      5'b01110:
        casez_tmp_272 = stq_14_bits_uop_lrs1;
      5'b01111:
        casez_tmp_272 = stq_15_bits_uop_lrs1;
      5'b10000:
        casez_tmp_272 = stq_16_bits_uop_lrs1;
      5'b10001:
        casez_tmp_272 = stq_17_bits_uop_lrs1;
      5'b10010:
        casez_tmp_272 = stq_18_bits_uop_lrs1;
      5'b10011:
        casez_tmp_272 = stq_19_bits_uop_lrs1;
      5'b10100:
        casez_tmp_272 = stq_20_bits_uop_lrs1;
      5'b10101:
        casez_tmp_272 = stq_21_bits_uop_lrs1;
      5'b10110:
        casez_tmp_272 = stq_22_bits_uop_lrs1;
      5'b10111:
        casez_tmp_272 = stq_23_bits_uop_lrs1;
      5'b11000:
        casez_tmp_272 = stq_24_bits_uop_lrs1;
      5'b11001:
        casez_tmp_272 = stq_25_bits_uop_lrs1;
      5'b11010:
        casez_tmp_272 = stq_26_bits_uop_lrs1;
      5'b11011:
        casez_tmp_272 = stq_27_bits_uop_lrs1;
      5'b11100:
        casez_tmp_272 = stq_28_bits_uop_lrs1;
      5'b11101:
        casez_tmp_272 = stq_29_bits_uop_lrs1;
      5'b11110:
        casez_tmp_272 = stq_30_bits_uop_lrs1;
      default:
        casez_tmp_272 = stq_31_bits_uop_lrs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_273;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_273 = stq_0_bits_uop_lrs2;
      5'b00001:
        casez_tmp_273 = stq_1_bits_uop_lrs2;
      5'b00010:
        casez_tmp_273 = stq_2_bits_uop_lrs2;
      5'b00011:
        casez_tmp_273 = stq_3_bits_uop_lrs2;
      5'b00100:
        casez_tmp_273 = stq_4_bits_uop_lrs2;
      5'b00101:
        casez_tmp_273 = stq_5_bits_uop_lrs2;
      5'b00110:
        casez_tmp_273 = stq_6_bits_uop_lrs2;
      5'b00111:
        casez_tmp_273 = stq_7_bits_uop_lrs2;
      5'b01000:
        casez_tmp_273 = stq_8_bits_uop_lrs2;
      5'b01001:
        casez_tmp_273 = stq_9_bits_uop_lrs2;
      5'b01010:
        casez_tmp_273 = stq_10_bits_uop_lrs2;
      5'b01011:
        casez_tmp_273 = stq_11_bits_uop_lrs2;
      5'b01100:
        casez_tmp_273 = stq_12_bits_uop_lrs2;
      5'b01101:
        casez_tmp_273 = stq_13_bits_uop_lrs2;
      5'b01110:
        casez_tmp_273 = stq_14_bits_uop_lrs2;
      5'b01111:
        casez_tmp_273 = stq_15_bits_uop_lrs2;
      5'b10000:
        casez_tmp_273 = stq_16_bits_uop_lrs2;
      5'b10001:
        casez_tmp_273 = stq_17_bits_uop_lrs2;
      5'b10010:
        casez_tmp_273 = stq_18_bits_uop_lrs2;
      5'b10011:
        casez_tmp_273 = stq_19_bits_uop_lrs2;
      5'b10100:
        casez_tmp_273 = stq_20_bits_uop_lrs2;
      5'b10101:
        casez_tmp_273 = stq_21_bits_uop_lrs2;
      5'b10110:
        casez_tmp_273 = stq_22_bits_uop_lrs2;
      5'b10111:
        casez_tmp_273 = stq_23_bits_uop_lrs2;
      5'b11000:
        casez_tmp_273 = stq_24_bits_uop_lrs2;
      5'b11001:
        casez_tmp_273 = stq_25_bits_uop_lrs2;
      5'b11010:
        casez_tmp_273 = stq_26_bits_uop_lrs2;
      5'b11011:
        casez_tmp_273 = stq_27_bits_uop_lrs2;
      5'b11100:
        casez_tmp_273 = stq_28_bits_uop_lrs2;
      5'b11101:
        casez_tmp_273 = stq_29_bits_uop_lrs2;
      5'b11110:
        casez_tmp_273 = stq_30_bits_uop_lrs2;
      default:
        casez_tmp_273 = stq_31_bits_uop_lrs2;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_274;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_274 = stq_0_bits_uop_lrs3;
      5'b00001:
        casez_tmp_274 = stq_1_bits_uop_lrs3;
      5'b00010:
        casez_tmp_274 = stq_2_bits_uop_lrs3;
      5'b00011:
        casez_tmp_274 = stq_3_bits_uop_lrs3;
      5'b00100:
        casez_tmp_274 = stq_4_bits_uop_lrs3;
      5'b00101:
        casez_tmp_274 = stq_5_bits_uop_lrs3;
      5'b00110:
        casez_tmp_274 = stq_6_bits_uop_lrs3;
      5'b00111:
        casez_tmp_274 = stq_7_bits_uop_lrs3;
      5'b01000:
        casez_tmp_274 = stq_8_bits_uop_lrs3;
      5'b01001:
        casez_tmp_274 = stq_9_bits_uop_lrs3;
      5'b01010:
        casez_tmp_274 = stq_10_bits_uop_lrs3;
      5'b01011:
        casez_tmp_274 = stq_11_bits_uop_lrs3;
      5'b01100:
        casez_tmp_274 = stq_12_bits_uop_lrs3;
      5'b01101:
        casez_tmp_274 = stq_13_bits_uop_lrs3;
      5'b01110:
        casez_tmp_274 = stq_14_bits_uop_lrs3;
      5'b01111:
        casez_tmp_274 = stq_15_bits_uop_lrs3;
      5'b10000:
        casez_tmp_274 = stq_16_bits_uop_lrs3;
      5'b10001:
        casez_tmp_274 = stq_17_bits_uop_lrs3;
      5'b10010:
        casez_tmp_274 = stq_18_bits_uop_lrs3;
      5'b10011:
        casez_tmp_274 = stq_19_bits_uop_lrs3;
      5'b10100:
        casez_tmp_274 = stq_20_bits_uop_lrs3;
      5'b10101:
        casez_tmp_274 = stq_21_bits_uop_lrs3;
      5'b10110:
        casez_tmp_274 = stq_22_bits_uop_lrs3;
      5'b10111:
        casez_tmp_274 = stq_23_bits_uop_lrs3;
      5'b11000:
        casez_tmp_274 = stq_24_bits_uop_lrs3;
      5'b11001:
        casez_tmp_274 = stq_25_bits_uop_lrs3;
      5'b11010:
        casez_tmp_274 = stq_26_bits_uop_lrs3;
      5'b11011:
        casez_tmp_274 = stq_27_bits_uop_lrs3;
      5'b11100:
        casez_tmp_274 = stq_28_bits_uop_lrs3;
      5'b11101:
        casez_tmp_274 = stq_29_bits_uop_lrs3;
      5'b11110:
        casez_tmp_274 = stq_30_bits_uop_lrs3;
      default:
        casez_tmp_274 = stq_31_bits_uop_lrs3;
    endcase
  end // always @(*)
  reg         casez_tmp_275;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_275 = stq_0_bits_uop_ldst_val;
      5'b00001:
        casez_tmp_275 = stq_1_bits_uop_ldst_val;
      5'b00010:
        casez_tmp_275 = stq_2_bits_uop_ldst_val;
      5'b00011:
        casez_tmp_275 = stq_3_bits_uop_ldst_val;
      5'b00100:
        casez_tmp_275 = stq_4_bits_uop_ldst_val;
      5'b00101:
        casez_tmp_275 = stq_5_bits_uop_ldst_val;
      5'b00110:
        casez_tmp_275 = stq_6_bits_uop_ldst_val;
      5'b00111:
        casez_tmp_275 = stq_7_bits_uop_ldst_val;
      5'b01000:
        casez_tmp_275 = stq_8_bits_uop_ldst_val;
      5'b01001:
        casez_tmp_275 = stq_9_bits_uop_ldst_val;
      5'b01010:
        casez_tmp_275 = stq_10_bits_uop_ldst_val;
      5'b01011:
        casez_tmp_275 = stq_11_bits_uop_ldst_val;
      5'b01100:
        casez_tmp_275 = stq_12_bits_uop_ldst_val;
      5'b01101:
        casez_tmp_275 = stq_13_bits_uop_ldst_val;
      5'b01110:
        casez_tmp_275 = stq_14_bits_uop_ldst_val;
      5'b01111:
        casez_tmp_275 = stq_15_bits_uop_ldst_val;
      5'b10000:
        casez_tmp_275 = stq_16_bits_uop_ldst_val;
      5'b10001:
        casez_tmp_275 = stq_17_bits_uop_ldst_val;
      5'b10010:
        casez_tmp_275 = stq_18_bits_uop_ldst_val;
      5'b10011:
        casez_tmp_275 = stq_19_bits_uop_ldst_val;
      5'b10100:
        casez_tmp_275 = stq_20_bits_uop_ldst_val;
      5'b10101:
        casez_tmp_275 = stq_21_bits_uop_ldst_val;
      5'b10110:
        casez_tmp_275 = stq_22_bits_uop_ldst_val;
      5'b10111:
        casez_tmp_275 = stq_23_bits_uop_ldst_val;
      5'b11000:
        casez_tmp_275 = stq_24_bits_uop_ldst_val;
      5'b11001:
        casez_tmp_275 = stq_25_bits_uop_ldst_val;
      5'b11010:
        casez_tmp_275 = stq_26_bits_uop_ldst_val;
      5'b11011:
        casez_tmp_275 = stq_27_bits_uop_ldst_val;
      5'b11100:
        casez_tmp_275 = stq_28_bits_uop_ldst_val;
      5'b11101:
        casez_tmp_275 = stq_29_bits_uop_ldst_val;
      5'b11110:
        casez_tmp_275 = stq_30_bits_uop_ldst_val;
      default:
        casez_tmp_275 = stq_31_bits_uop_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_276;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_276 = stq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_276 = stq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_276 = stq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_276 = stq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_276 = stq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_276 = stq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_276 = stq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_276 = stq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_276 = stq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_276 = stq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_276 = stq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_276 = stq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_276 = stq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_276 = stq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_276 = stq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_276 = stq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_276 = stq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_276 = stq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_276 = stq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_276 = stq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_276 = stq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_276 = stq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_276 = stq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_276 = stq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_276 = stq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_276 = stq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_276 = stq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_276 = stq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_276 = stq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_276 = stq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_276 = stq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_276 = stq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_277;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_277 = stq_0_bits_uop_lrs1_rtype;
      5'b00001:
        casez_tmp_277 = stq_1_bits_uop_lrs1_rtype;
      5'b00010:
        casez_tmp_277 = stq_2_bits_uop_lrs1_rtype;
      5'b00011:
        casez_tmp_277 = stq_3_bits_uop_lrs1_rtype;
      5'b00100:
        casez_tmp_277 = stq_4_bits_uop_lrs1_rtype;
      5'b00101:
        casez_tmp_277 = stq_5_bits_uop_lrs1_rtype;
      5'b00110:
        casez_tmp_277 = stq_6_bits_uop_lrs1_rtype;
      5'b00111:
        casez_tmp_277 = stq_7_bits_uop_lrs1_rtype;
      5'b01000:
        casez_tmp_277 = stq_8_bits_uop_lrs1_rtype;
      5'b01001:
        casez_tmp_277 = stq_9_bits_uop_lrs1_rtype;
      5'b01010:
        casez_tmp_277 = stq_10_bits_uop_lrs1_rtype;
      5'b01011:
        casez_tmp_277 = stq_11_bits_uop_lrs1_rtype;
      5'b01100:
        casez_tmp_277 = stq_12_bits_uop_lrs1_rtype;
      5'b01101:
        casez_tmp_277 = stq_13_bits_uop_lrs1_rtype;
      5'b01110:
        casez_tmp_277 = stq_14_bits_uop_lrs1_rtype;
      5'b01111:
        casez_tmp_277 = stq_15_bits_uop_lrs1_rtype;
      5'b10000:
        casez_tmp_277 = stq_16_bits_uop_lrs1_rtype;
      5'b10001:
        casez_tmp_277 = stq_17_bits_uop_lrs1_rtype;
      5'b10010:
        casez_tmp_277 = stq_18_bits_uop_lrs1_rtype;
      5'b10011:
        casez_tmp_277 = stq_19_bits_uop_lrs1_rtype;
      5'b10100:
        casez_tmp_277 = stq_20_bits_uop_lrs1_rtype;
      5'b10101:
        casez_tmp_277 = stq_21_bits_uop_lrs1_rtype;
      5'b10110:
        casez_tmp_277 = stq_22_bits_uop_lrs1_rtype;
      5'b10111:
        casez_tmp_277 = stq_23_bits_uop_lrs1_rtype;
      5'b11000:
        casez_tmp_277 = stq_24_bits_uop_lrs1_rtype;
      5'b11001:
        casez_tmp_277 = stq_25_bits_uop_lrs1_rtype;
      5'b11010:
        casez_tmp_277 = stq_26_bits_uop_lrs1_rtype;
      5'b11011:
        casez_tmp_277 = stq_27_bits_uop_lrs1_rtype;
      5'b11100:
        casez_tmp_277 = stq_28_bits_uop_lrs1_rtype;
      5'b11101:
        casez_tmp_277 = stq_29_bits_uop_lrs1_rtype;
      5'b11110:
        casez_tmp_277 = stq_30_bits_uop_lrs1_rtype;
      default:
        casez_tmp_277 = stq_31_bits_uop_lrs1_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_278;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_278 = stq_0_bits_uop_lrs2_rtype;
      5'b00001:
        casez_tmp_278 = stq_1_bits_uop_lrs2_rtype;
      5'b00010:
        casez_tmp_278 = stq_2_bits_uop_lrs2_rtype;
      5'b00011:
        casez_tmp_278 = stq_3_bits_uop_lrs2_rtype;
      5'b00100:
        casez_tmp_278 = stq_4_bits_uop_lrs2_rtype;
      5'b00101:
        casez_tmp_278 = stq_5_bits_uop_lrs2_rtype;
      5'b00110:
        casez_tmp_278 = stq_6_bits_uop_lrs2_rtype;
      5'b00111:
        casez_tmp_278 = stq_7_bits_uop_lrs2_rtype;
      5'b01000:
        casez_tmp_278 = stq_8_bits_uop_lrs2_rtype;
      5'b01001:
        casez_tmp_278 = stq_9_bits_uop_lrs2_rtype;
      5'b01010:
        casez_tmp_278 = stq_10_bits_uop_lrs2_rtype;
      5'b01011:
        casez_tmp_278 = stq_11_bits_uop_lrs2_rtype;
      5'b01100:
        casez_tmp_278 = stq_12_bits_uop_lrs2_rtype;
      5'b01101:
        casez_tmp_278 = stq_13_bits_uop_lrs2_rtype;
      5'b01110:
        casez_tmp_278 = stq_14_bits_uop_lrs2_rtype;
      5'b01111:
        casez_tmp_278 = stq_15_bits_uop_lrs2_rtype;
      5'b10000:
        casez_tmp_278 = stq_16_bits_uop_lrs2_rtype;
      5'b10001:
        casez_tmp_278 = stq_17_bits_uop_lrs2_rtype;
      5'b10010:
        casez_tmp_278 = stq_18_bits_uop_lrs2_rtype;
      5'b10011:
        casez_tmp_278 = stq_19_bits_uop_lrs2_rtype;
      5'b10100:
        casez_tmp_278 = stq_20_bits_uop_lrs2_rtype;
      5'b10101:
        casez_tmp_278 = stq_21_bits_uop_lrs2_rtype;
      5'b10110:
        casez_tmp_278 = stq_22_bits_uop_lrs2_rtype;
      5'b10111:
        casez_tmp_278 = stq_23_bits_uop_lrs2_rtype;
      5'b11000:
        casez_tmp_278 = stq_24_bits_uop_lrs2_rtype;
      5'b11001:
        casez_tmp_278 = stq_25_bits_uop_lrs2_rtype;
      5'b11010:
        casez_tmp_278 = stq_26_bits_uop_lrs2_rtype;
      5'b11011:
        casez_tmp_278 = stq_27_bits_uop_lrs2_rtype;
      5'b11100:
        casez_tmp_278 = stq_28_bits_uop_lrs2_rtype;
      5'b11101:
        casez_tmp_278 = stq_29_bits_uop_lrs2_rtype;
      5'b11110:
        casez_tmp_278 = stq_30_bits_uop_lrs2_rtype;
      default:
        casez_tmp_278 = stq_31_bits_uop_lrs2_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_279;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_279 = stq_0_bits_uop_frs3_en;
      5'b00001:
        casez_tmp_279 = stq_1_bits_uop_frs3_en;
      5'b00010:
        casez_tmp_279 = stq_2_bits_uop_frs3_en;
      5'b00011:
        casez_tmp_279 = stq_3_bits_uop_frs3_en;
      5'b00100:
        casez_tmp_279 = stq_4_bits_uop_frs3_en;
      5'b00101:
        casez_tmp_279 = stq_5_bits_uop_frs3_en;
      5'b00110:
        casez_tmp_279 = stq_6_bits_uop_frs3_en;
      5'b00111:
        casez_tmp_279 = stq_7_bits_uop_frs3_en;
      5'b01000:
        casez_tmp_279 = stq_8_bits_uop_frs3_en;
      5'b01001:
        casez_tmp_279 = stq_9_bits_uop_frs3_en;
      5'b01010:
        casez_tmp_279 = stq_10_bits_uop_frs3_en;
      5'b01011:
        casez_tmp_279 = stq_11_bits_uop_frs3_en;
      5'b01100:
        casez_tmp_279 = stq_12_bits_uop_frs3_en;
      5'b01101:
        casez_tmp_279 = stq_13_bits_uop_frs3_en;
      5'b01110:
        casez_tmp_279 = stq_14_bits_uop_frs3_en;
      5'b01111:
        casez_tmp_279 = stq_15_bits_uop_frs3_en;
      5'b10000:
        casez_tmp_279 = stq_16_bits_uop_frs3_en;
      5'b10001:
        casez_tmp_279 = stq_17_bits_uop_frs3_en;
      5'b10010:
        casez_tmp_279 = stq_18_bits_uop_frs3_en;
      5'b10011:
        casez_tmp_279 = stq_19_bits_uop_frs3_en;
      5'b10100:
        casez_tmp_279 = stq_20_bits_uop_frs3_en;
      5'b10101:
        casez_tmp_279 = stq_21_bits_uop_frs3_en;
      5'b10110:
        casez_tmp_279 = stq_22_bits_uop_frs3_en;
      5'b10111:
        casez_tmp_279 = stq_23_bits_uop_frs3_en;
      5'b11000:
        casez_tmp_279 = stq_24_bits_uop_frs3_en;
      5'b11001:
        casez_tmp_279 = stq_25_bits_uop_frs3_en;
      5'b11010:
        casez_tmp_279 = stq_26_bits_uop_frs3_en;
      5'b11011:
        casez_tmp_279 = stq_27_bits_uop_frs3_en;
      5'b11100:
        casez_tmp_279 = stq_28_bits_uop_frs3_en;
      5'b11101:
        casez_tmp_279 = stq_29_bits_uop_frs3_en;
      5'b11110:
        casez_tmp_279 = stq_30_bits_uop_frs3_en;
      default:
        casez_tmp_279 = stq_31_bits_uop_frs3_en;
    endcase
  end // always @(*)
  reg         casez_tmp_280;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_280 = stq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_280 = stq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_280 = stq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_280 = stq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_280 = stq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_280 = stq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_280 = stq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_280 = stq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_280 = stq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_280 = stq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_280 = stq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_280 = stq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_280 = stq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_280 = stq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_280 = stq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_280 = stq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_280 = stq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_280 = stq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_280 = stq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_280 = stq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_280 = stq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_280 = stq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_280 = stq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_280 = stq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_280 = stq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_280 = stq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_280 = stq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_280 = stq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_280 = stq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_280 = stq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_280 = stq_30_bits_uop_fp_val;
      default:
        casez_tmp_280 = stq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  reg         casez_tmp_281;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_281 = stq_0_bits_uop_fp_single;
      5'b00001:
        casez_tmp_281 = stq_1_bits_uop_fp_single;
      5'b00010:
        casez_tmp_281 = stq_2_bits_uop_fp_single;
      5'b00011:
        casez_tmp_281 = stq_3_bits_uop_fp_single;
      5'b00100:
        casez_tmp_281 = stq_4_bits_uop_fp_single;
      5'b00101:
        casez_tmp_281 = stq_5_bits_uop_fp_single;
      5'b00110:
        casez_tmp_281 = stq_6_bits_uop_fp_single;
      5'b00111:
        casez_tmp_281 = stq_7_bits_uop_fp_single;
      5'b01000:
        casez_tmp_281 = stq_8_bits_uop_fp_single;
      5'b01001:
        casez_tmp_281 = stq_9_bits_uop_fp_single;
      5'b01010:
        casez_tmp_281 = stq_10_bits_uop_fp_single;
      5'b01011:
        casez_tmp_281 = stq_11_bits_uop_fp_single;
      5'b01100:
        casez_tmp_281 = stq_12_bits_uop_fp_single;
      5'b01101:
        casez_tmp_281 = stq_13_bits_uop_fp_single;
      5'b01110:
        casez_tmp_281 = stq_14_bits_uop_fp_single;
      5'b01111:
        casez_tmp_281 = stq_15_bits_uop_fp_single;
      5'b10000:
        casez_tmp_281 = stq_16_bits_uop_fp_single;
      5'b10001:
        casez_tmp_281 = stq_17_bits_uop_fp_single;
      5'b10010:
        casez_tmp_281 = stq_18_bits_uop_fp_single;
      5'b10011:
        casez_tmp_281 = stq_19_bits_uop_fp_single;
      5'b10100:
        casez_tmp_281 = stq_20_bits_uop_fp_single;
      5'b10101:
        casez_tmp_281 = stq_21_bits_uop_fp_single;
      5'b10110:
        casez_tmp_281 = stq_22_bits_uop_fp_single;
      5'b10111:
        casez_tmp_281 = stq_23_bits_uop_fp_single;
      5'b11000:
        casez_tmp_281 = stq_24_bits_uop_fp_single;
      5'b11001:
        casez_tmp_281 = stq_25_bits_uop_fp_single;
      5'b11010:
        casez_tmp_281 = stq_26_bits_uop_fp_single;
      5'b11011:
        casez_tmp_281 = stq_27_bits_uop_fp_single;
      5'b11100:
        casez_tmp_281 = stq_28_bits_uop_fp_single;
      5'b11101:
        casez_tmp_281 = stq_29_bits_uop_fp_single;
      5'b11110:
        casez_tmp_281 = stq_30_bits_uop_fp_single;
      default:
        casez_tmp_281 = stq_31_bits_uop_fp_single;
    endcase
  end // always @(*)
  reg         casez_tmp_282;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_282 = stq_0_bits_uop_xcpt_pf_if;
      5'b00001:
        casez_tmp_282 = stq_1_bits_uop_xcpt_pf_if;
      5'b00010:
        casez_tmp_282 = stq_2_bits_uop_xcpt_pf_if;
      5'b00011:
        casez_tmp_282 = stq_3_bits_uop_xcpt_pf_if;
      5'b00100:
        casez_tmp_282 = stq_4_bits_uop_xcpt_pf_if;
      5'b00101:
        casez_tmp_282 = stq_5_bits_uop_xcpt_pf_if;
      5'b00110:
        casez_tmp_282 = stq_6_bits_uop_xcpt_pf_if;
      5'b00111:
        casez_tmp_282 = stq_7_bits_uop_xcpt_pf_if;
      5'b01000:
        casez_tmp_282 = stq_8_bits_uop_xcpt_pf_if;
      5'b01001:
        casez_tmp_282 = stq_9_bits_uop_xcpt_pf_if;
      5'b01010:
        casez_tmp_282 = stq_10_bits_uop_xcpt_pf_if;
      5'b01011:
        casez_tmp_282 = stq_11_bits_uop_xcpt_pf_if;
      5'b01100:
        casez_tmp_282 = stq_12_bits_uop_xcpt_pf_if;
      5'b01101:
        casez_tmp_282 = stq_13_bits_uop_xcpt_pf_if;
      5'b01110:
        casez_tmp_282 = stq_14_bits_uop_xcpt_pf_if;
      5'b01111:
        casez_tmp_282 = stq_15_bits_uop_xcpt_pf_if;
      5'b10000:
        casez_tmp_282 = stq_16_bits_uop_xcpt_pf_if;
      5'b10001:
        casez_tmp_282 = stq_17_bits_uop_xcpt_pf_if;
      5'b10010:
        casez_tmp_282 = stq_18_bits_uop_xcpt_pf_if;
      5'b10011:
        casez_tmp_282 = stq_19_bits_uop_xcpt_pf_if;
      5'b10100:
        casez_tmp_282 = stq_20_bits_uop_xcpt_pf_if;
      5'b10101:
        casez_tmp_282 = stq_21_bits_uop_xcpt_pf_if;
      5'b10110:
        casez_tmp_282 = stq_22_bits_uop_xcpt_pf_if;
      5'b10111:
        casez_tmp_282 = stq_23_bits_uop_xcpt_pf_if;
      5'b11000:
        casez_tmp_282 = stq_24_bits_uop_xcpt_pf_if;
      5'b11001:
        casez_tmp_282 = stq_25_bits_uop_xcpt_pf_if;
      5'b11010:
        casez_tmp_282 = stq_26_bits_uop_xcpt_pf_if;
      5'b11011:
        casez_tmp_282 = stq_27_bits_uop_xcpt_pf_if;
      5'b11100:
        casez_tmp_282 = stq_28_bits_uop_xcpt_pf_if;
      5'b11101:
        casez_tmp_282 = stq_29_bits_uop_xcpt_pf_if;
      5'b11110:
        casez_tmp_282 = stq_30_bits_uop_xcpt_pf_if;
      default:
        casez_tmp_282 = stq_31_bits_uop_xcpt_pf_if;
    endcase
  end // always @(*)
  reg         casez_tmp_283;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_283 = stq_0_bits_uop_xcpt_ae_if;
      5'b00001:
        casez_tmp_283 = stq_1_bits_uop_xcpt_ae_if;
      5'b00010:
        casez_tmp_283 = stq_2_bits_uop_xcpt_ae_if;
      5'b00011:
        casez_tmp_283 = stq_3_bits_uop_xcpt_ae_if;
      5'b00100:
        casez_tmp_283 = stq_4_bits_uop_xcpt_ae_if;
      5'b00101:
        casez_tmp_283 = stq_5_bits_uop_xcpt_ae_if;
      5'b00110:
        casez_tmp_283 = stq_6_bits_uop_xcpt_ae_if;
      5'b00111:
        casez_tmp_283 = stq_7_bits_uop_xcpt_ae_if;
      5'b01000:
        casez_tmp_283 = stq_8_bits_uop_xcpt_ae_if;
      5'b01001:
        casez_tmp_283 = stq_9_bits_uop_xcpt_ae_if;
      5'b01010:
        casez_tmp_283 = stq_10_bits_uop_xcpt_ae_if;
      5'b01011:
        casez_tmp_283 = stq_11_bits_uop_xcpt_ae_if;
      5'b01100:
        casez_tmp_283 = stq_12_bits_uop_xcpt_ae_if;
      5'b01101:
        casez_tmp_283 = stq_13_bits_uop_xcpt_ae_if;
      5'b01110:
        casez_tmp_283 = stq_14_bits_uop_xcpt_ae_if;
      5'b01111:
        casez_tmp_283 = stq_15_bits_uop_xcpt_ae_if;
      5'b10000:
        casez_tmp_283 = stq_16_bits_uop_xcpt_ae_if;
      5'b10001:
        casez_tmp_283 = stq_17_bits_uop_xcpt_ae_if;
      5'b10010:
        casez_tmp_283 = stq_18_bits_uop_xcpt_ae_if;
      5'b10011:
        casez_tmp_283 = stq_19_bits_uop_xcpt_ae_if;
      5'b10100:
        casez_tmp_283 = stq_20_bits_uop_xcpt_ae_if;
      5'b10101:
        casez_tmp_283 = stq_21_bits_uop_xcpt_ae_if;
      5'b10110:
        casez_tmp_283 = stq_22_bits_uop_xcpt_ae_if;
      5'b10111:
        casez_tmp_283 = stq_23_bits_uop_xcpt_ae_if;
      5'b11000:
        casez_tmp_283 = stq_24_bits_uop_xcpt_ae_if;
      5'b11001:
        casez_tmp_283 = stq_25_bits_uop_xcpt_ae_if;
      5'b11010:
        casez_tmp_283 = stq_26_bits_uop_xcpt_ae_if;
      5'b11011:
        casez_tmp_283 = stq_27_bits_uop_xcpt_ae_if;
      5'b11100:
        casez_tmp_283 = stq_28_bits_uop_xcpt_ae_if;
      5'b11101:
        casez_tmp_283 = stq_29_bits_uop_xcpt_ae_if;
      5'b11110:
        casez_tmp_283 = stq_30_bits_uop_xcpt_ae_if;
      default:
        casez_tmp_283 = stq_31_bits_uop_xcpt_ae_if;
    endcase
  end // always @(*)
  reg         casez_tmp_284;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_284 = stq_0_bits_uop_xcpt_ma_if;
      5'b00001:
        casez_tmp_284 = stq_1_bits_uop_xcpt_ma_if;
      5'b00010:
        casez_tmp_284 = stq_2_bits_uop_xcpt_ma_if;
      5'b00011:
        casez_tmp_284 = stq_3_bits_uop_xcpt_ma_if;
      5'b00100:
        casez_tmp_284 = stq_4_bits_uop_xcpt_ma_if;
      5'b00101:
        casez_tmp_284 = stq_5_bits_uop_xcpt_ma_if;
      5'b00110:
        casez_tmp_284 = stq_6_bits_uop_xcpt_ma_if;
      5'b00111:
        casez_tmp_284 = stq_7_bits_uop_xcpt_ma_if;
      5'b01000:
        casez_tmp_284 = stq_8_bits_uop_xcpt_ma_if;
      5'b01001:
        casez_tmp_284 = stq_9_bits_uop_xcpt_ma_if;
      5'b01010:
        casez_tmp_284 = stq_10_bits_uop_xcpt_ma_if;
      5'b01011:
        casez_tmp_284 = stq_11_bits_uop_xcpt_ma_if;
      5'b01100:
        casez_tmp_284 = stq_12_bits_uop_xcpt_ma_if;
      5'b01101:
        casez_tmp_284 = stq_13_bits_uop_xcpt_ma_if;
      5'b01110:
        casez_tmp_284 = stq_14_bits_uop_xcpt_ma_if;
      5'b01111:
        casez_tmp_284 = stq_15_bits_uop_xcpt_ma_if;
      5'b10000:
        casez_tmp_284 = stq_16_bits_uop_xcpt_ma_if;
      5'b10001:
        casez_tmp_284 = stq_17_bits_uop_xcpt_ma_if;
      5'b10010:
        casez_tmp_284 = stq_18_bits_uop_xcpt_ma_if;
      5'b10011:
        casez_tmp_284 = stq_19_bits_uop_xcpt_ma_if;
      5'b10100:
        casez_tmp_284 = stq_20_bits_uop_xcpt_ma_if;
      5'b10101:
        casez_tmp_284 = stq_21_bits_uop_xcpt_ma_if;
      5'b10110:
        casez_tmp_284 = stq_22_bits_uop_xcpt_ma_if;
      5'b10111:
        casez_tmp_284 = stq_23_bits_uop_xcpt_ma_if;
      5'b11000:
        casez_tmp_284 = stq_24_bits_uop_xcpt_ma_if;
      5'b11001:
        casez_tmp_284 = stq_25_bits_uop_xcpt_ma_if;
      5'b11010:
        casez_tmp_284 = stq_26_bits_uop_xcpt_ma_if;
      5'b11011:
        casez_tmp_284 = stq_27_bits_uop_xcpt_ma_if;
      5'b11100:
        casez_tmp_284 = stq_28_bits_uop_xcpt_ma_if;
      5'b11101:
        casez_tmp_284 = stq_29_bits_uop_xcpt_ma_if;
      5'b11110:
        casez_tmp_284 = stq_30_bits_uop_xcpt_ma_if;
      default:
        casez_tmp_284 = stq_31_bits_uop_xcpt_ma_if;
    endcase
  end // always @(*)
  reg         casez_tmp_285;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_285 = stq_0_bits_uop_bp_debug_if;
      5'b00001:
        casez_tmp_285 = stq_1_bits_uop_bp_debug_if;
      5'b00010:
        casez_tmp_285 = stq_2_bits_uop_bp_debug_if;
      5'b00011:
        casez_tmp_285 = stq_3_bits_uop_bp_debug_if;
      5'b00100:
        casez_tmp_285 = stq_4_bits_uop_bp_debug_if;
      5'b00101:
        casez_tmp_285 = stq_5_bits_uop_bp_debug_if;
      5'b00110:
        casez_tmp_285 = stq_6_bits_uop_bp_debug_if;
      5'b00111:
        casez_tmp_285 = stq_7_bits_uop_bp_debug_if;
      5'b01000:
        casez_tmp_285 = stq_8_bits_uop_bp_debug_if;
      5'b01001:
        casez_tmp_285 = stq_9_bits_uop_bp_debug_if;
      5'b01010:
        casez_tmp_285 = stq_10_bits_uop_bp_debug_if;
      5'b01011:
        casez_tmp_285 = stq_11_bits_uop_bp_debug_if;
      5'b01100:
        casez_tmp_285 = stq_12_bits_uop_bp_debug_if;
      5'b01101:
        casez_tmp_285 = stq_13_bits_uop_bp_debug_if;
      5'b01110:
        casez_tmp_285 = stq_14_bits_uop_bp_debug_if;
      5'b01111:
        casez_tmp_285 = stq_15_bits_uop_bp_debug_if;
      5'b10000:
        casez_tmp_285 = stq_16_bits_uop_bp_debug_if;
      5'b10001:
        casez_tmp_285 = stq_17_bits_uop_bp_debug_if;
      5'b10010:
        casez_tmp_285 = stq_18_bits_uop_bp_debug_if;
      5'b10011:
        casez_tmp_285 = stq_19_bits_uop_bp_debug_if;
      5'b10100:
        casez_tmp_285 = stq_20_bits_uop_bp_debug_if;
      5'b10101:
        casez_tmp_285 = stq_21_bits_uop_bp_debug_if;
      5'b10110:
        casez_tmp_285 = stq_22_bits_uop_bp_debug_if;
      5'b10111:
        casez_tmp_285 = stq_23_bits_uop_bp_debug_if;
      5'b11000:
        casez_tmp_285 = stq_24_bits_uop_bp_debug_if;
      5'b11001:
        casez_tmp_285 = stq_25_bits_uop_bp_debug_if;
      5'b11010:
        casez_tmp_285 = stq_26_bits_uop_bp_debug_if;
      5'b11011:
        casez_tmp_285 = stq_27_bits_uop_bp_debug_if;
      5'b11100:
        casez_tmp_285 = stq_28_bits_uop_bp_debug_if;
      5'b11101:
        casez_tmp_285 = stq_29_bits_uop_bp_debug_if;
      5'b11110:
        casez_tmp_285 = stq_30_bits_uop_bp_debug_if;
      default:
        casez_tmp_285 = stq_31_bits_uop_bp_debug_if;
    endcase
  end // always @(*)
  reg         casez_tmp_286;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_286 = stq_0_bits_uop_bp_xcpt_if;
      5'b00001:
        casez_tmp_286 = stq_1_bits_uop_bp_xcpt_if;
      5'b00010:
        casez_tmp_286 = stq_2_bits_uop_bp_xcpt_if;
      5'b00011:
        casez_tmp_286 = stq_3_bits_uop_bp_xcpt_if;
      5'b00100:
        casez_tmp_286 = stq_4_bits_uop_bp_xcpt_if;
      5'b00101:
        casez_tmp_286 = stq_5_bits_uop_bp_xcpt_if;
      5'b00110:
        casez_tmp_286 = stq_6_bits_uop_bp_xcpt_if;
      5'b00111:
        casez_tmp_286 = stq_7_bits_uop_bp_xcpt_if;
      5'b01000:
        casez_tmp_286 = stq_8_bits_uop_bp_xcpt_if;
      5'b01001:
        casez_tmp_286 = stq_9_bits_uop_bp_xcpt_if;
      5'b01010:
        casez_tmp_286 = stq_10_bits_uop_bp_xcpt_if;
      5'b01011:
        casez_tmp_286 = stq_11_bits_uop_bp_xcpt_if;
      5'b01100:
        casez_tmp_286 = stq_12_bits_uop_bp_xcpt_if;
      5'b01101:
        casez_tmp_286 = stq_13_bits_uop_bp_xcpt_if;
      5'b01110:
        casez_tmp_286 = stq_14_bits_uop_bp_xcpt_if;
      5'b01111:
        casez_tmp_286 = stq_15_bits_uop_bp_xcpt_if;
      5'b10000:
        casez_tmp_286 = stq_16_bits_uop_bp_xcpt_if;
      5'b10001:
        casez_tmp_286 = stq_17_bits_uop_bp_xcpt_if;
      5'b10010:
        casez_tmp_286 = stq_18_bits_uop_bp_xcpt_if;
      5'b10011:
        casez_tmp_286 = stq_19_bits_uop_bp_xcpt_if;
      5'b10100:
        casez_tmp_286 = stq_20_bits_uop_bp_xcpt_if;
      5'b10101:
        casez_tmp_286 = stq_21_bits_uop_bp_xcpt_if;
      5'b10110:
        casez_tmp_286 = stq_22_bits_uop_bp_xcpt_if;
      5'b10111:
        casez_tmp_286 = stq_23_bits_uop_bp_xcpt_if;
      5'b11000:
        casez_tmp_286 = stq_24_bits_uop_bp_xcpt_if;
      5'b11001:
        casez_tmp_286 = stq_25_bits_uop_bp_xcpt_if;
      5'b11010:
        casez_tmp_286 = stq_26_bits_uop_bp_xcpt_if;
      5'b11011:
        casez_tmp_286 = stq_27_bits_uop_bp_xcpt_if;
      5'b11100:
        casez_tmp_286 = stq_28_bits_uop_bp_xcpt_if;
      5'b11101:
        casez_tmp_286 = stq_29_bits_uop_bp_xcpt_if;
      5'b11110:
        casez_tmp_286 = stq_30_bits_uop_bp_xcpt_if;
      default:
        casez_tmp_286 = stq_31_bits_uop_bp_xcpt_if;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_287;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_287 = stq_0_bits_uop_debug_fsrc;
      5'b00001:
        casez_tmp_287 = stq_1_bits_uop_debug_fsrc;
      5'b00010:
        casez_tmp_287 = stq_2_bits_uop_debug_fsrc;
      5'b00011:
        casez_tmp_287 = stq_3_bits_uop_debug_fsrc;
      5'b00100:
        casez_tmp_287 = stq_4_bits_uop_debug_fsrc;
      5'b00101:
        casez_tmp_287 = stq_5_bits_uop_debug_fsrc;
      5'b00110:
        casez_tmp_287 = stq_6_bits_uop_debug_fsrc;
      5'b00111:
        casez_tmp_287 = stq_7_bits_uop_debug_fsrc;
      5'b01000:
        casez_tmp_287 = stq_8_bits_uop_debug_fsrc;
      5'b01001:
        casez_tmp_287 = stq_9_bits_uop_debug_fsrc;
      5'b01010:
        casez_tmp_287 = stq_10_bits_uop_debug_fsrc;
      5'b01011:
        casez_tmp_287 = stq_11_bits_uop_debug_fsrc;
      5'b01100:
        casez_tmp_287 = stq_12_bits_uop_debug_fsrc;
      5'b01101:
        casez_tmp_287 = stq_13_bits_uop_debug_fsrc;
      5'b01110:
        casez_tmp_287 = stq_14_bits_uop_debug_fsrc;
      5'b01111:
        casez_tmp_287 = stq_15_bits_uop_debug_fsrc;
      5'b10000:
        casez_tmp_287 = stq_16_bits_uop_debug_fsrc;
      5'b10001:
        casez_tmp_287 = stq_17_bits_uop_debug_fsrc;
      5'b10010:
        casez_tmp_287 = stq_18_bits_uop_debug_fsrc;
      5'b10011:
        casez_tmp_287 = stq_19_bits_uop_debug_fsrc;
      5'b10100:
        casez_tmp_287 = stq_20_bits_uop_debug_fsrc;
      5'b10101:
        casez_tmp_287 = stq_21_bits_uop_debug_fsrc;
      5'b10110:
        casez_tmp_287 = stq_22_bits_uop_debug_fsrc;
      5'b10111:
        casez_tmp_287 = stq_23_bits_uop_debug_fsrc;
      5'b11000:
        casez_tmp_287 = stq_24_bits_uop_debug_fsrc;
      5'b11001:
        casez_tmp_287 = stq_25_bits_uop_debug_fsrc;
      5'b11010:
        casez_tmp_287 = stq_26_bits_uop_debug_fsrc;
      5'b11011:
        casez_tmp_287 = stq_27_bits_uop_debug_fsrc;
      5'b11100:
        casez_tmp_287 = stq_28_bits_uop_debug_fsrc;
      5'b11101:
        casez_tmp_287 = stq_29_bits_uop_debug_fsrc;
      5'b11110:
        casez_tmp_287 = stq_30_bits_uop_debug_fsrc;
      default:
        casez_tmp_287 = stq_31_bits_uop_debug_fsrc;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_288;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_288 = stq_0_bits_uop_debug_tsrc;
      5'b00001:
        casez_tmp_288 = stq_1_bits_uop_debug_tsrc;
      5'b00010:
        casez_tmp_288 = stq_2_bits_uop_debug_tsrc;
      5'b00011:
        casez_tmp_288 = stq_3_bits_uop_debug_tsrc;
      5'b00100:
        casez_tmp_288 = stq_4_bits_uop_debug_tsrc;
      5'b00101:
        casez_tmp_288 = stq_5_bits_uop_debug_tsrc;
      5'b00110:
        casez_tmp_288 = stq_6_bits_uop_debug_tsrc;
      5'b00111:
        casez_tmp_288 = stq_7_bits_uop_debug_tsrc;
      5'b01000:
        casez_tmp_288 = stq_8_bits_uop_debug_tsrc;
      5'b01001:
        casez_tmp_288 = stq_9_bits_uop_debug_tsrc;
      5'b01010:
        casez_tmp_288 = stq_10_bits_uop_debug_tsrc;
      5'b01011:
        casez_tmp_288 = stq_11_bits_uop_debug_tsrc;
      5'b01100:
        casez_tmp_288 = stq_12_bits_uop_debug_tsrc;
      5'b01101:
        casez_tmp_288 = stq_13_bits_uop_debug_tsrc;
      5'b01110:
        casez_tmp_288 = stq_14_bits_uop_debug_tsrc;
      5'b01111:
        casez_tmp_288 = stq_15_bits_uop_debug_tsrc;
      5'b10000:
        casez_tmp_288 = stq_16_bits_uop_debug_tsrc;
      5'b10001:
        casez_tmp_288 = stq_17_bits_uop_debug_tsrc;
      5'b10010:
        casez_tmp_288 = stq_18_bits_uop_debug_tsrc;
      5'b10011:
        casez_tmp_288 = stq_19_bits_uop_debug_tsrc;
      5'b10100:
        casez_tmp_288 = stq_20_bits_uop_debug_tsrc;
      5'b10101:
        casez_tmp_288 = stq_21_bits_uop_debug_tsrc;
      5'b10110:
        casez_tmp_288 = stq_22_bits_uop_debug_tsrc;
      5'b10111:
        casez_tmp_288 = stq_23_bits_uop_debug_tsrc;
      5'b11000:
        casez_tmp_288 = stq_24_bits_uop_debug_tsrc;
      5'b11001:
        casez_tmp_288 = stq_25_bits_uop_debug_tsrc;
      5'b11010:
        casez_tmp_288 = stq_26_bits_uop_debug_tsrc;
      5'b11011:
        casez_tmp_288 = stq_27_bits_uop_debug_tsrc;
      5'b11100:
        casez_tmp_288 = stq_28_bits_uop_debug_tsrc;
      5'b11101:
        casez_tmp_288 = stq_29_bits_uop_debug_tsrc;
      5'b11110:
        casez_tmp_288 = stq_30_bits_uop_debug_tsrc;
      default:
        casez_tmp_288 = stq_31_bits_uop_debug_tsrc;
    endcase
  end // always @(*)
  reg         casez_tmp_289;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_289 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_289 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_289 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_289 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_289 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_289 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_289 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_289 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_289 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_289 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_289 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_289 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_289 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_289 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_289 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_289 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_289 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_289 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_289 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_289 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_289 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_289 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_289 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_289 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_289 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_289 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_289 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_289 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_289 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_289 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_289 = stq_30_bits_addr_valid;
      default:
        casez_tmp_289 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_290;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_290 = stq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_290 = stq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_290 = stq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_290 = stq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_290 = stq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_290 = stq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_290 = stq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_290 = stq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_290 = stq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_290 = stq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_290 = stq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_290 = stq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_290 = stq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_290 = stq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_290 = stq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_290 = stq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_290 = stq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_290 = stq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_290 = stq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_290 = stq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_290 = stq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_290 = stq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_290 = stq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_290 = stq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_290 = stq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_290 = stq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_290 = stq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_290 = stq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_290 = stq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_290 = stq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_290 = stq_30_bits_addr_bits;
      default:
        casez_tmp_290 = stq_31_bits_addr_bits;
    endcase
  end // always @(*)
  reg         casez_tmp_291;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_291 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_291 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_291 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_291 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_291 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_291 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_291 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_291 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_291 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_291 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_291 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_291 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_291 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_291 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_291 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_291 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_291 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_291 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_291 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_291 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_291 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_291 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_291 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_291 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_291 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_291 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_291 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_291 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_291 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_291 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_291 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_291 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         casez_tmp_292;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_292 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_292 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_292 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_292 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_292 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_292 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_292 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_292 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_292 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_292 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_292 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_292 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_292 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_292 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_292 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_292 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_292 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_292 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_292 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_292 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_292 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_292 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_292 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_292 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_292 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_292 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_292 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_292 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_292 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_292 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_292 = stq_30_bits_data_valid;
      default:
        casez_tmp_292 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg         can_fire_sta_retry_REG_1;
  reg         casez_tmp_293;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_293 = ldq_0_valid;
      5'b00001:
        casez_tmp_293 = ldq_1_valid;
      5'b00010:
        casez_tmp_293 = ldq_2_valid;
      5'b00011:
        casez_tmp_293 = ldq_3_valid;
      5'b00100:
        casez_tmp_293 = ldq_4_valid;
      5'b00101:
        casez_tmp_293 = ldq_5_valid;
      5'b00110:
        casez_tmp_293 = ldq_6_valid;
      5'b00111:
        casez_tmp_293 = ldq_7_valid;
      5'b01000:
        casez_tmp_293 = ldq_8_valid;
      5'b01001:
        casez_tmp_293 = ldq_9_valid;
      5'b01010:
        casez_tmp_293 = ldq_10_valid;
      5'b01011:
        casez_tmp_293 = ldq_11_valid;
      5'b01100:
        casez_tmp_293 = ldq_12_valid;
      5'b01101:
        casez_tmp_293 = ldq_13_valid;
      5'b01110:
        casez_tmp_293 = ldq_14_valid;
      5'b01111:
        casez_tmp_293 = ldq_15_valid;
      5'b10000:
        casez_tmp_293 = ldq_16_valid;
      5'b10001:
        casez_tmp_293 = ldq_17_valid;
      5'b10010:
        casez_tmp_293 = ldq_18_valid;
      5'b10011:
        casez_tmp_293 = ldq_19_valid;
      5'b10100:
        casez_tmp_293 = ldq_20_valid;
      5'b10101:
        casez_tmp_293 = ldq_21_valid;
      5'b10110:
        casez_tmp_293 = ldq_22_valid;
      5'b10111:
        casez_tmp_293 = ldq_23_valid;
      5'b11000:
        casez_tmp_293 = ldq_24_valid;
      5'b11001:
        casez_tmp_293 = ldq_25_valid;
      5'b11010:
        casez_tmp_293 = ldq_26_valid;
      5'b11011:
        casez_tmp_293 = ldq_27_valid;
      5'b11100:
        casez_tmp_293 = ldq_28_valid;
      5'b11101:
        casez_tmp_293 = ldq_29_valid;
      5'b11110:
        casez_tmp_293 = ldq_30_valid;
      default:
        casez_tmp_293 = ldq_31_valid;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_294;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_294 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_294 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_294 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_294 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_294 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_294 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_294 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_294 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_294 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_294 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_294 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_294 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_294 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_294 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_294 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_294 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_294 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_294 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_294 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_294 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_294 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_294 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_294 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_294 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_294 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_294 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_294 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_294 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_294 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_294 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_294 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_294 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_295;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_295 = ldq_0_bits_uop_inst;
      5'b00001:
        casez_tmp_295 = ldq_1_bits_uop_inst;
      5'b00010:
        casez_tmp_295 = ldq_2_bits_uop_inst;
      5'b00011:
        casez_tmp_295 = ldq_3_bits_uop_inst;
      5'b00100:
        casez_tmp_295 = ldq_4_bits_uop_inst;
      5'b00101:
        casez_tmp_295 = ldq_5_bits_uop_inst;
      5'b00110:
        casez_tmp_295 = ldq_6_bits_uop_inst;
      5'b00111:
        casez_tmp_295 = ldq_7_bits_uop_inst;
      5'b01000:
        casez_tmp_295 = ldq_8_bits_uop_inst;
      5'b01001:
        casez_tmp_295 = ldq_9_bits_uop_inst;
      5'b01010:
        casez_tmp_295 = ldq_10_bits_uop_inst;
      5'b01011:
        casez_tmp_295 = ldq_11_bits_uop_inst;
      5'b01100:
        casez_tmp_295 = ldq_12_bits_uop_inst;
      5'b01101:
        casez_tmp_295 = ldq_13_bits_uop_inst;
      5'b01110:
        casez_tmp_295 = ldq_14_bits_uop_inst;
      5'b01111:
        casez_tmp_295 = ldq_15_bits_uop_inst;
      5'b10000:
        casez_tmp_295 = ldq_16_bits_uop_inst;
      5'b10001:
        casez_tmp_295 = ldq_17_bits_uop_inst;
      5'b10010:
        casez_tmp_295 = ldq_18_bits_uop_inst;
      5'b10011:
        casez_tmp_295 = ldq_19_bits_uop_inst;
      5'b10100:
        casez_tmp_295 = ldq_20_bits_uop_inst;
      5'b10101:
        casez_tmp_295 = ldq_21_bits_uop_inst;
      5'b10110:
        casez_tmp_295 = ldq_22_bits_uop_inst;
      5'b10111:
        casez_tmp_295 = ldq_23_bits_uop_inst;
      5'b11000:
        casez_tmp_295 = ldq_24_bits_uop_inst;
      5'b11001:
        casez_tmp_295 = ldq_25_bits_uop_inst;
      5'b11010:
        casez_tmp_295 = ldq_26_bits_uop_inst;
      5'b11011:
        casez_tmp_295 = ldq_27_bits_uop_inst;
      5'b11100:
        casez_tmp_295 = ldq_28_bits_uop_inst;
      5'b11101:
        casez_tmp_295 = ldq_29_bits_uop_inst;
      5'b11110:
        casez_tmp_295 = ldq_30_bits_uop_inst;
      default:
        casez_tmp_295 = ldq_31_bits_uop_inst;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_296;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_296 = ldq_0_bits_uop_debug_inst;
      5'b00001:
        casez_tmp_296 = ldq_1_bits_uop_debug_inst;
      5'b00010:
        casez_tmp_296 = ldq_2_bits_uop_debug_inst;
      5'b00011:
        casez_tmp_296 = ldq_3_bits_uop_debug_inst;
      5'b00100:
        casez_tmp_296 = ldq_4_bits_uop_debug_inst;
      5'b00101:
        casez_tmp_296 = ldq_5_bits_uop_debug_inst;
      5'b00110:
        casez_tmp_296 = ldq_6_bits_uop_debug_inst;
      5'b00111:
        casez_tmp_296 = ldq_7_bits_uop_debug_inst;
      5'b01000:
        casez_tmp_296 = ldq_8_bits_uop_debug_inst;
      5'b01001:
        casez_tmp_296 = ldq_9_bits_uop_debug_inst;
      5'b01010:
        casez_tmp_296 = ldq_10_bits_uop_debug_inst;
      5'b01011:
        casez_tmp_296 = ldq_11_bits_uop_debug_inst;
      5'b01100:
        casez_tmp_296 = ldq_12_bits_uop_debug_inst;
      5'b01101:
        casez_tmp_296 = ldq_13_bits_uop_debug_inst;
      5'b01110:
        casez_tmp_296 = ldq_14_bits_uop_debug_inst;
      5'b01111:
        casez_tmp_296 = ldq_15_bits_uop_debug_inst;
      5'b10000:
        casez_tmp_296 = ldq_16_bits_uop_debug_inst;
      5'b10001:
        casez_tmp_296 = ldq_17_bits_uop_debug_inst;
      5'b10010:
        casez_tmp_296 = ldq_18_bits_uop_debug_inst;
      5'b10011:
        casez_tmp_296 = ldq_19_bits_uop_debug_inst;
      5'b10100:
        casez_tmp_296 = ldq_20_bits_uop_debug_inst;
      5'b10101:
        casez_tmp_296 = ldq_21_bits_uop_debug_inst;
      5'b10110:
        casez_tmp_296 = ldq_22_bits_uop_debug_inst;
      5'b10111:
        casez_tmp_296 = ldq_23_bits_uop_debug_inst;
      5'b11000:
        casez_tmp_296 = ldq_24_bits_uop_debug_inst;
      5'b11001:
        casez_tmp_296 = ldq_25_bits_uop_debug_inst;
      5'b11010:
        casez_tmp_296 = ldq_26_bits_uop_debug_inst;
      5'b11011:
        casez_tmp_296 = ldq_27_bits_uop_debug_inst;
      5'b11100:
        casez_tmp_296 = ldq_28_bits_uop_debug_inst;
      5'b11101:
        casez_tmp_296 = ldq_29_bits_uop_debug_inst;
      5'b11110:
        casez_tmp_296 = ldq_30_bits_uop_debug_inst;
      default:
        casez_tmp_296 = ldq_31_bits_uop_debug_inst;
    endcase
  end // always @(*)
  reg         casez_tmp_297;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_297 = ldq_0_bits_uop_is_rvc;
      5'b00001:
        casez_tmp_297 = ldq_1_bits_uop_is_rvc;
      5'b00010:
        casez_tmp_297 = ldq_2_bits_uop_is_rvc;
      5'b00011:
        casez_tmp_297 = ldq_3_bits_uop_is_rvc;
      5'b00100:
        casez_tmp_297 = ldq_4_bits_uop_is_rvc;
      5'b00101:
        casez_tmp_297 = ldq_5_bits_uop_is_rvc;
      5'b00110:
        casez_tmp_297 = ldq_6_bits_uop_is_rvc;
      5'b00111:
        casez_tmp_297 = ldq_7_bits_uop_is_rvc;
      5'b01000:
        casez_tmp_297 = ldq_8_bits_uop_is_rvc;
      5'b01001:
        casez_tmp_297 = ldq_9_bits_uop_is_rvc;
      5'b01010:
        casez_tmp_297 = ldq_10_bits_uop_is_rvc;
      5'b01011:
        casez_tmp_297 = ldq_11_bits_uop_is_rvc;
      5'b01100:
        casez_tmp_297 = ldq_12_bits_uop_is_rvc;
      5'b01101:
        casez_tmp_297 = ldq_13_bits_uop_is_rvc;
      5'b01110:
        casez_tmp_297 = ldq_14_bits_uop_is_rvc;
      5'b01111:
        casez_tmp_297 = ldq_15_bits_uop_is_rvc;
      5'b10000:
        casez_tmp_297 = ldq_16_bits_uop_is_rvc;
      5'b10001:
        casez_tmp_297 = ldq_17_bits_uop_is_rvc;
      5'b10010:
        casez_tmp_297 = ldq_18_bits_uop_is_rvc;
      5'b10011:
        casez_tmp_297 = ldq_19_bits_uop_is_rvc;
      5'b10100:
        casez_tmp_297 = ldq_20_bits_uop_is_rvc;
      5'b10101:
        casez_tmp_297 = ldq_21_bits_uop_is_rvc;
      5'b10110:
        casez_tmp_297 = ldq_22_bits_uop_is_rvc;
      5'b10111:
        casez_tmp_297 = ldq_23_bits_uop_is_rvc;
      5'b11000:
        casez_tmp_297 = ldq_24_bits_uop_is_rvc;
      5'b11001:
        casez_tmp_297 = ldq_25_bits_uop_is_rvc;
      5'b11010:
        casez_tmp_297 = ldq_26_bits_uop_is_rvc;
      5'b11011:
        casez_tmp_297 = ldq_27_bits_uop_is_rvc;
      5'b11100:
        casez_tmp_297 = ldq_28_bits_uop_is_rvc;
      5'b11101:
        casez_tmp_297 = ldq_29_bits_uop_is_rvc;
      5'b11110:
        casez_tmp_297 = ldq_30_bits_uop_is_rvc;
      default:
        casez_tmp_297 = ldq_31_bits_uop_is_rvc;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_298;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_298 = ldq_0_bits_uop_debug_pc;
      5'b00001:
        casez_tmp_298 = ldq_1_bits_uop_debug_pc;
      5'b00010:
        casez_tmp_298 = ldq_2_bits_uop_debug_pc;
      5'b00011:
        casez_tmp_298 = ldq_3_bits_uop_debug_pc;
      5'b00100:
        casez_tmp_298 = ldq_4_bits_uop_debug_pc;
      5'b00101:
        casez_tmp_298 = ldq_5_bits_uop_debug_pc;
      5'b00110:
        casez_tmp_298 = ldq_6_bits_uop_debug_pc;
      5'b00111:
        casez_tmp_298 = ldq_7_bits_uop_debug_pc;
      5'b01000:
        casez_tmp_298 = ldq_8_bits_uop_debug_pc;
      5'b01001:
        casez_tmp_298 = ldq_9_bits_uop_debug_pc;
      5'b01010:
        casez_tmp_298 = ldq_10_bits_uop_debug_pc;
      5'b01011:
        casez_tmp_298 = ldq_11_bits_uop_debug_pc;
      5'b01100:
        casez_tmp_298 = ldq_12_bits_uop_debug_pc;
      5'b01101:
        casez_tmp_298 = ldq_13_bits_uop_debug_pc;
      5'b01110:
        casez_tmp_298 = ldq_14_bits_uop_debug_pc;
      5'b01111:
        casez_tmp_298 = ldq_15_bits_uop_debug_pc;
      5'b10000:
        casez_tmp_298 = ldq_16_bits_uop_debug_pc;
      5'b10001:
        casez_tmp_298 = ldq_17_bits_uop_debug_pc;
      5'b10010:
        casez_tmp_298 = ldq_18_bits_uop_debug_pc;
      5'b10011:
        casez_tmp_298 = ldq_19_bits_uop_debug_pc;
      5'b10100:
        casez_tmp_298 = ldq_20_bits_uop_debug_pc;
      5'b10101:
        casez_tmp_298 = ldq_21_bits_uop_debug_pc;
      5'b10110:
        casez_tmp_298 = ldq_22_bits_uop_debug_pc;
      5'b10111:
        casez_tmp_298 = ldq_23_bits_uop_debug_pc;
      5'b11000:
        casez_tmp_298 = ldq_24_bits_uop_debug_pc;
      5'b11001:
        casez_tmp_298 = ldq_25_bits_uop_debug_pc;
      5'b11010:
        casez_tmp_298 = ldq_26_bits_uop_debug_pc;
      5'b11011:
        casez_tmp_298 = ldq_27_bits_uop_debug_pc;
      5'b11100:
        casez_tmp_298 = ldq_28_bits_uop_debug_pc;
      5'b11101:
        casez_tmp_298 = ldq_29_bits_uop_debug_pc;
      5'b11110:
        casez_tmp_298 = ldq_30_bits_uop_debug_pc;
      default:
        casez_tmp_298 = ldq_31_bits_uop_debug_pc;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_299;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_299 = ldq_0_bits_uop_iq_type;
      5'b00001:
        casez_tmp_299 = ldq_1_bits_uop_iq_type;
      5'b00010:
        casez_tmp_299 = ldq_2_bits_uop_iq_type;
      5'b00011:
        casez_tmp_299 = ldq_3_bits_uop_iq_type;
      5'b00100:
        casez_tmp_299 = ldq_4_bits_uop_iq_type;
      5'b00101:
        casez_tmp_299 = ldq_5_bits_uop_iq_type;
      5'b00110:
        casez_tmp_299 = ldq_6_bits_uop_iq_type;
      5'b00111:
        casez_tmp_299 = ldq_7_bits_uop_iq_type;
      5'b01000:
        casez_tmp_299 = ldq_8_bits_uop_iq_type;
      5'b01001:
        casez_tmp_299 = ldq_9_bits_uop_iq_type;
      5'b01010:
        casez_tmp_299 = ldq_10_bits_uop_iq_type;
      5'b01011:
        casez_tmp_299 = ldq_11_bits_uop_iq_type;
      5'b01100:
        casez_tmp_299 = ldq_12_bits_uop_iq_type;
      5'b01101:
        casez_tmp_299 = ldq_13_bits_uop_iq_type;
      5'b01110:
        casez_tmp_299 = ldq_14_bits_uop_iq_type;
      5'b01111:
        casez_tmp_299 = ldq_15_bits_uop_iq_type;
      5'b10000:
        casez_tmp_299 = ldq_16_bits_uop_iq_type;
      5'b10001:
        casez_tmp_299 = ldq_17_bits_uop_iq_type;
      5'b10010:
        casez_tmp_299 = ldq_18_bits_uop_iq_type;
      5'b10011:
        casez_tmp_299 = ldq_19_bits_uop_iq_type;
      5'b10100:
        casez_tmp_299 = ldq_20_bits_uop_iq_type;
      5'b10101:
        casez_tmp_299 = ldq_21_bits_uop_iq_type;
      5'b10110:
        casez_tmp_299 = ldq_22_bits_uop_iq_type;
      5'b10111:
        casez_tmp_299 = ldq_23_bits_uop_iq_type;
      5'b11000:
        casez_tmp_299 = ldq_24_bits_uop_iq_type;
      5'b11001:
        casez_tmp_299 = ldq_25_bits_uop_iq_type;
      5'b11010:
        casez_tmp_299 = ldq_26_bits_uop_iq_type;
      5'b11011:
        casez_tmp_299 = ldq_27_bits_uop_iq_type;
      5'b11100:
        casez_tmp_299 = ldq_28_bits_uop_iq_type;
      5'b11101:
        casez_tmp_299 = ldq_29_bits_uop_iq_type;
      5'b11110:
        casez_tmp_299 = ldq_30_bits_uop_iq_type;
      default:
        casez_tmp_299 = ldq_31_bits_uop_iq_type;
    endcase
  end // always @(*)
  reg  [9:0]  casez_tmp_300;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_300 = ldq_0_bits_uop_fu_code;
      5'b00001:
        casez_tmp_300 = ldq_1_bits_uop_fu_code;
      5'b00010:
        casez_tmp_300 = ldq_2_bits_uop_fu_code;
      5'b00011:
        casez_tmp_300 = ldq_3_bits_uop_fu_code;
      5'b00100:
        casez_tmp_300 = ldq_4_bits_uop_fu_code;
      5'b00101:
        casez_tmp_300 = ldq_5_bits_uop_fu_code;
      5'b00110:
        casez_tmp_300 = ldq_6_bits_uop_fu_code;
      5'b00111:
        casez_tmp_300 = ldq_7_bits_uop_fu_code;
      5'b01000:
        casez_tmp_300 = ldq_8_bits_uop_fu_code;
      5'b01001:
        casez_tmp_300 = ldq_9_bits_uop_fu_code;
      5'b01010:
        casez_tmp_300 = ldq_10_bits_uop_fu_code;
      5'b01011:
        casez_tmp_300 = ldq_11_bits_uop_fu_code;
      5'b01100:
        casez_tmp_300 = ldq_12_bits_uop_fu_code;
      5'b01101:
        casez_tmp_300 = ldq_13_bits_uop_fu_code;
      5'b01110:
        casez_tmp_300 = ldq_14_bits_uop_fu_code;
      5'b01111:
        casez_tmp_300 = ldq_15_bits_uop_fu_code;
      5'b10000:
        casez_tmp_300 = ldq_16_bits_uop_fu_code;
      5'b10001:
        casez_tmp_300 = ldq_17_bits_uop_fu_code;
      5'b10010:
        casez_tmp_300 = ldq_18_bits_uop_fu_code;
      5'b10011:
        casez_tmp_300 = ldq_19_bits_uop_fu_code;
      5'b10100:
        casez_tmp_300 = ldq_20_bits_uop_fu_code;
      5'b10101:
        casez_tmp_300 = ldq_21_bits_uop_fu_code;
      5'b10110:
        casez_tmp_300 = ldq_22_bits_uop_fu_code;
      5'b10111:
        casez_tmp_300 = ldq_23_bits_uop_fu_code;
      5'b11000:
        casez_tmp_300 = ldq_24_bits_uop_fu_code;
      5'b11001:
        casez_tmp_300 = ldq_25_bits_uop_fu_code;
      5'b11010:
        casez_tmp_300 = ldq_26_bits_uop_fu_code;
      5'b11011:
        casez_tmp_300 = ldq_27_bits_uop_fu_code;
      5'b11100:
        casez_tmp_300 = ldq_28_bits_uop_fu_code;
      5'b11101:
        casez_tmp_300 = ldq_29_bits_uop_fu_code;
      5'b11110:
        casez_tmp_300 = ldq_30_bits_uop_fu_code;
      default:
        casez_tmp_300 = ldq_31_bits_uop_fu_code;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_301;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_301 = ldq_0_bits_uop_ctrl_br_type;
      5'b00001:
        casez_tmp_301 = ldq_1_bits_uop_ctrl_br_type;
      5'b00010:
        casez_tmp_301 = ldq_2_bits_uop_ctrl_br_type;
      5'b00011:
        casez_tmp_301 = ldq_3_bits_uop_ctrl_br_type;
      5'b00100:
        casez_tmp_301 = ldq_4_bits_uop_ctrl_br_type;
      5'b00101:
        casez_tmp_301 = ldq_5_bits_uop_ctrl_br_type;
      5'b00110:
        casez_tmp_301 = ldq_6_bits_uop_ctrl_br_type;
      5'b00111:
        casez_tmp_301 = ldq_7_bits_uop_ctrl_br_type;
      5'b01000:
        casez_tmp_301 = ldq_8_bits_uop_ctrl_br_type;
      5'b01001:
        casez_tmp_301 = ldq_9_bits_uop_ctrl_br_type;
      5'b01010:
        casez_tmp_301 = ldq_10_bits_uop_ctrl_br_type;
      5'b01011:
        casez_tmp_301 = ldq_11_bits_uop_ctrl_br_type;
      5'b01100:
        casez_tmp_301 = ldq_12_bits_uop_ctrl_br_type;
      5'b01101:
        casez_tmp_301 = ldq_13_bits_uop_ctrl_br_type;
      5'b01110:
        casez_tmp_301 = ldq_14_bits_uop_ctrl_br_type;
      5'b01111:
        casez_tmp_301 = ldq_15_bits_uop_ctrl_br_type;
      5'b10000:
        casez_tmp_301 = ldq_16_bits_uop_ctrl_br_type;
      5'b10001:
        casez_tmp_301 = ldq_17_bits_uop_ctrl_br_type;
      5'b10010:
        casez_tmp_301 = ldq_18_bits_uop_ctrl_br_type;
      5'b10011:
        casez_tmp_301 = ldq_19_bits_uop_ctrl_br_type;
      5'b10100:
        casez_tmp_301 = ldq_20_bits_uop_ctrl_br_type;
      5'b10101:
        casez_tmp_301 = ldq_21_bits_uop_ctrl_br_type;
      5'b10110:
        casez_tmp_301 = ldq_22_bits_uop_ctrl_br_type;
      5'b10111:
        casez_tmp_301 = ldq_23_bits_uop_ctrl_br_type;
      5'b11000:
        casez_tmp_301 = ldq_24_bits_uop_ctrl_br_type;
      5'b11001:
        casez_tmp_301 = ldq_25_bits_uop_ctrl_br_type;
      5'b11010:
        casez_tmp_301 = ldq_26_bits_uop_ctrl_br_type;
      5'b11011:
        casez_tmp_301 = ldq_27_bits_uop_ctrl_br_type;
      5'b11100:
        casez_tmp_301 = ldq_28_bits_uop_ctrl_br_type;
      5'b11101:
        casez_tmp_301 = ldq_29_bits_uop_ctrl_br_type;
      5'b11110:
        casez_tmp_301 = ldq_30_bits_uop_ctrl_br_type;
      default:
        casez_tmp_301 = ldq_31_bits_uop_ctrl_br_type;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_302;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_302 = ldq_0_bits_uop_ctrl_op1_sel;
      5'b00001:
        casez_tmp_302 = ldq_1_bits_uop_ctrl_op1_sel;
      5'b00010:
        casez_tmp_302 = ldq_2_bits_uop_ctrl_op1_sel;
      5'b00011:
        casez_tmp_302 = ldq_3_bits_uop_ctrl_op1_sel;
      5'b00100:
        casez_tmp_302 = ldq_4_bits_uop_ctrl_op1_sel;
      5'b00101:
        casez_tmp_302 = ldq_5_bits_uop_ctrl_op1_sel;
      5'b00110:
        casez_tmp_302 = ldq_6_bits_uop_ctrl_op1_sel;
      5'b00111:
        casez_tmp_302 = ldq_7_bits_uop_ctrl_op1_sel;
      5'b01000:
        casez_tmp_302 = ldq_8_bits_uop_ctrl_op1_sel;
      5'b01001:
        casez_tmp_302 = ldq_9_bits_uop_ctrl_op1_sel;
      5'b01010:
        casez_tmp_302 = ldq_10_bits_uop_ctrl_op1_sel;
      5'b01011:
        casez_tmp_302 = ldq_11_bits_uop_ctrl_op1_sel;
      5'b01100:
        casez_tmp_302 = ldq_12_bits_uop_ctrl_op1_sel;
      5'b01101:
        casez_tmp_302 = ldq_13_bits_uop_ctrl_op1_sel;
      5'b01110:
        casez_tmp_302 = ldq_14_bits_uop_ctrl_op1_sel;
      5'b01111:
        casez_tmp_302 = ldq_15_bits_uop_ctrl_op1_sel;
      5'b10000:
        casez_tmp_302 = ldq_16_bits_uop_ctrl_op1_sel;
      5'b10001:
        casez_tmp_302 = ldq_17_bits_uop_ctrl_op1_sel;
      5'b10010:
        casez_tmp_302 = ldq_18_bits_uop_ctrl_op1_sel;
      5'b10011:
        casez_tmp_302 = ldq_19_bits_uop_ctrl_op1_sel;
      5'b10100:
        casez_tmp_302 = ldq_20_bits_uop_ctrl_op1_sel;
      5'b10101:
        casez_tmp_302 = ldq_21_bits_uop_ctrl_op1_sel;
      5'b10110:
        casez_tmp_302 = ldq_22_bits_uop_ctrl_op1_sel;
      5'b10111:
        casez_tmp_302 = ldq_23_bits_uop_ctrl_op1_sel;
      5'b11000:
        casez_tmp_302 = ldq_24_bits_uop_ctrl_op1_sel;
      5'b11001:
        casez_tmp_302 = ldq_25_bits_uop_ctrl_op1_sel;
      5'b11010:
        casez_tmp_302 = ldq_26_bits_uop_ctrl_op1_sel;
      5'b11011:
        casez_tmp_302 = ldq_27_bits_uop_ctrl_op1_sel;
      5'b11100:
        casez_tmp_302 = ldq_28_bits_uop_ctrl_op1_sel;
      5'b11101:
        casez_tmp_302 = ldq_29_bits_uop_ctrl_op1_sel;
      5'b11110:
        casez_tmp_302 = ldq_30_bits_uop_ctrl_op1_sel;
      default:
        casez_tmp_302 = ldq_31_bits_uop_ctrl_op1_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_303;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_303 = ldq_0_bits_uop_ctrl_op2_sel;
      5'b00001:
        casez_tmp_303 = ldq_1_bits_uop_ctrl_op2_sel;
      5'b00010:
        casez_tmp_303 = ldq_2_bits_uop_ctrl_op2_sel;
      5'b00011:
        casez_tmp_303 = ldq_3_bits_uop_ctrl_op2_sel;
      5'b00100:
        casez_tmp_303 = ldq_4_bits_uop_ctrl_op2_sel;
      5'b00101:
        casez_tmp_303 = ldq_5_bits_uop_ctrl_op2_sel;
      5'b00110:
        casez_tmp_303 = ldq_6_bits_uop_ctrl_op2_sel;
      5'b00111:
        casez_tmp_303 = ldq_7_bits_uop_ctrl_op2_sel;
      5'b01000:
        casez_tmp_303 = ldq_8_bits_uop_ctrl_op2_sel;
      5'b01001:
        casez_tmp_303 = ldq_9_bits_uop_ctrl_op2_sel;
      5'b01010:
        casez_tmp_303 = ldq_10_bits_uop_ctrl_op2_sel;
      5'b01011:
        casez_tmp_303 = ldq_11_bits_uop_ctrl_op2_sel;
      5'b01100:
        casez_tmp_303 = ldq_12_bits_uop_ctrl_op2_sel;
      5'b01101:
        casez_tmp_303 = ldq_13_bits_uop_ctrl_op2_sel;
      5'b01110:
        casez_tmp_303 = ldq_14_bits_uop_ctrl_op2_sel;
      5'b01111:
        casez_tmp_303 = ldq_15_bits_uop_ctrl_op2_sel;
      5'b10000:
        casez_tmp_303 = ldq_16_bits_uop_ctrl_op2_sel;
      5'b10001:
        casez_tmp_303 = ldq_17_bits_uop_ctrl_op2_sel;
      5'b10010:
        casez_tmp_303 = ldq_18_bits_uop_ctrl_op2_sel;
      5'b10011:
        casez_tmp_303 = ldq_19_bits_uop_ctrl_op2_sel;
      5'b10100:
        casez_tmp_303 = ldq_20_bits_uop_ctrl_op2_sel;
      5'b10101:
        casez_tmp_303 = ldq_21_bits_uop_ctrl_op2_sel;
      5'b10110:
        casez_tmp_303 = ldq_22_bits_uop_ctrl_op2_sel;
      5'b10111:
        casez_tmp_303 = ldq_23_bits_uop_ctrl_op2_sel;
      5'b11000:
        casez_tmp_303 = ldq_24_bits_uop_ctrl_op2_sel;
      5'b11001:
        casez_tmp_303 = ldq_25_bits_uop_ctrl_op2_sel;
      5'b11010:
        casez_tmp_303 = ldq_26_bits_uop_ctrl_op2_sel;
      5'b11011:
        casez_tmp_303 = ldq_27_bits_uop_ctrl_op2_sel;
      5'b11100:
        casez_tmp_303 = ldq_28_bits_uop_ctrl_op2_sel;
      5'b11101:
        casez_tmp_303 = ldq_29_bits_uop_ctrl_op2_sel;
      5'b11110:
        casez_tmp_303 = ldq_30_bits_uop_ctrl_op2_sel;
      default:
        casez_tmp_303 = ldq_31_bits_uop_ctrl_op2_sel;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_304;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_304 = ldq_0_bits_uop_ctrl_imm_sel;
      5'b00001:
        casez_tmp_304 = ldq_1_bits_uop_ctrl_imm_sel;
      5'b00010:
        casez_tmp_304 = ldq_2_bits_uop_ctrl_imm_sel;
      5'b00011:
        casez_tmp_304 = ldq_3_bits_uop_ctrl_imm_sel;
      5'b00100:
        casez_tmp_304 = ldq_4_bits_uop_ctrl_imm_sel;
      5'b00101:
        casez_tmp_304 = ldq_5_bits_uop_ctrl_imm_sel;
      5'b00110:
        casez_tmp_304 = ldq_6_bits_uop_ctrl_imm_sel;
      5'b00111:
        casez_tmp_304 = ldq_7_bits_uop_ctrl_imm_sel;
      5'b01000:
        casez_tmp_304 = ldq_8_bits_uop_ctrl_imm_sel;
      5'b01001:
        casez_tmp_304 = ldq_9_bits_uop_ctrl_imm_sel;
      5'b01010:
        casez_tmp_304 = ldq_10_bits_uop_ctrl_imm_sel;
      5'b01011:
        casez_tmp_304 = ldq_11_bits_uop_ctrl_imm_sel;
      5'b01100:
        casez_tmp_304 = ldq_12_bits_uop_ctrl_imm_sel;
      5'b01101:
        casez_tmp_304 = ldq_13_bits_uop_ctrl_imm_sel;
      5'b01110:
        casez_tmp_304 = ldq_14_bits_uop_ctrl_imm_sel;
      5'b01111:
        casez_tmp_304 = ldq_15_bits_uop_ctrl_imm_sel;
      5'b10000:
        casez_tmp_304 = ldq_16_bits_uop_ctrl_imm_sel;
      5'b10001:
        casez_tmp_304 = ldq_17_bits_uop_ctrl_imm_sel;
      5'b10010:
        casez_tmp_304 = ldq_18_bits_uop_ctrl_imm_sel;
      5'b10011:
        casez_tmp_304 = ldq_19_bits_uop_ctrl_imm_sel;
      5'b10100:
        casez_tmp_304 = ldq_20_bits_uop_ctrl_imm_sel;
      5'b10101:
        casez_tmp_304 = ldq_21_bits_uop_ctrl_imm_sel;
      5'b10110:
        casez_tmp_304 = ldq_22_bits_uop_ctrl_imm_sel;
      5'b10111:
        casez_tmp_304 = ldq_23_bits_uop_ctrl_imm_sel;
      5'b11000:
        casez_tmp_304 = ldq_24_bits_uop_ctrl_imm_sel;
      5'b11001:
        casez_tmp_304 = ldq_25_bits_uop_ctrl_imm_sel;
      5'b11010:
        casez_tmp_304 = ldq_26_bits_uop_ctrl_imm_sel;
      5'b11011:
        casez_tmp_304 = ldq_27_bits_uop_ctrl_imm_sel;
      5'b11100:
        casez_tmp_304 = ldq_28_bits_uop_ctrl_imm_sel;
      5'b11101:
        casez_tmp_304 = ldq_29_bits_uop_ctrl_imm_sel;
      5'b11110:
        casez_tmp_304 = ldq_30_bits_uop_ctrl_imm_sel;
      default:
        casez_tmp_304 = ldq_31_bits_uop_ctrl_imm_sel;
    endcase
  end // always @(*)
  reg  [3:0]  casez_tmp_305;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_305 = ldq_0_bits_uop_ctrl_op_fcn;
      5'b00001:
        casez_tmp_305 = ldq_1_bits_uop_ctrl_op_fcn;
      5'b00010:
        casez_tmp_305 = ldq_2_bits_uop_ctrl_op_fcn;
      5'b00011:
        casez_tmp_305 = ldq_3_bits_uop_ctrl_op_fcn;
      5'b00100:
        casez_tmp_305 = ldq_4_bits_uop_ctrl_op_fcn;
      5'b00101:
        casez_tmp_305 = ldq_5_bits_uop_ctrl_op_fcn;
      5'b00110:
        casez_tmp_305 = ldq_6_bits_uop_ctrl_op_fcn;
      5'b00111:
        casez_tmp_305 = ldq_7_bits_uop_ctrl_op_fcn;
      5'b01000:
        casez_tmp_305 = ldq_8_bits_uop_ctrl_op_fcn;
      5'b01001:
        casez_tmp_305 = ldq_9_bits_uop_ctrl_op_fcn;
      5'b01010:
        casez_tmp_305 = ldq_10_bits_uop_ctrl_op_fcn;
      5'b01011:
        casez_tmp_305 = ldq_11_bits_uop_ctrl_op_fcn;
      5'b01100:
        casez_tmp_305 = ldq_12_bits_uop_ctrl_op_fcn;
      5'b01101:
        casez_tmp_305 = ldq_13_bits_uop_ctrl_op_fcn;
      5'b01110:
        casez_tmp_305 = ldq_14_bits_uop_ctrl_op_fcn;
      5'b01111:
        casez_tmp_305 = ldq_15_bits_uop_ctrl_op_fcn;
      5'b10000:
        casez_tmp_305 = ldq_16_bits_uop_ctrl_op_fcn;
      5'b10001:
        casez_tmp_305 = ldq_17_bits_uop_ctrl_op_fcn;
      5'b10010:
        casez_tmp_305 = ldq_18_bits_uop_ctrl_op_fcn;
      5'b10011:
        casez_tmp_305 = ldq_19_bits_uop_ctrl_op_fcn;
      5'b10100:
        casez_tmp_305 = ldq_20_bits_uop_ctrl_op_fcn;
      5'b10101:
        casez_tmp_305 = ldq_21_bits_uop_ctrl_op_fcn;
      5'b10110:
        casez_tmp_305 = ldq_22_bits_uop_ctrl_op_fcn;
      5'b10111:
        casez_tmp_305 = ldq_23_bits_uop_ctrl_op_fcn;
      5'b11000:
        casez_tmp_305 = ldq_24_bits_uop_ctrl_op_fcn;
      5'b11001:
        casez_tmp_305 = ldq_25_bits_uop_ctrl_op_fcn;
      5'b11010:
        casez_tmp_305 = ldq_26_bits_uop_ctrl_op_fcn;
      5'b11011:
        casez_tmp_305 = ldq_27_bits_uop_ctrl_op_fcn;
      5'b11100:
        casez_tmp_305 = ldq_28_bits_uop_ctrl_op_fcn;
      5'b11101:
        casez_tmp_305 = ldq_29_bits_uop_ctrl_op_fcn;
      5'b11110:
        casez_tmp_305 = ldq_30_bits_uop_ctrl_op_fcn;
      default:
        casez_tmp_305 = ldq_31_bits_uop_ctrl_op_fcn;
    endcase
  end // always @(*)
  reg         casez_tmp_306;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_306 = ldq_0_bits_uop_ctrl_fcn_dw;
      5'b00001:
        casez_tmp_306 = ldq_1_bits_uop_ctrl_fcn_dw;
      5'b00010:
        casez_tmp_306 = ldq_2_bits_uop_ctrl_fcn_dw;
      5'b00011:
        casez_tmp_306 = ldq_3_bits_uop_ctrl_fcn_dw;
      5'b00100:
        casez_tmp_306 = ldq_4_bits_uop_ctrl_fcn_dw;
      5'b00101:
        casez_tmp_306 = ldq_5_bits_uop_ctrl_fcn_dw;
      5'b00110:
        casez_tmp_306 = ldq_6_bits_uop_ctrl_fcn_dw;
      5'b00111:
        casez_tmp_306 = ldq_7_bits_uop_ctrl_fcn_dw;
      5'b01000:
        casez_tmp_306 = ldq_8_bits_uop_ctrl_fcn_dw;
      5'b01001:
        casez_tmp_306 = ldq_9_bits_uop_ctrl_fcn_dw;
      5'b01010:
        casez_tmp_306 = ldq_10_bits_uop_ctrl_fcn_dw;
      5'b01011:
        casez_tmp_306 = ldq_11_bits_uop_ctrl_fcn_dw;
      5'b01100:
        casez_tmp_306 = ldq_12_bits_uop_ctrl_fcn_dw;
      5'b01101:
        casez_tmp_306 = ldq_13_bits_uop_ctrl_fcn_dw;
      5'b01110:
        casez_tmp_306 = ldq_14_bits_uop_ctrl_fcn_dw;
      5'b01111:
        casez_tmp_306 = ldq_15_bits_uop_ctrl_fcn_dw;
      5'b10000:
        casez_tmp_306 = ldq_16_bits_uop_ctrl_fcn_dw;
      5'b10001:
        casez_tmp_306 = ldq_17_bits_uop_ctrl_fcn_dw;
      5'b10010:
        casez_tmp_306 = ldq_18_bits_uop_ctrl_fcn_dw;
      5'b10011:
        casez_tmp_306 = ldq_19_bits_uop_ctrl_fcn_dw;
      5'b10100:
        casez_tmp_306 = ldq_20_bits_uop_ctrl_fcn_dw;
      5'b10101:
        casez_tmp_306 = ldq_21_bits_uop_ctrl_fcn_dw;
      5'b10110:
        casez_tmp_306 = ldq_22_bits_uop_ctrl_fcn_dw;
      5'b10111:
        casez_tmp_306 = ldq_23_bits_uop_ctrl_fcn_dw;
      5'b11000:
        casez_tmp_306 = ldq_24_bits_uop_ctrl_fcn_dw;
      5'b11001:
        casez_tmp_306 = ldq_25_bits_uop_ctrl_fcn_dw;
      5'b11010:
        casez_tmp_306 = ldq_26_bits_uop_ctrl_fcn_dw;
      5'b11011:
        casez_tmp_306 = ldq_27_bits_uop_ctrl_fcn_dw;
      5'b11100:
        casez_tmp_306 = ldq_28_bits_uop_ctrl_fcn_dw;
      5'b11101:
        casez_tmp_306 = ldq_29_bits_uop_ctrl_fcn_dw;
      5'b11110:
        casez_tmp_306 = ldq_30_bits_uop_ctrl_fcn_dw;
      default:
        casez_tmp_306 = ldq_31_bits_uop_ctrl_fcn_dw;
    endcase
  end // always @(*)
  reg  [2:0]  casez_tmp_307;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_307 = ldq_0_bits_uop_ctrl_csr_cmd;
      5'b00001:
        casez_tmp_307 = ldq_1_bits_uop_ctrl_csr_cmd;
      5'b00010:
        casez_tmp_307 = ldq_2_bits_uop_ctrl_csr_cmd;
      5'b00011:
        casez_tmp_307 = ldq_3_bits_uop_ctrl_csr_cmd;
      5'b00100:
        casez_tmp_307 = ldq_4_bits_uop_ctrl_csr_cmd;
      5'b00101:
        casez_tmp_307 = ldq_5_bits_uop_ctrl_csr_cmd;
      5'b00110:
        casez_tmp_307 = ldq_6_bits_uop_ctrl_csr_cmd;
      5'b00111:
        casez_tmp_307 = ldq_7_bits_uop_ctrl_csr_cmd;
      5'b01000:
        casez_tmp_307 = ldq_8_bits_uop_ctrl_csr_cmd;
      5'b01001:
        casez_tmp_307 = ldq_9_bits_uop_ctrl_csr_cmd;
      5'b01010:
        casez_tmp_307 = ldq_10_bits_uop_ctrl_csr_cmd;
      5'b01011:
        casez_tmp_307 = ldq_11_bits_uop_ctrl_csr_cmd;
      5'b01100:
        casez_tmp_307 = ldq_12_bits_uop_ctrl_csr_cmd;
      5'b01101:
        casez_tmp_307 = ldq_13_bits_uop_ctrl_csr_cmd;
      5'b01110:
        casez_tmp_307 = ldq_14_bits_uop_ctrl_csr_cmd;
      5'b01111:
        casez_tmp_307 = ldq_15_bits_uop_ctrl_csr_cmd;
      5'b10000:
        casez_tmp_307 = ldq_16_bits_uop_ctrl_csr_cmd;
      5'b10001:
        casez_tmp_307 = ldq_17_bits_uop_ctrl_csr_cmd;
      5'b10010:
        casez_tmp_307 = ldq_18_bits_uop_ctrl_csr_cmd;
      5'b10011:
        casez_tmp_307 = ldq_19_bits_uop_ctrl_csr_cmd;
      5'b10100:
        casez_tmp_307 = ldq_20_bits_uop_ctrl_csr_cmd;
      5'b10101:
        casez_tmp_307 = ldq_21_bits_uop_ctrl_csr_cmd;
      5'b10110:
        casez_tmp_307 = ldq_22_bits_uop_ctrl_csr_cmd;
      5'b10111:
        casez_tmp_307 = ldq_23_bits_uop_ctrl_csr_cmd;
      5'b11000:
        casez_tmp_307 = ldq_24_bits_uop_ctrl_csr_cmd;
      5'b11001:
        casez_tmp_307 = ldq_25_bits_uop_ctrl_csr_cmd;
      5'b11010:
        casez_tmp_307 = ldq_26_bits_uop_ctrl_csr_cmd;
      5'b11011:
        casez_tmp_307 = ldq_27_bits_uop_ctrl_csr_cmd;
      5'b11100:
        casez_tmp_307 = ldq_28_bits_uop_ctrl_csr_cmd;
      5'b11101:
        casez_tmp_307 = ldq_29_bits_uop_ctrl_csr_cmd;
      5'b11110:
        casez_tmp_307 = ldq_30_bits_uop_ctrl_csr_cmd;
      default:
        casez_tmp_307 = ldq_31_bits_uop_ctrl_csr_cmd;
    endcase
  end // always @(*)
  reg         casez_tmp_308;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_308 = ldq_0_bits_uop_ctrl_is_load;
      5'b00001:
        casez_tmp_308 = ldq_1_bits_uop_ctrl_is_load;
      5'b00010:
        casez_tmp_308 = ldq_2_bits_uop_ctrl_is_load;
      5'b00011:
        casez_tmp_308 = ldq_3_bits_uop_ctrl_is_load;
      5'b00100:
        casez_tmp_308 = ldq_4_bits_uop_ctrl_is_load;
      5'b00101:
        casez_tmp_308 = ldq_5_bits_uop_ctrl_is_load;
      5'b00110:
        casez_tmp_308 = ldq_6_bits_uop_ctrl_is_load;
      5'b00111:
        casez_tmp_308 = ldq_7_bits_uop_ctrl_is_load;
      5'b01000:
        casez_tmp_308 = ldq_8_bits_uop_ctrl_is_load;
      5'b01001:
        casez_tmp_308 = ldq_9_bits_uop_ctrl_is_load;
      5'b01010:
        casez_tmp_308 = ldq_10_bits_uop_ctrl_is_load;
      5'b01011:
        casez_tmp_308 = ldq_11_bits_uop_ctrl_is_load;
      5'b01100:
        casez_tmp_308 = ldq_12_bits_uop_ctrl_is_load;
      5'b01101:
        casez_tmp_308 = ldq_13_bits_uop_ctrl_is_load;
      5'b01110:
        casez_tmp_308 = ldq_14_bits_uop_ctrl_is_load;
      5'b01111:
        casez_tmp_308 = ldq_15_bits_uop_ctrl_is_load;
      5'b10000:
        casez_tmp_308 = ldq_16_bits_uop_ctrl_is_load;
      5'b10001:
        casez_tmp_308 = ldq_17_bits_uop_ctrl_is_load;
      5'b10010:
        casez_tmp_308 = ldq_18_bits_uop_ctrl_is_load;
      5'b10011:
        casez_tmp_308 = ldq_19_bits_uop_ctrl_is_load;
      5'b10100:
        casez_tmp_308 = ldq_20_bits_uop_ctrl_is_load;
      5'b10101:
        casez_tmp_308 = ldq_21_bits_uop_ctrl_is_load;
      5'b10110:
        casez_tmp_308 = ldq_22_bits_uop_ctrl_is_load;
      5'b10111:
        casez_tmp_308 = ldq_23_bits_uop_ctrl_is_load;
      5'b11000:
        casez_tmp_308 = ldq_24_bits_uop_ctrl_is_load;
      5'b11001:
        casez_tmp_308 = ldq_25_bits_uop_ctrl_is_load;
      5'b11010:
        casez_tmp_308 = ldq_26_bits_uop_ctrl_is_load;
      5'b11011:
        casez_tmp_308 = ldq_27_bits_uop_ctrl_is_load;
      5'b11100:
        casez_tmp_308 = ldq_28_bits_uop_ctrl_is_load;
      5'b11101:
        casez_tmp_308 = ldq_29_bits_uop_ctrl_is_load;
      5'b11110:
        casez_tmp_308 = ldq_30_bits_uop_ctrl_is_load;
      default:
        casez_tmp_308 = ldq_31_bits_uop_ctrl_is_load;
    endcase
  end // always @(*)
  reg         casez_tmp_309;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_309 = ldq_0_bits_uop_ctrl_is_sta;
      5'b00001:
        casez_tmp_309 = ldq_1_bits_uop_ctrl_is_sta;
      5'b00010:
        casez_tmp_309 = ldq_2_bits_uop_ctrl_is_sta;
      5'b00011:
        casez_tmp_309 = ldq_3_bits_uop_ctrl_is_sta;
      5'b00100:
        casez_tmp_309 = ldq_4_bits_uop_ctrl_is_sta;
      5'b00101:
        casez_tmp_309 = ldq_5_bits_uop_ctrl_is_sta;
      5'b00110:
        casez_tmp_309 = ldq_6_bits_uop_ctrl_is_sta;
      5'b00111:
        casez_tmp_309 = ldq_7_bits_uop_ctrl_is_sta;
      5'b01000:
        casez_tmp_309 = ldq_8_bits_uop_ctrl_is_sta;
      5'b01001:
        casez_tmp_309 = ldq_9_bits_uop_ctrl_is_sta;
      5'b01010:
        casez_tmp_309 = ldq_10_bits_uop_ctrl_is_sta;
      5'b01011:
        casez_tmp_309 = ldq_11_bits_uop_ctrl_is_sta;
      5'b01100:
        casez_tmp_309 = ldq_12_bits_uop_ctrl_is_sta;
      5'b01101:
        casez_tmp_309 = ldq_13_bits_uop_ctrl_is_sta;
      5'b01110:
        casez_tmp_309 = ldq_14_bits_uop_ctrl_is_sta;
      5'b01111:
        casez_tmp_309 = ldq_15_bits_uop_ctrl_is_sta;
      5'b10000:
        casez_tmp_309 = ldq_16_bits_uop_ctrl_is_sta;
      5'b10001:
        casez_tmp_309 = ldq_17_bits_uop_ctrl_is_sta;
      5'b10010:
        casez_tmp_309 = ldq_18_bits_uop_ctrl_is_sta;
      5'b10011:
        casez_tmp_309 = ldq_19_bits_uop_ctrl_is_sta;
      5'b10100:
        casez_tmp_309 = ldq_20_bits_uop_ctrl_is_sta;
      5'b10101:
        casez_tmp_309 = ldq_21_bits_uop_ctrl_is_sta;
      5'b10110:
        casez_tmp_309 = ldq_22_bits_uop_ctrl_is_sta;
      5'b10111:
        casez_tmp_309 = ldq_23_bits_uop_ctrl_is_sta;
      5'b11000:
        casez_tmp_309 = ldq_24_bits_uop_ctrl_is_sta;
      5'b11001:
        casez_tmp_309 = ldq_25_bits_uop_ctrl_is_sta;
      5'b11010:
        casez_tmp_309 = ldq_26_bits_uop_ctrl_is_sta;
      5'b11011:
        casez_tmp_309 = ldq_27_bits_uop_ctrl_is_sta;
      5'b11100:
        casez_tmp_309 = ldq_28_bits_uop_ctrl_is_sta;
      5'b11101:
        casez_tmp_309 = ldq_29_bits_uop_ctrl_is_sta;
      5'b11110:
        casez_tmp_309 = ldq_30_bits_uop_ctrl_is_sta;
      default:
        casez_tmp_309 = ldq_31_bits_uop_ctrl_is_sta;
    endcase
  end // always @(*)
  reg         casez_tmp_310;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_310 = ldq_0_bits_uop_ctrl_is_std;
      5'b00001:
        casez_tmp_310 = ldq_1_bits_uop_ctrl_is_std;
      5'b00010:
        casez_tmp_310 = ldq_2_bits_uop_ctrl_is_std;
      5'b00011:
        casez_tmp_310 = ldq_3_bits_uop_ctrl_is_std;
      5'b00100:
        casez_tmp_310 = ldq_4_bits_uop_ctrl_is_std;
      5'b00101:
        casez_tmp_310 = ldq_5_bits_uop_ctrl_is_std;
      5'b00110:
        casez_tmp_310 = ldq_6_bits_uop_ctrl_is_std;
      5'b00111:
        casez_tmp_310 = ldq_7_bits_uop_ctrl_is_std;
      5'b01000:
        casez_tmp_310 = ldq_8_bits_uop_ctrl_is_std;
      5'b01001:
        casez_tmp_310 = ldq_9_bits_uop_ctrl_is_std;
      5'b01010:
        casez_tmp_310 = ldq_10_bits_uop_ctrl_is_std;
      5'b01011:
        casez_tmp_310 = ldq_11_bits_uop_ctrl_is_std;
      5'b01100:
        casez_tmp_310 = ldq_12_bits_uop_ctrl_is_std;
      5'b01101:
        casez_tmp_310 = ldq_13_bits_uop_ctrl_is_std;
      5'b01110:
        casez_tmp_310 = ldq_14_bits_uop_ctrl_is_std;
      5'b01111:
        casez_tmp_310 = ldq_15_bits_uop_ctrl_is_std;
      5'b10000:
        casez_tmp_310 = ldq_16_bits_uop_ctrl_is_std;
      5'b10001:
        casez_tmp_310 = ldq_17_bits_uop_ctrl_is_std;
      5'b10010:
        casez_tmp_310 = ldq_18_bits_uop_ctrl_is_std;
      5'b10011:
        casez_tmp_310 = ldq_19_bits_uop_ctrl_is_std;
      5'b10100:
        casez_tmp_310 = ldq_20_bits_uop_ctrl_is_std;
      5'b10101:
        casez_tmp_310 = ldq_21_bits_uop_ctrl_is_std;
      5'b10110:
        casez_tmp_310 = ldq_22_bits_uop_ctrl_is_std;
      5'b10111:
        casez_tmp_310 = ldq_23_bits_uop_ctrl_is_std;
      5'b11000:
        casez_tmp_310 = ldq_24_bits_uop_ctrl_is_std;
      5'b11001:
        casez_tmp_310 = ldq_25_bits_uop_ctrl_is_std;
      5'b11010:
        casez_tmp_310 = ldq_26_bits_uop_ctrl_is_std;
      5'b11011:
        casez_tmp_310 = ldq_27_bits_uop_ctrl_is_std;
      5'b11100:
        casez_tmp_310 = ldq_28_bits_uop_ctrl_is_std;
      5'b11101:
        casez_tmp_310 = ldq_29_bits_uop_ctrl_is_std;
      5'b11110:
        casez_tmp_310 = ldq_30_bits_uop_ctrl_is_std;
      default:
        casez_tmp_310 = ldq_31_bits_uop_ctrl_is_std;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_311;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_311 = ldq_0_bits_uop_iw_state;
      5'b00001:
        casez_tmp_311 = ldq_1_bits_uop_iw_state;
      5'b00010:
        casez_tmp_311 = ldq_2_bits_uop_iw_state;
      5'b00011:
        casez_tmp_311 = ldq_3_bits_uop_iw_state;
      5'b00100:
        casez_tmp_311 = ldq_4_bits_uop_iw_state;
      5'b00101:
        casez_tmp_311 = ldq_5_bits_uop_iw_state;
      5'b00110:
        casez_tmp_311 = ldq_6_bits_uop_iw_state;
      5'b00111:
        casez_tmp_311 = ldq_7_bits_uop_iw_state;
      5'b01000:
        casez_tmp_311 = ldq_8_bits_uop_iw_state;
      5'b01001:
        casez_tmp_311 = ldq_9_bits_uop_iw_state;
      5'b01010:
        casez_tmp_311 = ldq_10_bits_uop_iw_state;
      5'b01011:
        casez_tmp_311 = ldq_11_bits_uop_iw_state;
      5'b01100:
        casez_tmp_311 = ldq_12_bits_uop_iw_state;
      5'b01101:
        casez_tmp_311 = ldq_13_bits_uop_iw_state;
      5'b01110:
        casez_tmp_311 = ldq_14_bits_uop_iw_state;
      5'b01111:
        casez_tmp_311 = ldq_15_bits_uop_iw_state;
      5'b10000:
        casez_tmp_311 = ldq_16_bits_uop_iw_state;
      5'b10001:
        casez_tmp_311 = ldq_17_bits_uop_iw_state;
      5'b10010:
        casez_tmp_311 = ldq_18_bits_uop_iw_state;
      5'b10011:
        casez_tmp_311 = ldq_19_bits_uop_iw_state;
      5'b10100:
        casez_tmp_311 = ldq_20_bits_uop_iw_state;
      5'b10101:
        casez_tmp_311 = ldq_21_bits_uop_iw_state;
      5'b10110:
        casez_tmp_311 = ldq_22_bits_uop_iw_state;
      5'b10111:
        casez_tmp_311 = ldq_23_bits_uop_iw_state;
      5'b11000:
        casez_tmp_311 = ldq_24_bits_uop_iw_state;
      5'b11001:
        casez_tmp_311 = ldq_25_bits_uop_iw_state;
      5'b11010:
        casez_tmp_311 = ldq_26_bits_uop_iw_state;
      5'b11011:
        casez_tmp_311 = ldq_27_bits_uop_iw_state;
      5'b11100:
        casez_tmp_311 = ldq_28_bits_uop_iw_state;
      5'b11101:
        casez_tmp_311 = ldq_29_bits_uop_iw_state;
      5'b11110:
        casez_tmp_311 = ldq_30_bits_uop_iw_state;
      default:
        casez_tmp_311 = ldq_31_bits_uop_iw_state;
    endcase
  end // always @(*)
  reg         casez_tmp_312;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_312 = ldq_0_bits_uop_iw_p1_poisoned;
      5'b00001:
        casez_tmp_312 = ldq_1_bits_uop_iw_p1_poisoned;
      5'b00010:
        casez_tmp_312 = ldq_2_bits_uop_iw_p1_poisoned;
      5'b00011:
        casez_tmp_312 = ldq_3_bits_uop_iw_p1_poisoned;
      5'b00100:
        casez_tmp_312 = ldq_4_bits_uop_iw_p1_poisoned;
      5'b00101:
        casez_tmp_312 = ldq_5_bits_uop_iw_p1_poisoned;
      5'b00110:
        casez_tmp_312 = ldq_6_bits_uop_iw_p1_poisoned;
      5'b00111:
        casez_tmp_312 = ldq_7_bits_uop_iw_p1_poisoned;
      5'b01000:
        casez_tmp_312 = ldq_8_bits_uop_iw_p1_poisoned;
      5'b01001:
        casez_tmp_312 = ldq_9_bits_uop_iw_p1_poisoned;
      5'b01010:
        casez_tmp_312 = ldq_10_bits_uop_iw_p1_poisoned;
      5'b01011:
        casez_tmp_312 = ldq_11_bits_uop_iw_p1_poisoned;
      5'b01100:
        casez_tmp_312 = ldq_12_bits_uop_iw_p1_poisoned;
      5'b01101:
        casez_tmp_312 = ldq_13_bits_uop_iw_p1_poisoned;
      5'b01110:
        casez_tmp_312 = ldq_14_bits_uop_iw_p1_poisoned;
      5'b01111:
        casez_tmp_312 = ldq_15_bits_uop_iw_p1_poisoned;
      5'b10000:
        casez_tmp_312 = ldq_16_bits_uop_iw_p1_poisoned;
      5'b10001:
        casez_tmp_312 = ldq_17_bits_uop_iw_p1_poisoned;
      5'b10010:
        casez_tmp_312 = ldq_18_bits_uop_iw_p1_poisoned;
      5'b10011:
        casez_tmp_312 = ldq_19_bits_uop_iw_p1_poisoned;
      5'b10100:
        casez_tmp_312 = ldq_20_bits_uop_iw_p1_poisoned;
      5'b10101:
        casez_tmp_312 = ldq_21_bits_uop_iw_p1_poisoned;
      5'b10110:
        casez_tmp_312 = ldq_22_bits_uop_iw_p1_poisoned;
      5'b10111:
        casez_tmp_312 = ldq_23_bits_uop_iw_p1_poisoned;
      5'b11000:
        casez_tmp_312 = ldq_24_bits_uop_iw_p1_poisoned;
      5'b11001:
        casez_tmp_312 = ldq_25_bits_uop_iw_p1_poisoned;
      5'b11010:
        casez_tmp_312 = ldq_26_bits_uop_iw_p1_poisoned;
      5'b11011:
        casez_tmp_312 = ldq_27_bits_uop_iw_p1_poisoned;
      5'b11100:
        casez_tmp_312 = ldq_28_bits_uop_iw_p1_poisoned;
      5'b11101:
        casez_tmp_312 = ldq_29_bits_uop_iw_p1_poisoned;
      5'b11110:
        casez_tmp_312 = ldq_30_bits_uop_iw_p1_poisoned;
      default:
        casez_tmp_312 = ldq_31_bits_uop_iw_p1_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_313;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_313 = ldq_0_bits_uop_iw_p2_poisoned;
      5'b00001:
        casez_tmp_313 = ldq_1_bits_uop_iw_p2_poisoned;
      5'b00010:
        casez_tmp_313 = ldq_2_bits_uop_iw_p2_poisoned;
      5'b00011:
        casez_tmp_313 = ldq_3_bits_uop_iw_p2_poisoned;
      5'b00100:
        casez_tmp_313 = ldq_4_bits_uop_iw_p2_poisoned;
      5'b00101:
        casez_tmp_313 = ldq_5_bits_uop_iw_p2_poisoned;
      5'b00110:
        casez_tmp_313 = ldq_6_bits_uop_iw_p2_poisoned;
      5'b00111:
        casez_tmp_313 = ldq_7_bits_uop_iw_p2_poisoned;
      5'b01000:
        casez_tmp_313 = ldq_8_bits_uop_iw_p2_poisoned;
      5'b01001:
        casez_tmp_313 = ldq_9_bits_uop_iw_p2_poisoned;
      5'b01010:
        casez_tmp_313 = ldq_10_bits_uop_iw_p2_poisoned;
      5'b01011:
        casez_tmp_313 = ldq_11_bits_uop_iw_p2_poisoned;
      5'b01100:
        casez_tmp_313 = ldq_12_bits_uop_iw_p2_poisoned;
      5'b01101:
        casez_tmp_313 = ldq_13_bits_uop_iw_p2_poisoned;
      5'b01110:
        casez_tmp_313 = ldq_14_bits_uop_iw_p2_poisoned;
      5'b01111:
        casez_tmp_313 = ldq_15_bits_uop_iw_p2_poisoned;
      5'b10000:
        casez_tmp_313 = ldq_16_bits_uop_iw_p2_poisoned;
      5'b10001:
        casez_tmp_313 = ldq_17_bits_uop_iw_p2_poisoned;
      5'b10010:
        casez_tmp_313 = ldq_18_bits_uop_iw_p2_poisoned;
      5'b10011:
        casez_tmp_313 = ldq_19_bits_uop_iw_p2_poisoned;
      5'b10100:
        casez_tmp_313 = ldq_20_bits_uop_iw_p2_poisoned;
      5'b10101:
        casez_tmp_313 = ldq_21_bits_uop_iw_p2_poisoned;
      5'b10110:
        casez_tmp_313 = ldq_22_bits_uop_iw_p2_poisoned;
      5'b10111:
        casez_tmp_313 = ldq_23_bits_uop_iw_p2_poisoned;
      5'b11000:
        casez_tmp_313 = ldq_24_bits_uop_iw_p2_poisoned;
      5'b11001:
        casez_tmp_313 = ldq_25_bits_uop_iw_p2_poisoned;
      5'b11010:
        casez_tmp_313 = ldq_26_bits_uop_iw_p2_poisoned;
      5'b11011:
        casez_tmp_313 = ldq_27_bits_uop_iw_p2_poisoned;
      5'b11100:
        casez_tmp_313 = ldq_28_bits_uop_iw_p2_poisoned;
      5'b11101:
        casez_tmp_313 = ldq_29_bits_uop_iw_p2_poisoned;
      5'b11110:
        casez_tmp_313 = ldq_30_bits_uop_iw_p2_poisoned;
      default:
        casez_tmp_313 = ldq_31_bits_uop_iw_p2_poisoned;
    endcase
  end // always @(*)
  reg         casez_tmp_314;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_314 = ldq_0_bits_uop_is_br;
      5'b00001:
        casez_tmp_314 = ldq_1_bits_uop_is_br;
      5'b00010:
        casez_tmp_314 = ldq_2_bits_uop_is_br;
      5'b00011:
        casez_tmp_314 = ldq_3_bits_uop_is_br;
      5'b00100:
        casez_tmp_314 = ldq_4_bits_uop_is_br;
      5'b00101:
        casez_tmp_314 = ldq_5_bits_uop_is_br;
      5'b00110:
        casez_tmp_314 = ldq_6_bits_uop_is_br;
      5'b00111:
        casez_tmp_314 = ldq_7_bits_uop_is_br;
      5'b01000:
        casez_tmp_314 = ldq_8_bits_uop_is_br;
      5'b01001:
        casez_tmp_314 = ldq_9_bits_uop_is_br;
      5'b01010:
        casez_tmp_314 = ldq_10_bits_uop_is_br;
      5'b01011:
        casez_tmp_314 = ldq_11_bits_uop_is_br;
      5'b01100:
        casez_tmp_314 = ldq_12_bits_uop_is_br;
      5'b01101:
        casez_tmp_314 = ldq_13_bits_uop_is_br;
      5'b01110:
        casez_tmp_314 = ldq_14_bits_uop_is_br;
      5'b01111:
        casez_tmp_314 = ldq_15_bits_uop_is_br;
      5'b10000:
        casez_tmp_314 = ldq_16_bits_uop_is_br;
      5'b10001:
        casez_tmp_314 = ldq_17_bits_uop_is_br;
      5'b10010:
        casez_tmp_314 = ldq_18_bits_uop_is_br;
      5'b10011:
        casez_tmp_314 = ldq_19_bits_uop_is_br;
      5'b10100:
        casez_tmp_314 = ldq_20_bits_uop_is_br;
      5'b10101:
        casez_tmp_314 = ldq_21_bits_uop_is_br;
      5'b10110:
        casez_tmp_314 = ldq_22_bits_uop_is_br;
      5'b10111:
        casez_tmp_314 = ldq_23_bits_uop_is_br;
      5'b11000:
        casez_tmp_314 = ldq_24_bits_uop_is_br;
      5'b11001:
        casez_tmp_314 = ldq_25_bits_uop_is_br;
      5'b11010:
        casez_tmp_314 = ldq_26_bits_uop_is_br;
      5'b11011:
        casez_tmp_314 = ldq_27_bits_uop_is_br;
      5'b11100:
        casez_tmp_314 = ldq_28_bits_uop_is_br;
      5'b11101:
        casez_tmp_314 = ldq_29_bits_uop_is_br;
      5'b11110:
        casez_tmp_314 = ldq_30_bits_uop_is_br;
      default:
        casez_tmp_314 = ldq_31_bits_uop_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_315;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_315 = ldq_0_bits_uop_is_jalr;
      5'b00001:
        casez_tmp_315 = ldq_1_bits_uop_is_jalr;
      5'b00010:
        casez_tmp_315 = ldq_2_bits_uop_is_jalr;
      5'b00011:
        casez_tmp_315 = ldq_3_bits_uop_is_jalr;
      5'b00100:
        casez_tmp_315 = ldq_4_bits_uop_is_jalr;
      5'b00101:
        casez_tmp_315 = ldq_5_bits_uop_is_jalr;
      5'b00110:
        casez_tmp_315 = ldq_6_bits_uop_is_jalr;
      5'b00111:
        casez_tmp_315 = ldq_7_bits_uop_is_jalr;
      5'b01000:
        casez_tmp_315 = ldq_8_bits_uop_is_jalr;
      5'b01001:
        casez_tmp_315 = ldq_9_bits_uop_is_jalr;
      5'b01010:
        casez_tmp_315 = ldq_10_bits_uop_is_jalr;
      5'b01011:
        casez_tmp_315 = ldq_11_bits_uop_is_jalr;
      5'b01100:
        casez_tmp_315 = ldq_12_bits_uop_is_jalr;
      5'b01101:
        casez_tmp_315 = ldq_13_bits_uop_is_jalr;
      5'b01110:
        casez_tmp_315 = ldq_14_bits_uop_is_jalr;
      5'b01111:
        casez_tmp_315 = ldq_15_bits_uop_is_jalr;
      5'b10000:
        casez_tmp_315 = ldq_16_bits_uop_is_jalr;
      5'b10001:
        casez_tmp_315 = ldq_17_bits_uop_is_jalr;
      5'b10010:
        casez_tmp_315 = ldq_18_bits_uop_is_jalr;
      5'b10011:
        casez_tmp_315 = ldq_19_bits_uop_is_jalr;
      5'b10100:
        casez_tmp_315 = ldq_20_bits_uop_is_jalr;
      5'b10101:
        casez_tmp_315 = ldq_21_bits_uop_is_jalr;
      5'b10110:
        casez_tmp_315 = ldq_22_bits_uop_is_jalr;
      5'b10111:
        casez_tmp_315 = ldq_23_bits_uop_is_jalr;
      5'b11000:
        casez_tmp_315 = ldq_24_bits_uop_is_jalr;
      5'b11001:
        casez_tmp_315 = ldq_25_bits_uop_is_jalr;
      5'b11010:
        casez_tmp_315 = ldq_26_bits_uop_is_jalr;
      5'b11011:
        casez_tmp_315 = ldq_27_bits_uop_is_jalr;
      5'b11100:
        casez_tmp_315 = ldq_28_bits_uop_is_jalr;
      5'b11101:
        casez_tmp_315 = ldq_29_bits_uop_is_jalr;
      5'b11110:
        casez_tmp_315 = ldq_30_bits_uop_is_jalr;
      default:
        casez_tmp_315 = ldq_31_bits_uop_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_316;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_316 = ldq_0_bits_uop_is_jal;
      5'b00001:
        casez_tmp_316 = ldq_1_bits_uop_is_jal;
      5'b00010:
        casez_tmp_316 = ldq_2_bits_uop_is_jal;
      5'b00011:
        casez_tmp_316 = ldq_3_bits_uop_is_jal;
      5'b00100:
        casez_tmp_316 = ldq_4_bits_uop_is_jal;
      5'b00101:
        casez_tmp_316 = ldq_5_bits_uop_is_jal;
      5'b00110:
        casez_tmp_316 = ldq_6_bits_uop_is_jal;
      5'b00111:
        casez_tmp_316 = ldq_7_bits_uop_is_jal;
      5'b01000:
        casez_tmp_316 = ldq_8_bits_uop_is_jal;
      5'b01001:
        casez_tmp_316 = ldq_9_bits_uop_is_jal;
      5'b01010:
        casez_tmp_316 = ldq_10_bits_uop_is_jal;
      5'b01011:
        casez_tmp_316 = ldq_11_bits_uop_is_jal;
      5'b01100:
        casez_tmp_316 = ldq_12_bits_uop_is_jal;
      5'b01101:
        casez_tmp_316 = ldq_13_bits_uop_is_jal;
      5'b01110:
        casez_tmp_316 = ldq_14_bits_uop_is_jal;
      5'b01111:
        casez_tmp_316 = ldq_15_bits_uop_is_jal;
      5'b10000:
        casez_tmp_316 = ldq_16_bits_uop_is_jal;
      5'b10001:
        casez_tmp_316 = ldq_17_bits_uop_is_jal;
      5'b10010:
        casez_tmp_316 = ldq_18_bits_uop_is_jal;
      5'b10011:
        casez_tmp_316 = ldq_19_bits_uop_is_jal;
      5'b10100:
        casez_tmp_316 = ldq_20_bits_uop_is_jal;
      5'b10101:
        casez_tmp_316 = ldq_21_bits_uop_is_jal;
      5'b10110:
        casez_tmp_316 = ldq_22_bits_uop_is_jal;
      5'b10111:
        casez_tmp_316 = ldq_23_bits_uop_is_jal;
      5'b11000:
        casez_tmp_316 = ldq_24_bits_uop_is_jal;
      5'b11001:
        casez_tmp_316 = ldq_25_bits_uop_is_jal;
      5'b11010:
        casez_tmp_316 = ldq_26_bits_uop_is_jal;
      5'b11011:
        casez_tmp_316 = ldq_27_bits_uop_is_jal;
      5'b11100:
        casez_tmp_316 = ldq_28_bits_uop_is_jal;
      5'b11101:
        casez_tmp_316 = ldq_29_bits_uop_is_jal;
      5'b11110:
        casez_tmp_316 = ldq_30_bits_uop_is_jal;
      default:
        casez_tmp_316 = ldq_31_bits_uop_is_jal;
    endcase
  end // always @(*)
  reg         casez_tmp_317;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_317 = ldq_0_bits_uop_is_sfb;
      5'b00001:
        casez_tmp_317 = ldq_1_bits_uop_is_sfb;
      5'b00010:
        casez_tmp_317 = ldq_2_bits_uop_is_sfb;
      5'b00011:
        casez_tmp_317 = ldq_3_bits_uop_is_sfb;
      5'b00100:
        casez_tmp_317 = ldq_4_bits_uop_is_sfb;
      5'b00101:
        casez_tmp_317 = ldq_5_bits_uop_is_sfb;
      5'b00110:
        casez_tmp_317 = ldq_6_bits_uop_is_sfb;
      5'b00111:
        casez_tmp_317 = ldq_7_bits_uop_is_sfb;
      5'b01000:
        casez_tmp_317 = ldq_8_bits_uop_is_sfb;
      5'b01001:
        casez_tmp_317 = ldq_9_bits_uop_is_sfb;
      5'b01010:
        casez_tmp_317 = ldq_10_bits_uop_is_sfb;
      5'b01011:
        casez_tmp_317 = ldq_11_bits_uop_is_sfb;
      5'b01100:
        casez_tmp_317 = ldq_12_bits_uop_is_sfb;
      5'b01101:
        casez_tmp_317 = ldq_13_bits_uop_is_sfb;
      5'b01110:
        casez_tmp_317 = ldq_14_bits_uop_is_sfb;
      5'b01111:
        casez_tmp_317 = ldq_15_bits_uop_is_sfb;
      5'b10000:
        casez_tmp_317 = ldq_16_bits_uop_is_sfb;
      5'b10001:
        casez_tmp_317 = ldq_17_bits_uop_is_sfb;
      5'b10010:
        casez_tmp_317 = ldq_18_bits_uop_is_sfb;
      5'b10011:
        casez_tmp_317 = ldq_19_bits_uop_is_sfb;
      5'b10100:
        casez_tmp_317 = ldq_20_bits_uop_is_sfb;
      5'b10101:
        casez_tmp_317 = ldq_21_bits_uop_is_sfb;
      5'b10110:
        casez_tmp_317 = ldq_22_bits_uop_is_sfb;
      5'b10111:
        casez_tmp_317 = ldq_23_bits_uop_is_sfb;
      5'b11000:
        casez_tmp_317 = ldq_24_bits_uop_is_sfb;
      5'b11001:
        casez_tmp_317 = ldq_25_bits_uop_is_sfb;
      5'b11010:
        casez_tmp_317 = ldq_26_bits_uop_is_sfb;
      5'b11011:
        casez_tmp_317 = ldq_27_bits_uop_is_sfb;
      5'b11100:
        casez_tmp_317 = ldq_28_bits_uop_is_sfb;
      5'b11101:
        casez_tmp_317 = ldq_29_bits_uop_is_sfb;
      5'b11110:
        casez_tmp_317 = ldq_30_bits_uop_is_sfb;
      default:
        casez_tmp_317 = ldq_31_bits_uop_is_sfb;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_318;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_318 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_318 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_318 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_318 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_318 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_318 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_318 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_318 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_318 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_318 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_318 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_318 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_318 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_318 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_318 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_318 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_318 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_318 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_318 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_318 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_318 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_318 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_318 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_318 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_318 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_318 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_318 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_318 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_318 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_318 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_318 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_318 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_319;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_319 = ldq_0_bits_uop_br_tag;
      5'b00001:
        casez_tmp_319 = ldq_1_bits_uop_br_tag;
      5'b00010:
        casez_tmp_319 = ldq_2_bits_uop_br_tag;
      5'b00011:
        casez_tmp_319 = ldq_3_bits_uop_br_tag;
      5'b00100:
        casez_tmp_319 = ldq_4_bits_uop_br_tag;
      5'b00101:
        casez_tmp_319 = ldq_5_bits_uop_br_tag;
      5'b00110:
        casez_tmp_319 = ldq_6_bits_uop_br_tag;
      5'b00111:
        casez_tmp_319 = ldq_7_bits_uop_br_tag;
      5'b01000:
        casez_tmp_319 = ldq_8_bits_uop_br_tag;
      5'b01001:
        casez_tmp_319 = ldq_9_bits_uop_br_tag;
      5'b01010:
        casez_tmp_319 = ldq_10_bits_uop_br_tag;
      5'b01011:
        casez_tmp_319 = ldq_11_bits_uop_br_tag;
      5'b01100:
        casez_tmp_319 = ldq_12_bits_uop_br_tag;
      5'b01101:
        casez_tmp_319 = ldq_13_bits_uop_br_tag;
      5'b01110:
        casez_tmp_319 = ldq_14_bits_uop_br_tag;
      5'b01111:
        casez_tmp_319 = ldq_15_bits_uop_br_tag;
      5'b10000:
        casez_tmp_319 = ldq_16_bits_uop_br_tag;
      5'b10001:
        casez_tmp_319 = ldq_17_bits_uop_br_tag;
      5'b10010:
        casez_tmp_319 = ldq_18_bits_uop_br_tag;
      5'b10011:
        casez_tmp_319 = ldq_19_bits_uop_br_tag;
      5'b10100:
        casez_tmp_319 = ldq_20_bits_uop_br_tag;
      5'b10101:
        casez_tmp_319 = ldq_21_bits_uop_br_tag;
      5'b10110:
        casez_tmp_319 = ldq_22_bits_uop_br_tag;
      5'b10111:
        casez_tmp_319 = ldq_23_bits_uop_br_tag;
      5'b11000:
        casez_tmp_319 = ldq_24_bits_uop_br_tag;
      5'b11001:
        casez_tmp_319 = ldq_25_bits_uop_br_tag;
      5'b11010:
        casez_tmp_319 = ldq_26_bits_uop_br_tag;
      5'b11011:
        casez_tmp_319 = ldq_27_bits_uop_br_tag;
      5'b11100:
        casez_tmp_319 = ldq_28_bits_uop_br_tag;
      5'b11101:
        casez_tmp_319 = ldq_29_bits_uop_br_tag;
      5'b11110:
        casez_tmp_319 = ldq_30_bits_uop_br_tag;
      default:
        casez_tmp_319 = ldq_31_bits_uop_br_tag;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_320;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_320 = ldq_0_bits_uop_ftq_idx;
      5'b00001:
        casez_tmp_320 = ldq_1_bits_uop_ftq_idx;
      5'b00010:
        casez_tmp_320 = ldq_2_bits_uop_ftq_idx;
      5'b00011:
        casez_tmp_320 = ldq_3_bits_uop_ftq_idx;
      5'b00100:
        casez_tmp_320 = ldq_4_bits_uop_ftq_idx;
      5'b00101:
        casez_tmp_320 = ldq_5_bits_uop_ftq_idx;
      5'b00110:
        casez_tmp_320 = ldq_6_bits_uop_ftq_idx;
      5'b00111:
        casez_tmp_320 = ldq_7_bits_uop_ftq_idx;
      5'b01000:
        casez_tmp_320 = ldq_8_bits_uop_ftq_idx;
      5'b01001:
        casez_tmp_320 = ldq_9_bits_uop_ftq_idx;
      5'b01010:
        casez_tmp_320 = ldq_10_bits_uop_ftq_idx;
      5'b01011:
        casez_tmp_320 = ldq_11_bits_uop_ftq_idx;
      5'b01100:
        casez_tmp_320 = ldq_12_bits_uop_ftq_idx;
      5'b01101:
        casez_tmp_320 = ldq_13_bits_uop_ftq_idx;
      5'b01110:
        casez_tmp_320 = ldq_14_bits_uop_ftq_idx;
      5'b01111:
        casez_tmp_320 = ldq_15_bits_uop_ftq_idx;
      5'b10000:
        casez_tmp_320 = ldq_16_bits_uop_ftq_idx;
      5'b10001:
        casez_tmp_320 = ldq_17_bits_uop_ftq_idx;
      5'b10010:
        casez_tmp_320 = ldq_18_bits_uop_ftq_idx;
      5'b10011:
        casez_tmp_320 = ldq_19_bits_uop_ftq_idx;
      5'b10100:
        casez_tmp_320 = ldq_20_bits_uop_ftq_idx;
      5'b10101:
        casez_tmp_320 = ldq_21_bits_uop_ftq_idx;
      5'b10110:
        casez_tmp_320 = ldq_22_bits_uop_ftq_idx;
      5'b10111:
        casez_tmp_320 = ldq_23_bits_uop_ftq_idx;
      5'b11000:
        casez_tmp_320 = ldq_24_bits_uop_ftq_idx;
      5'b11001:
        casez_tmp_320 = ldq_25_bits_uop_ftq_idx;
      5'b11010:
        casez_tmp_320 = ldq_26_bits_uop_ftq_idx;
      5'b11011:
        casez_tmp_320 = ldq_27_bits_uop_ftq_idx;
      5'b11100:
        casez_tmp_320 = ldq_28_bits_uop_ftq_idx;
      5'b11101:
        casez_tmp_320 = ldq_29_bits_uop_ftq_idx;
      5'b11110:
        casez_tmp_320 = ldq_30_bits_uop_ftq_idx;
      default:
        casez_tmp_320 = ldq_31_bits_uop_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_321;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_321 = ldq_0_bits_uop_edge_inst;
      5'b00001:
        casez_tmp_321 = ldq_1_bits_uop_edge_inst;
      5'b00010:
        casez_tmp_321 = ldq_2_bits_uop_edge_inst;
      5'b00011:
        casez_tmp_321 = ldq_3_bits_uop_edge_inst;
      5'b00100:
        casez_tmp_321 = ldq_4_bits_uop_edge_inst;
      5'b00101:
        casez_tmp_321 = ldq_5_bits_uop_edge_inst;
      5'b00110:
        casez_tmp_321 = ldq_6_bits_uop_edge_inst;
      5'b00111:
        casez_tmp_321 = ldq_7_bits_uop_edge_inst;
      5'b01000:
        casez_tmp_321 = ldq_8_bits_uop_edge_inst;
      5'b01001:
        casez_tmp_321 = ldq_9_bits_uop_edge_inst;
      5'b01010:
        casez_tmp_321 = ldq_10_bits_uop_edge_inst;
      5'b01011:
        casez_tmp_321 = ldq_11_bits_uop_edge_inst;
      5'b01100:
        casez_tmp_321 = ldq_12_bits_uop_edge_inst;
      5'b01101:
        casez_tmp_321 = ldq_13_bits_uop_edge_inst;
      5'b01110:
        casez_tmp_321 = ldq_14_bits_uop_edge_inst;
      5'b01111:
        casez_tmp_321 = ldq_15_bits_uop_edge_inst;
      5'b10000:
        casez_tmp_321 = ldq_16_bits_uop_edge_inst;
      5'b10001:
        casez_tmp_321 = ldq_17_bits_uop_edge_inst;
      5'b10010:
        casez_tmp_321 = ldq_18_bits_uop_edge_inst;
      5'b10011:
        casez_tmp_321 = ldq_19_bits_uop_edge_inst;
      5'b10100:
        casez_tmp_321 = ldq_20_bits_uop_edge_inst;
      5'b10101:
        casez_tmp_321 = ldq_21_bits_uop_edge_inst;
      5'b10110:
        casez_tmp_321 = ldq_22_bits_uop_edge_inst;
      5'b10111:
        casez_tmp_321 = ldq_23_bits_uop_edge_inst;
      5'b11000:
        casez_tmp_321 = ldq_24_bits_uop_edge_inst;
      5'b11001:
        casez_tmp_321 = ldq_25_bits_uop_edge_inst;
      5'b11010:
        casez_tmp_321 = ldq_26_bits_uop_edge_inst;
      5'b11011:
        casez_tmp_321 = ldq_27_bits_uop_edge_inst;
      5'b11100:
        casez_tmp_321 = ldq_28_bits_uop_edge_inst;
      5'b11101:
        casez_tmp_321 = ldq_29_bits_uop_edge_inst;
      5'b11110:
        casez_tmp_321 = ldq_30_bits_uop_edge_inst;
      default:
        casez_tmp_321 = ldq_31_bits_uop_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_322;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_322 = ldq_0_bits_uop_pc_lob;
      5'b00001:
        casez_tmp_322 = ldq_1_bits_uop_pc_lob;
      5'b00010:
        casez_tmp_322 = ldq_2_bits_uop_pc_lob;
      5'b00011:
        casez_tmp_322 = ldq_3_bits_uop_pc_lob;
      5'b00100:
        casez_tmp_322 = ldq_4_bits_uop_pc_lob;
      5'b00101:
        casez_tmp_322 = ldq_5_bits_uop_pc_lob;
      5'b00110:
        casez_tmp_322 = ldq_6_bits_uop_pc_lob;
      5'b00111:
        casez_tmp_322 = ldq_7_bits_uop_pc_lob;
      5'b01000:
        casez_tmp_322 = ldq_8_bits_uop_pc_lob;
      5'b01001:
        casez_tmp_322 = ldq_9_bits_uop_pc_lob;
      5'b01010:
        casez_tmp_322 = ldq_10_bits_uop_pc_lob;
      5'b01011:
        casez_tmp_322 = ldq_11_bits_uop_pc_lob;
      5'b01100:
        casez_tmp_322 = ldq_12_bits_uop_pc_lob;
      5'b01101:
        casez_tmp_322 = ldq_13_bits_uop_pc_lob;
      5'b01110:
        casez_tmp_322 = ldq_14_bits_uop_pc_lob;
      5'b01111:
        casez_tmp_322 = ldq_15_bits_uop_pc_lob;
      5'b10000:
        casez_tmp_322 = ldq_16_bits_uop_pc_lob;
      5'b10001:
        casez_tmp_322 = ldq_17_bits_uop_pc_lob;
      5'b10010:
        casez_tmp_322 = ldq_18_bits_uop_pc_lob;
      5'b10011:
        casez_tmp_322 = ldq_19_bits_uop_pc_lob;
      5'b10100:
        casez_tmp_322 = ldq_20_bits_uop_pc_lob;
      5'b10101:
        casez_tmp_322 = ldq_21_bits_uop_pc_lob;
      5'b10110:
        casez_tmp_322 = ldq_22_bits_uop_pc_lob;
      5'b10111:
        casez_tmp_322 = ldq_23_bits_uop_pc_lob;
      5'b11000:
        casez_tmp_322 = ldq_24_bits_uop_pc_lob;
      5'b11001:
        casez_tmp_322 = ldq_25_bits_uop_pc_lob;
      5'b11010:
        casez_tmp_322 = ldq_26_bits_uop_pc_lob;
      5'b11011:
        casez_tmp_322 = ldq_27_bits_uop_pc_lob;
      5'b11100:
        casez_tmp_322 = ldq_28_bits_uop_pc_lob;
      5'b11101:
        casez_tmp_322 = ldq_29_bits_uop_pc_lob;
      5'b11110:
        casez_tmp_322 = ldq_30_bits_uop_pc_lob;
      default:
        casez_tmp_322 = ldq_31_bits_uop_pc_lob;
    endcase
  end // always @(*)
  reg         casez_tmp_323;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_323 = ldq_0_bits_uop_taken;
      5'b00001:
        casez_tmp_323 = ldq_1_bits_uop_taken;
      5'b00010:
        casez_tmp_323 = ldq_2_bits_uop_taken;
      5'b00011:
        casez_tmp_323 = ldq_3_bits_uop_taken;
      5'b00100:
        casez_tmp_323 = ldq_4_bits_uop_taken;
      5'b00101:
        casez_tmp_323 = ldq_5_bits_uop_taken;
      5'b00110:
        casez_tmp_323 = ldq_6_bits_uop_taken;
      5'b00111:
        casez_tmp_323 = ldq_7_bits_uop_taken;
      5'b01000:
        casez_tmp_323 = ldq_8_bits_uop_taken;
      5'b01001:
        casez_tmp_323 = ldq_9_bits_uop_taken;
      5'b01010:
        casez_tmp_323 = ldq_10_bits_uop_taken;
      5'b01011:
        casez_tmp_323 = ldq_11_bits_uop_taken;
      5'b01100:
        casez_tmp_323 = ldq_12_bits_uop_taken;
      5'b01101:
        casez_tmp_323 = ldq_13_bits_uop_taken;
      5'b01110:
        casez_tmp_323 = ldq_14_bits_uop_taken;
      5'b01111:
        casez_tmp_323 = ldq_15_bits_uop_taken;
      5'b10000:
        casez_tmp_323 = ldq_16_bits_uop_taken;
      5'b10001:
        casez_tmp_323 = ldq_17_bits_uop_taken;
      5'b10010:
        casez_tmp_323 = ldq_18_bits_uop_taken;
      5'b10011:
        casez_tmp_323 = ldq_19_bits_uop_taken;
      5'b10100:
        casez_tmp_323 = ldq_20_bits_uop_taken;
      5'b10101:
        casez_tmp_323 = ldq_21_bits_uop_taken;
      5'b10110:
        casez_tmp_323 = ldq_22_bits_uop_taken;
      5'b10111:
        casez_tmp_323 = ldq_23_bits_uop_taken;
      5'b11000:
        casez_tmp_323 = ldq_24_bits_uop_taken;
      5'b11001:
        casez_tmp_323 = ldq_25_bits_uop_taken;
      5'b11010:
        casez_tmp_323 = ldq_26_bits_uop_taken;
      5'b11011:
        casez_tmp_323 = ldq_27_bits_uop_taken;
      5'b11100:
        casez_tmp_323 = ldq_28_bits_uop_taken;
      5'b11101:
        casez_tmp_323 = ldq_29_bits_uop_taken;
      5'b11110:
        casez_tmp_323 = ldq_30_bits_uop_taken;
      default:
        casez_tmp_323 = ldq_31_bits_uop_taken;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_324;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_324 = ldq_0_bits_uop_imm_packed;
      5'b00001:
        casez_tmp_324 = ldq_1_bits_uop_imm_packed;
      5'b00010:
        casez_tmp_324 = ldq_2_bits_uop_imm_packed;
      5'b00011:
        casez_tmp_324 = ldq_3_bits_uop_imm_packed;
      5'b00100:
        casez_tmp_324 = ldq_4_bits_uop_imm_packed;
      5'b00101:
        casez_tmp_324 = ldq_5_bits_uop_imm_packed;
      5'b00110:
        casez_tmp_324 = ldq_6_bits_uop_imm_packed;
      5'b00111:
        casez_tmp_324 = ldq_7_bits_uop_imm_packed;
      5'b01000:
        casez_tmp_324 = ldq_8_bits_uop_imm_packed;
      5'b01001:
        casez_tmp_324 = ldq_9_bits_uop_imm_packed;
      5'b01010:
        casez_tmp_324 = ldq_10_bits_uop_imm_packed;
      5'b01011:
        casez_tmp_324 = ldq_11_bits_uop_imm_packed;
      5'b01100:
        casez_tmp_324 = ldq_12_bits_uop_imm_packed;
      5'b01101:
        casez_tmp_324 = ldq_13_bits_uop_imm_packed;
      5'b01110:
        casez_tmp_324 = ldq_14_bits_uop_imm_packed;
      5'b01111:
        casez_tmp_324 = ldq_15_bits_uop_imm_packed;
      5'b10000:
        casez_tmp_324 = ldq_16_bits_uop_imm_packed;
      5'b10001:
        casez_tmp_324 = ldq_17_bits_uop_imm_packed;
      5'b10010:
        casez_tmp_324 = ldq_18_bits_uop_imm_packed;
      5'b10011:
        casez_tmp_324 = ldq_19_bits_uop_imm_packed;
      5'b10100:
        casez_tmp_324 = ldq_20_bits_uop_imm_packed;
      5'b10101:
        casez_tmp_324 = ldq_21_bits_uop_imm_packed;
      5'b10110:
        casez_tmp_324 = ldq_22_bits_uop_imm_packed;
      5'b10111:
        casez_tmp_324 = ldq_23_bits_uop_imm_packed;
      5'b11000:
        casez_tmp_324 = ldq_24_bits_uop_imm_packed;
      5'b11001:
        casez_tmp_324 = ldq_25_bits_uop_imm_packed;
      5'b11010:
        casez_tmp_324 = ldq_26_bits_uop_imm_packed;
      5'b11011:
        casez_tmp_324 = ldq_27_bits_uop_imm_packed;
      5'b11100:
        casez_tmp_324 = ldq_28_bits_uop_imm_packed;
      5'b11101:
        casez_tmp_324 = ldq_29_bits_uop_imm_packed;
      5'b11110:
        casez_tmp_324 = ldq_30_bits_uop_imm_packed;
      default:
        casez_tmp_324 = ldq_31_bits_uop_imm_packed;
    endcase
  end // always @(*)
  reg  [11:0] casez_tmp_325;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_325 = ldq_0_bits_uop_csr_addr;
      5'b00001:
        casez_tmp_325 = ldq_1_bits_uop_csr_addr;
      5'b00010:
        casez_tmp_325 = ldq_2_bits_uop_csr_addr;
      5'b00011:
        casez_tmp_325 = ldq_3_bits_uop_csr_addr;
      5'b00100:
        casez_tmp_325 = ldq_4_bits_uop_csr_addr;
      5'b00101:
        casez_tmp_325 = ldq_5_bits_uop_csr_addr;
      5'b00110:
        casez_tmp_325 = ldq_6_bits_uop_csr_addr;
      5'b00111:
        casez_tmp_325 = ldq_7_bits_uop_csr_addr;
      5'b01000:
        casez_tmp_325 = ldq_8_bits_uop_csr_addr;
      5'b01001:
        casez_tmp_325 = ldq_9_bits_uop_csr_addr;
      5'b01010:
        casez_tmp_325 = ldq_10_bits_uop_csr_addr;
      5'b01011:
        casez_tmp_325 = ldq_11_bits_uop_csr_addr;
      5'b01100:
        casez_tmp_325 = ldq_12_bits_uop_csr_addr;
      5'b01101:
        casez_tmp_325 = ldq_13_bits_uop_csr_addr;
      5'b01110:
        casez_tmp_325 = ldq_14_bits_uop_csr_addr;
      5'b01111:
        casez_tmp_325 = ldq_15_bits_uop_csr_addr;
      5'b10000:
        casez_tmp_325 = ldq_16_bits_uop_csr_addr;
      5'b10001:
        casez_tmp_325 = ldq_17_bits_uop_csr_addr;
      5'b10010:
        casez_tmp_325 = ldq_18_bits_uop_csr_addr;
      5'b10011:
        casez_tmp_325 = ldq_19_bits_uop_csr_addr;
      5'b10100:
        casez_tmp_325 = ldq_20_bits_uop_csr_addr;
      5'b10101:
        casez_tmp_325 = ldq_21_bits_uop_csr_addr;
      5'b10110:
        casez_tmp_325 = ldq_22_bits_uop_csr_addr;
      5'b10111:
        casez_tmp_325 = ldq_23_bits_uop_csr_addr;
      5'b11000:
        casez_tmp_325 = ldq_24_bits_uop_csr_addr;
      5'b11001:
        casez_tmp_325 = ldq_25_bits_uop_csr_addr;
      5'b11010:
        casez_tmp_325 = ldq_26_bits_uop_csr_addr;
      5'b11011:
        casez_tmp_325 = ldq_27_bits_uop_csr_addr;
      5'b11100:
        casez_tmp_325 = ldq_28_bits_uop_csr_addr;
      5'b11101:
        casez_tmp_325 = ldq_29_bits_uop_csr_addr;
      5'b11110:
        casez_tmp_325 = ldq_30_bits_uop_csr_addr;
      default:
        casez_tmp_325 = ldq_31_bits_uop_csr_addr;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_326;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_326 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_326 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_326 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_326 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_326 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_326 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_326 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_326 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_326 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_326 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_326 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_326 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_326 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_326 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_326 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_326 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_326 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_326 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_326 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_326 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_326 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_326 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_326 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_326 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_326 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_326 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_326 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_326 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_326 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_326 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_326 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_326 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_327;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_327 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_327 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_327 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_327 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_327 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_327 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_327 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_327 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_327 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_327 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_327 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_327 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_327 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_327 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_327 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_327 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_327 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_327 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_327 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_327 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_327 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_327 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_327 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_327 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_327 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_327 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_327 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_327 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_327 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_327 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_327 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_327 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_328;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_328 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_328 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_328 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_328 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_328 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_328 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_328 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_328 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_328 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_328 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_328 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_328 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_328 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_328 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_328 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_328 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_328 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_328 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_328 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_328 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_328 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_328 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_328 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_328 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_328 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_328 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_328 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_328 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_328 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_328 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_328 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_328 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_329;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_329 = ldq_0_bits_uop_rxq_idx;
      5'b00001:
        casez_tmp_329 = ldq_1_bits_uop_rxq_idx;
      5'b00010:
        casez_tmp_329 = ldq_2_bits_uop_rxq_idx;
      5'b00011:
        casez_tmp_329 = ldq_3_bits_uop_rxq_idx;
      5'b00100:
        casez_tmp_329 = ldq_4_bits_uop_rxq_idx;
      5'b00101:
        casez_tmp_329 = ldq_5_bits_uop_rxq_idx;
      5'b00110:
        casez_tmp_329 = ldq_6_bits_uop_rxq_idx;
      5'b00111:
        casez_tmp_329 = ldq_7_bits_uop_rxq_idx;
      5'b01000:
        casez_tmp_329 = ldq_8_bits_uop_rxq_idx;
      5'b01001:
        casez_tmp_329 = ldq_9_bits_uop_rxq_idx;
      5'b01010:
        casez_tmp_329 = ldq_10_bits_uop_rxq_idx;
      5'b01011:
        casez_tmp_329 = ldq_11_bits_uop_rxq_idx;
      5'b01100:
        casez_tmp_329 = ldq_12_bits_uop_rxq_idx;
      5'b01101:
        casez_tmp_329 = ldq_13_bits_uop_rxq_idx;
      5'b01110:
        casez_tmp_329 = ldq_14_bits_uop_rxq_idx;
      5'b01111:
        casez_tmp_329 = ldq_15_bits_uop_rxq_idx;
      5'b10000:
        casez_tmp_329 = ldq_16_bits_uop_rxq_idx;
      5'b10001:
        casez_tmp_329 = ldq_17_bits_uop_rxq_idx;
      5'b10010:
        casez_tmp_329 = ldq_18_bits_uop_rxq_idx;
      5'b10011:
        casez_tmp_329 = ldq_19_bits_uop_rxq_idx;
      5'b10100:
        casez_tmp_329 = ldq_20_bits_uop_rxq_idx;
      5'b10101:
        casez_tmp_329 = ldq_21_bits_uop_rxq_idx;
      5'b10110:
        casez_tmp_329 = ldq_22_bits_uop_rxq_idx;
      5'b10111:
        casez_tmp_329 = ldq_23_bits_uop_rxq_idx;
      5'b11000:
        casez_tmp_329 = ldq_24_bits_uop_rxq_idx;
      5'b11001:
        casez_tmp_329 = ldq_25_bits_uop_rxq_idx;
      5'b11010:
        casez_tmp_329 = ldq_26_bits_uop_rxq_idx;
      5'b11011:
        casez_tmp_329 = ldq_27_bits_uop_rxq_idx;
      5'b11100:
        casez_tmp_329 = ldq_28_bits_uop_rxq_idx;
      5'b11101:
        casez_tmp_329 = ldq_29_bits_uop_rxq_idx;
      5'b11110:
        casez_tmp_329 = ldq_30_bits_uop_rxq_idx;
      default:
        casez_tmp_329 = ldq_31_bits_uop_rxq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_330;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_330 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_330 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_330 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_330 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_330 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_330 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_330 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_330 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_330 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_330 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_330 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_330 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_330 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_330 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_330 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_330 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_330 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_330 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_330 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_330 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_330 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_330 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_330 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_330 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_330 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_330 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_330 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_330 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_330 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_330 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_330 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_330 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_331;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_331 = ldq_0_bits_uop_prs1;
      5'b00001:
        casez_tmp_331 = ldq_1_bits_uop_prs1;
      5'b00010:
        casez_tmp_331 = ldq_2_bits_uop_prs1;
      5'b00011:
        casez_tmp_331 = ldq_3_bits_uop_prs1;
      5'b00100:
        casez_tmp_331 = ldq_4_bits_uop_prs1;
      5'b00101:
        casez_tmp_331 = ldq_5_bits_uop_prs1;
      5'b00110:
        casez_tmp_331 = ldq_6_bits_uop_prs1;
      5'b00111:
        casez_tmp_331 = ldq_7_bits_uop_prs1;
      5'b01000:
        casez_tmp_331 = ldq_8_bits_uop_prs1;
      5'b01001:
        casez_tmp_331 = ldq_9_bits_uop_prs1;
      5'b01010:
        casez_tmp_331 = ldq_10_bits_uop_prs1;
      5'b01011:
        casez_tmp_331 = ldq_11_bits_uop_prs1;
      5'b01100:
        casez_tmp_331 = ldq_12_bits_uop_prs1;
      5'b01101:
        casez_tmp_331 = ldq_13_bits_uop_prs1;
      5'b01110:
        casez_tmp_331 = ldq_14_bits_uop_prs1;
      5'b01111:
        casez_tmp_331 = ldq_15_bits_uop_prs1;
      5'b10000:
        casez_tmp_331 = ldq_16_bits_uop_prs1;
      5'b10001:
        casez_tmp_331 = ldq_17_bits_uop_prs1;
      5'b10010:
        casez_tmp_331 = ldq_18_bits_uop_prs1;
      5'b10011:
        casez_tmp_331 = ldq_19_bits_uop_prs1;
      5'b10100:
        casez_tmp_331 = ldq_20_bits_uop_prs1;
      5'b10101:
        casez_tmp_331 = ldq_21_bits_uop_prs1;
      5'b10110:
        casez_tmp_331 = ldq_22_bits_uop_prs1;
      5'b10111:
        casez_tmp_331 = ldq_23_bits_uop_prs1;
      5'b11000:
        casez_tmp_331 = ldq_24_bits_uop_prs1;
      5'b11001:
        casez_tmp_331 = ldq_25_bits_uop_prs1;
      5'b11010:
        casez_tmp_331 = ldq_26_bits_uop_prs1;
      5'b11011:
        casez_tmp_331 = ldq_27_bits_uop_prs1;
      5'b11100:
        casez_tmp_331 = ldq_28_bits_uop_prs1;
      5'b11101:
        casez_tmp_331 = ldq_29_bits_uop_prs1;
      5'b11110:
        casez_tmp_331 = ldq_30_bits_uop_prs1;
      default:
        casez_tmp_331 = ldq_31_bits_uop_prs1;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_332;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_332 = ldq_0_bits_uop_prs2;
      5'b00001:
        casez_tmp_332 = ldq_1_bits_uop_prs2;
      5'b00010:
        casez_tmp_332 = ldq_2_bits_uop_prs2;
      5'b00011:
        casez_tmp_332 = ldq_3_bits_uop_prs2;
      5'b00100:
        casez_tmp_332 = ldq_4_bits_uop_prs2;
      5'b00101:
        casez_tmp_332 = ldq_5_bits_uop_prs2;
      5'b00110:
        casez_tmp_332 = ldq_6_bits_uop_prs2;
      5'b00111:
        casez_tmp_332 = ldq_7_bits_uop_prs2;
      5'b01000:
        casez_tmp_332 = ldq_8_bits_uop_prs2;
      5'b01001:
        casez_tmp_332 = ldq_9_bits_uop_prs2;
      5'b01010:
        casez_tmp_332 = ldq_10_bits_uop_prs2;
      5'b01011:
        casez_tmp_332 = ldq_11_bits_uop_prs2;
      5'b01100:
        casez_tmp_332 = ldq_12_bits_uop_prs2;
      5'b01101:
        casez_tmp_332 = ldq_13_bits_uop_prs2;
      5'b01110:
        casez_tmp_332 = ldq_14_bits_uop_prs2;
      5'b01111:
        casez_tmp_332 = ldq_15_bits_uop_prs2;
      5'b10000:
        casez_tmp_332 = ldq_16_bits_uop_prs2;
      5'b10001:
        casez_tmp_332 = ldq_17_bits_uop_prs2;
      5'b10010:
        casez_tmp_332 = ldq_18_bits_uop_prs2;
      5'b10011:
        casez_tmp_332 = ldq_19_bits_uop_prs2;
      5'b10100:
        casez_tmp_332 = ldq_20_bits_uop_prs2;
      5'b10101:
        casez_tmp_332 = ldq_21_bits_uop_prs2;
      5'b10110:
        casez_tmp_332 = ldq_22_bits_uop_prs2;
      5'b10111:
        casez_tmp_332 = ldq_23_bits_uop_prs2;
      5'b11000:
        casez_tmp_332 = ldq_24_bits_uop_prs2;
      5'b11001:
        casez_tmp_332 = ldq_25_bits_uop_prs2;
      5'b11010:
        casez_tmp_332 = ldq_26_bits_uop_prs2;
      5'b11011:
        casez_tmp_332 = ldq_27_bits_uop_prs2;
      5'b11100:
        casez_tmp_332 = ldq_28_bits_uop_prs2;
      5'b11101:
        casez_tmp_332 = ldq_29_bits_uop_prs2;
      5'b11110:
        casez_tmp_332 = ldq_30_bits_uop_prs2;
      default:
        casez_tmp_332 = ldq_31_bits_uop_prs2;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_333;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_333 = ldq_0_bits_uop_prs3;
      5'b00001:
        casez_tmp_333 = ldq_1_bits_uop_prs3;
      5'b00010:
        casez_tmp_333 = ldq_2_bits_uop_prs3;
      5'b00011:
        casez_tmp_333 = ldq_3_bits_uop_prs3;
      5'b00100:
        casez_tmp_333 = ldq_4_bits_uop_prs3;
      5'b00101:
        casez_tmp_333 = ldq_5_bits_uop_prs3;
      5'b00110:
        casez_tmp_333 = ldq_6_bits_uop_prs3;
      5'b00111:
        casez_tmp_333 = ldq_7_bits_uop_prs3;
      5'b01000:
        casez_tmp_333 = ldq_8_bits_uop_prs3;
      5'b01001:
        casez_tmp_333 = ldq_9_bits_uop_prs3;
      5'b01010:
        casez_tmp_333 = ldq_10_bits_uop_prs3;
      5'b01011:
        casez_tmp_333 = ldq_11_bits_uop_prs3;
      5'b01100:
        casez_tmp_333 = ldq_12_bits_uop_prs3;
      5'b01101:
        casez_tmp_333 = ldq_13_bits_uop_prs3;
      5'b01110:
        casez_tmp_333 = ldq_14_bits_uop_prs3;
      5'b01111:
        casez_tmp_333 = ldq_15_bits_uop_prs3;
      5'b10000:
        casez_tmp_333 = ldq_16_bits_uop_prs3;
      5'b10001:
        casez_tmp_333 = ldq_17_bits_uop_prs3;
      5'b10010:
        casez_tmp_333 = ldq_18_bits_uop_prs3;
      5'b10011:
        casez_tmp_333 = ldq_19_bits_uop_prs3;
      5'b10100:
        casez_tmp_333 = ldq_20_bits_uop_prs3;
      5'b10101:
        casez_tmp_333 = ldq_21_bits_uop_prs3;
      5'b10110:
        casez_tmp_333 = ldq_22_bits_uop_prs3;
      5'b10111:
        casez_tmp_333 = ldq_23_bits_uop_prs3;
      5'b11000:
        casez_tmp_333 = ldq_24_bits_uop_prs3;
      5'b11001:
        casez_tmp_333 = ldq_25_bits_uop_prs3;
      5'b11010:
        casez_tmp_333 = ldq_26_bits_uop_prs3;
      5'b11011:
        casez_tmp_333 = ldq_27_bits_uop_prs3;
      5'b11100:
        casez_tmp_333 = ldq_28_bits_uop_prs3;
      5'b11101:
        casez_tmp_333 = ldq_29_bits_uop_prs3;
      5'b11110:
        casez_tmp_333 = ldq_30_bits_uop_prs3;
      default:
        casez_tmp_333 = ldq_31_bits_uop_prs3;
    endcase
  end // always @(*)
  reg         casez_tmp_334;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_334 = ldq_0_bits_uop_prs1_busy;
      5'b00001:
        casez_tmp_334 = ldq_1_bits_uop_prs1_busy;
      5'b00010:
        casez_tmp_334 = ldq_2_bits_uop_prs1_busy;
      5'b00011:
        casez_tmp_334 = ldq_3_bits_uop_prs1_busy;
      5'b00100:
        casez_tmp_334 = ldq_4_bits_uop_prs1_busy;
      5'b00101:
        casez_tmp_334 = ldq_5_bits_uop_prs1_busy;
      5'b00110:
        casez_tmp_334 = ldq_6_bits_uop_prs1_busy;
      5'b00111:
        casez_tmp_334 = ldq_7_bits_uop_prs1_busy;
      5'b01000:
        casez_tmp_334 = ldq_8_bits_uop_prs1_busy;
      5'b01001:
        casez_tmp_334 = ldq_9_bits_uop_prs1_busy;
      5'b01010:
        casez_tmp_334 = ldq_10_bits_uop_prs1_busy;
      5'b01011:
        casez_tmp_334 = ldq_11_bits_uop_prs1_busy;
      5'b01100:
        casez_tmp_334 = ldq_12_bits_uop_prs1_busy;
      5'b01101:
        casez_tmp_334 = ldq_13_bits_uop_prs1_busy;
      5'b01110:
        casez_tmp_334 = ldq_14_bits_uop_prs1_busy;
      5'b01111:
        casez_tmp_334 = ldq_15_bits_uop_prs1_busy;
      5'b10000:
        casez_tmp_334 = ldq_16_bits_uop_prs1_busy;
      5'b10001:
        casez_tmp_334 = ldq_17_bits_uop_prs1_busy;
      5'b10010:
        casez_tmp_334 = ldq_18_bits_uop_prs1_busy;
      5'b10011:
        casez_tmp_334 = ldq_19_bits_uop_prs1_busy;
      5'b10100:
        casez_tmp_334 = ldq_20_bits_uop_prs1_busy;
      5'b10101:
        casez_tmp_334 = ldq_21_bits_uop_prs1_busy;
      5'b10110:
        casez_tmp_334 = ldq_22_bits_uop_prs1_busy;
      5'b10111:
        casez_tmp_334 = ldq_23_bits_uop_prs1_busy;
      5'b11000:
        casez_tmp_334 = ldq_24_bits_uop_prs1_busy;
      5'b11001:
        casez_tmp_334 = ldq_25_bits_uop_prs1_busy;
      5'b11010:
        casez_tmp_334 = ldq_26_bits_uop_prs1_busy;
      5'b11011:
        casez_tmp_334 = ldq_27_bits_uop_prs1_busy;
      5'b11100:
        casez_tmp_334 = ldq_28_bits_uop_prs1_busy;
      5'b11101:
        casez_tmp_334 = ldq_29_bits_uop_prs1_busy;
      5'b11110:
        casez_tmp_334 = ldq_30_bits_uop_prs1_busy;
      default:
        casez_tmp_334 = ldq_31_bits_uop_prs1_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_335;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_335 = ldq_0_bits_uop_prs2_busy;
      5'b00001:
        casez_tmp_335 = ldq_1_bits_uop_prs2_busy;
      5'b00010:
        casez_tmp_335 = ldq_2_bits_uop_prs2_busy;
      5'b00011:
        casez_tmp_335 = ldq_3_bits_uop_prs2_busy;
      5'b00100:
        casez_tmp_335 = ldq_4_bits_uop_prs2_busy;
      5'b00101:
        casez_tmp_335 = ldq_5_bits_uop_prs2_busy;
      5'b00110:
        casez_tmp_335 = ldq_6_bits_uop_prs2_busy;
      5'b00111:
        casez_tmp_335 = ldq_7_bits_uop_prs2_busy;
      5'b01000:
        casez_tmp_335 = ldq_8_bits_uop_prs2_busy;
      5'b01001:
        casez_tmp_335 = ldq_9_bits_uop_prs2_busy;
      5'b01010:
        casez_tmp_335 = ldq_10_bits_uop_prs2_busy;
      5'b01011:
        casez_tmp_335 = ldq_11_bits_uop_prs2_busy;
      5'b01100:
        casez_tmp_335 = ldq_12_bits_uop_prs2_busy;
      5'b01101:
        casez_tmp_335 = ldq_13_bits_uop_prs2_busy;
      5'b01110:
        casez_tmp_335 = ldq_14_bits_uop_prs2_busy;
      5'b01111:
        casez_tmp_335 = ldq_15_bits_uop_prs2_busy;
      5'b10000:
        casez_tmp_335 = ldq_16_bits_uop_prs2_busy;
      5'b10001:
        casez_tmp_335 = ldq_17_bits_uop_prs2_busy;
      5'b10010:
        casez_tmp_335 = ldq_18_bits_uop_prs2_busy;
      5'b10011:
        casez_tmp_335 = ldq_19_bits_uop_prs2_busy;
      5'b10100:
        casez_tmp_335 = ldq_20_bits_uop_prs2_busy;
      5'b10101:
        casez_tmp_335 = ldq_21_bits_uop_prs2_busy;
      5'b10110:
        casez_tmp_335 = ldq_22_bits_uop_prs2_busy;
      5'b10111:
        casez_tmp_335 = ldq_23_bits_uop_prs2_busy;
      5'b11000:
        casez_tmp_335 = ldq_24_bits_uop_prs2_busy;
      5'b11001:
        casez_tmp_335 = ldq_25_bits_uop_prs2_busy;
      5'b11010:
        casez_tmp_335 = ldq_26_bits_uop_prs2_busy;
      5'b11011:
        casez_tmp_335 = ldq_27_bits_uop_prs2_busy;
      5'b11100:
        casez_tmp_335 = ldq_28_bits_uop_prs2_busy;
      5'b11101:
        casez_tmp_335 = ldq_29_bits_uop_prs2_busy;
      5'b11110:
        casez_tmp_335 = ldq_30_bits_uop_prs2_busy;
      default:
        casez_tmp_335 = ldq_31_bits_uop_prs2_busy;
    endcase
  end // always @(*)
  reg         casez_tmp_336;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_336 = ldq_0_bits_uop_prs3_busy;
      5'b00001:
        casez_tmp_336 = ldq_1_bits_uop_prs3_busy;
      5'b00010:
        casez_tmp_336 = ldq_2_bits_uop_prs3_busy;
      5'b00011:
        casez_tmp_336 = ldq_3_bits_uop_prs3_busy;
      5'b00100:
        casez_tmp_336 = ldq_4_bits_uop_prs3_busy;
      5'b00101:
        casez_tmp_336 = ldq_5_bits_uop_prs3_busy;
      5'b00110:
        casez_tmp_336 = ldq_6_bits_uop_prs3_busy;
      5'b00111:
        casez_tmp_336 = ldq_7_bits_uop_prs3_busy;
      5'b01000:
        casez_tmp_336 = ldq_8_bits_uop_prs3_busy;
      5'b01001:
        casez_tmp_336 = ldq_9_bits_uop_prs3_busy;
      5'b01010:
        casez_tmp_336 = ldq_10_bits_uop_prs3_busy;
      5'b01011:
        casez_tmp_336 = ldq_11_bits_uop_prs3_busy;
      5'b01100:
        casez_tmp_336 = ldq_12_bits_uop_prs3_busy;
      5'b01101:
        casez_tmp_336 = ldq_13_bits_uop_prs3_busy;
      5'b01110:
        casez_tmp_336 = ldq_14_bits_uop_prs3_busy;
      5'b01111:
        casez_tmp_336 = ldq_15_bits_uop_prs3_busy;
      5'b10000:
        casez_tmp_336 = ldq_16_bits_uop_prs3_busy;
      5'b10001:
        casez_tmp_336 = ldq_17_bits_uop_prs3_busy;
      5'b10010:
        casez_tmp_336 = ldq_18_bits_uop_prs3_busy;
      5'b10011:
        casez_tmp_336 = ldq_19_bits_uop_prs3_busy;
      5'b10100:
        casez_tmp_336 = ldq_20_bits_uop_prs3_busy;
      5'b10101:
        casez_tmp_336 = ldq_21_bits_uop_prs3_busy;
      5'b10110:
        casez_tmp_336 = ldq_22_bits_uop_prs3_busy;
      5'b10111:
        casez_tmp_336 = ldq_23_bits_uop_prs3_busy;
      5'b11000:
        casez_tmp_336 = ldq_24_bits_uop_prs3_busy;
      5'b11001:
        casez_tmp_336 = ldq_25_bits_uop_prs3_busy;
      5'b11010:
        casez_tmp_336 = ldq_26_bits_uop_prs3_busy;
      5'b11011:
        casez_tmp_336 = ldq_27_bits_uop_prs3_busy;
      5'b11100:
        casez_tmp_336 = ldq_28_bits_uop_prs3_busy;
      5'b11101:
        casez_tmp_336 = ldq_29_bits_uop_prs3_busy;
      5'b11110:
        casez_tmp_336 = ldq_30_bits_uop_prs3_busy;
      default:
        casez_tmp_336 = ldq_31_bits_uop_prs3_busy;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_337;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_337 = ldq_0_bits_uop_stale_pdst;
      5'b00001:
        casez_tmp_337 = ldq_1_bits_uop_stale_pdst;
      5'b00010:
        casez_tmp_337 = ldq_2_bits_uop_stale_pdst;
      5'b00011:
        casez_tmp_337 = ldq_3_bits_uop_stale_pdst;
      5'b00100:
        casez_tmp_337 = ldq_4_bits_uop_stale_pdst;
      5'b00101:
        casez_tmp_337 = ldq_5_bits_uop_stale_pdst;
      5'b00110:
        casez_tmp_337 = ldq_6_bits_uop_stale_pdst;
      5'b00111:
        casez_tmp_337 = ldq_7_bits_uop_stale_pdst;
      5'b01000:
        casez_tmp_337 = ldq_8_bits_uop_stale_pdst;
      5'b01001:
        casez_tmp_337 = ldq_9_bits_uop_stale_pdst;
      5'b01010:
        casez_tmp_337 = ldq_10_bits_uop_stale_pdst;
      5'b01011:
        casez_tmp_337 = ldq_11_bits_uop_stale_pdst;
      5'b01100:
        casez_tmp_337 = ldq_12_bits_uop_stale_pdst;
      5'b01101:
        casez_tmp_337 = ldq_13_bits_uop_stale_pdst;
      5'b01110:
        casez_tmp_337 = ldq_14_bits_uop_stale_pdst;
      5'b01111:
        casez_tmp_337 = ldq_15_bits_uop_stale_pdst;
      5'b10000:
        casez_tmp_337 = ldq_16_bits_uop_stale_pdst;
      5'b10001:
        casez_tmp_337 = ldq_17_bits_uop_stale_pdst;
      5'b10010:
        casez_tmp_337 = ldq_18_bits_uop_stale_pdst;
      5'b10011:
        casez_tmp_337 = ldq_19_bits_uop_stale_pdst;
      5'b10100:
        casez_tmp_337 = ldq_20_bits_uop_stale_pdst;
      5'b10101:
        casez_tmp_337 = ldq_21_bits_uop_stale_pdst;
      5'b10110:
        casez_tmp_337 = ldq_22_bits_uop_stale_pdst;
      5'b10111:
        casez_tmp_337 = ldq_23_bits_uop_stale_pdst;
      5'b11000:
        casez_tmp_337 = ldq_24_bits_uop_stale_pdst;
      5'b11001:
        casez_tmp_337 = ldq_25_bits_uop_stale_pdst;
      5'b11010:
        casez_tmp_337 = ldq_26_bits_uop_stale_pdst;
      5'b11011:
        casez_tmp_337 = ldq_27_bits_uop_stale_pdst;
      5'b11100:
        casez_tmp_337 = ldq_28_bits_uop_stale_pdst;
      5'b11101:
        casez_tmp_337 = ldq_29_bits_uop_stale_pdst;
      5'b11110:
        casez_tmp_337 = ldq_30_bits_uop_stale_pdst;
      default:
        casez_tmp_337 = ldq_31_bits_uop_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_338;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_338 = ldq_0_bits_uop_exception;
      5'b00001:
        casez_tmp_338 = ldq_1_bits_uop_exception;
      5'b00010:
        casez_tmp_338 = ldq_2_bits_uop_exception;
      5'b00011:
        casez_tmp_338 = ldq_3_bits_uop_exception;
      5'b00100:
        casez_tmp_338 = ldq_4_bits_uop_exception;
      5'b00101:
        casez_tmp_338 = ldq_5_bits_uop_exception;
      5'b00110:
        casez_tmp_338 = ldq_6_bits_uop_exception;
      5'b00111:
        casez_tmp_338 = ldq_7_bits_uop_exception;
      5'b01000:
        casez_tmp_338 = ldq_8_bits_uop_exception;
      5'b01001:
        casez_tmp_338 = ldq_9_bits_uop_exception;
      5'b01010:
        casez_tmp_338 = ldq_10_bits_uop_exception;
      5'b01011:
        casez_tmp_338 = ldq_11_bits_uop_exception;
      5'b01100:
        casez_tmp_338 = ldq_12_bits_uop_exception;
      5'b01101:
        casez_tmp_338 = ldq_13_bits_uop_exception;
      5'b01110:
        casez_tmp_338 = ldq_14_bits_uop_exception;
      5'b01111:
        casez_tmp_338 = ldq_15_bits_uop_exception;
      5'b10000:
        casez_tmp_338 = ldq_16_bits_uop_exception;
      5'b10001:
        casez_tmp_338 = ldq_17_bits_uop_exception;
      5'b10010:
        casez_tmp_338 = ldq_18_bits_uop_exception;
      5'b10011:
        casez_tmp_338 = ldq_19_bits_uop_exception;
      5'b10100:
        casez_tmp_338 = ldq_20_bits_uop_exception;
      5'b10101:
        casez_tmp_338 = ldq_21_bits_uop_exception;
      5'b10110:
        casez_tmp_338 = ldq_22_bits_uop_exception;
      5'b10111:
        casez_tmp_338 = ldq_23_bits_uop_exception;
      5'b11000:
        casez_tmp_338 = ldq_24_bits_uop_exception;
      5'b11001:
        casez_tmp_338 = ldq_25_bits_uop_exception;
      5'b11010:
        casez_tmp_338 = ldq_26_bits_uop_exception;
      5'b11011:
        casez_tmp_338 = ldq_27_bits_uop_exception;
      5'b11100:
        casez_tmp_338 = ldq_28_bits_uop_exception;
      5'b11101:
        casez_tmp_338 = ldq_29_bits_uop_exception;
      5'b11110:
        casez_tmp_338 = ldq_30_bits_uop_exception;
      default:
        casez_tmp_338 = ldq_31_bits_uop_exception;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_339;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_339 = ldq_0_bits_uop_exc_cause;
      5'b00001:
        casez_tmp_339 = ldq_1_bits_uop_exc_cause;
      5'b00010:
        casez_tmp_339 = ldq_2_bits_uop_exc_cause;
      5'b00011:
        casez_tmp_339 = ldq_3_bits_uop_exc_cause;
      5'b00100:
        casez_tmp_339 = ldq_4_bits_uop_exc_cause;
      5'b00101:
        casez_tmp_339 = ldq_5_bits_uop_exc_cause;
      5'b00110:
        casez_tmp_339 = ldq_6_bits_uop_exc_cause;
      5'b00111:
        casez_tmp_339 = ldq_7_bits_uop_exc_cause;
      5'b01000:
        casez_tmp_339 = ldq_8_bits_uop_exc_cause;
      5'b01001:
        casez_tmp_339 = ldq_9_bits_uop_exc_cause;
      5'b01010:
        casez_tmp_339 = ldq_10_bits_uop_exc_cause;
      5'b01011:
        casez_tmp_339 = ldq_11_bits_uop_exc_cause;
      5'b01100:
        casez_tmp_339 = ldq_12_bits_uop_exc_cause;
      5'b01101:
        casez_tmp_339 = ldq_13_bits_uop_exc_cause;
      5'b01110:
        casez_tmp_339 = ldq_14_bits_uop_exc_cause;
      5'b01111:
        casez_tmp_339 = ldq_15_bits_uop_exc_cause;
      5'b10000:
        casez_tmp_339 = ldq_16_bits_uop_exc_cause;
      5'b10001:
        casez_tmp_339 = ldq_17_bits_uop_exc_cause;
      5'b10010:
        casez_tmp_339 = ldq_18_bits_uop_exc_cause;
      5'b10011:
        casez_tmp_339 = ldq_19_bits_uop_exc_cause;
      5'b10100:
        casez_tmp_339 = ldq_20_bits_uop_exc_cause;
      5'b10101:
        casez_tmp_339 = ldq_21_bits_uop_exc_cause;
      5'b10110:
        casez_tmp_339 = ldq_22_bits_uop_exc_cause;
      5'b10111:
        casez_tmp_339 = ldq_23_bits_uop_exc_cause;
      5'b11000:
        casez_tmp_339 = ldq_24_bits_uop_exc_cause;
      5'b11001:
        casez_tmp_339 = ldq_25_bits_uop_exc_cause;
      5'b11010:
        casez_tmp_339 = ldq_26_bits_uop_exc_cause;
      5'b11011:
        casez_tmp_339 = ldq_27_bits_uop_exc_cause;
      5'b11100:
        casez_tmp_339 = ldq_28_bits_uop_exc_cause;
      5'b11101:
        casez_tmp_339 = ldq_29_bits_uop_exc_cause;
      5'b11110:
        casez_tmp_339 = ldq_30_bits_uop_exc_cause;
      default:
        casez_tmp_339 = ldq_31_bits_uop_exc_cause;
    endcase
  end // always @(*)
  reg         casez_tmp_340;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_340 = ldq_0_bits_uop_bypassable;
      5'b00001:
        casez_tmp_340 = ldq_1_bits_uop_bypassable;
      5'b00010:
        casez_tmp_340 = ldq_2_bits_uop_bypassable;
      5'b00011:
        casez_tmp_340 = ldq_3_bits_uop_bypassable;
      5'b00100:
        casez_tmp_340 = ldq_4_bits_uop_bypassable;
      5'b00101:
        casez_tmp_340 = ldq_5_bits_uop_bypassable;
      5'b00110:
        casez_tmp_340 = ldq_6_bits_uop_bypassable;
      5'b00111:
        casez_tmp_340 = ldq_7_bits_uop_bypassable;
      5'b01000:
        casez_tmp_340 = ldq_8_bits_uop_bypassable;
      5'b01001:
        casez_tmp_340 = ldq_9_bits_uop_bypassable;
      5'b01010:
        casez_tmp_340 = ldq_10_bits_uop_bypassable;
      5'b01011:
        casez_tmp_340 = ldq_11_bits_uop_bypassable;
      5'b01100:
        casez_tmp_340 = ldq_12_bits_uop_bypassable;
      5'b01101:
        casez_tmp_340 = ldq_13_bits_uop_bypassable;
      5'b01110:
        casez_tmp_340 = ldq_14_bits_uop_bypassable;
      5'b01111:
        casez_tmp_340 = ldq_15_bits_uop_bypassable;
      5'b10000:
        casez_tmp_340 = ldq_16_bits_uop_bypassable;
      5'b10001:
        casez_tmp_340 = ldq_17_bits_uop_bypassable;
      5'b10010:
        casez_tmp_340 = ldq_18_bits_uop_bypassable;
      5'b10011:
        casez_tmp_340 = ldq_19_bits_uop_bypassable;
      5'b10100:
        casez_tmp_340 = ldq_20_bits_uop_bypassable;
      5'b10101:
        casez_tmp_340 = ldq_21_bits_uop_bypassable;
      5'b10110:
        casez_tmp_340 = ldq_22_bits_uop_bypassable;
      5'b10111:
        casez_tmp_340 = ldq_23_bits_uop_bypassable;
      5'b11000:
        casez_tmp_340 = ldq_24_bits_uop_bypassable;
      5'b11001:
        casez_tmp_340 = ldq_25_bits_uop_bypassable;
      5'b11010:
        casez_tmp_340 = ldq_26_bits_uop_bypassable;
      5'b11011:
        casez_tmp_340 = ldq_27_bits_uop_bypassable;
      5'b11100:
        casez_tmp_340 = ldq_28_bits_uop_bypassable;
      5'b11101:
        casez_tmp_340 = ldq_29_bits_uop_bypassable;
      5'b11110:
        casez_tmp_340 = ldq_30_bits_uop_bypassable;
      default:
        casez_tmp_340 = ldq_31_bits_uop_bypassable;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_341;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_341 = ldq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_341 = ldq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_341 = ldq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_341 = ldq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_341 = ldq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_341 = ldq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_341 = ldq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_341 = ldq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_341 = ldq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_341 = ldq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_341 = ldq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_341 = ldq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_341 = ldq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_341 = ldq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_341 = ldq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_341 = ldq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_341 = ldq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_341 = ldq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_341 = ldq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_341 = ldq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_341 = ldq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_341 = ldq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_341 = ldq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_341 = ldq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_341 = ldq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_341 = ldq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_341 = ldq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_341 = ldq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_341 = ldq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_341 = ldq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_341 = ldq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_341 = ldq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_342;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_342 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_342 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_342 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_342 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_342 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_342 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_342 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_342 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_342 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_342 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_342 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_342 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_342 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_342 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_342 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_342 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_342 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_342 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_342 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_342 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_342 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_342 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_342 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_342 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_342 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_342 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_342 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_342 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_342 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_342 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_342 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_342 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_343;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_343 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_343 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_343 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_343 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_343 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_343 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_343 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_343 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_343 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_343 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_343 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_343 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_343 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_343 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_343 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_343 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_343 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_343 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_343 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_343 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_343 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_343 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_343 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_343 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_343 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_343 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_343 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_343 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_343 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_343 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_343 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_343 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  reg         casez_tmp_344;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_344 = ldq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_344 = ldq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_344 = ldq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_344 = ldq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_344 = ldq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_344 = ldq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_344 = ldq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_344 = ldq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_344 = ldq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_344 = ldq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_344 = ldq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_344 = ldq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_344 = ldq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_344 = ldq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_344 = ldq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_344 = ldq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_344 = ldq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_344 = ldq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_344 = ldq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_344 = ldq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_344 = ldq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_344 = ldq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_344 = ldq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_344 = ldq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_344 = ldq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_344 = ldq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_344 = ldq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_344 = ldq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_344 = ldq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_344 = ldq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_344 = ldq_30_bits_uop_is_fence;
      default:
        casez_tmp_344 = ldq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  reg         casez_tmp_345;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_345 = ldq_0_bits_uop_is_fencei;
      5'b00001:
        casez_tmp_345 = ldq_1_bits_uop_is_fencei;
      5'b00010:
        casez_tmp_345 = ldq_2_bits_uop_is_fencei;
      5'b00011:
        casez_tmp_345 = ldq_3_bits_uop_is_fencei;
      5'b00100:
        casez_tmp_345 = ldq_4_bits_uop_is_fencei;
      5'b00101:
        casez_tmp_345 = ldq_5_bits_uop_is_fencei;
      5'b00110:
        casez_tmp_345 = ldq_6_bits_uop_is_fencei;
      5'b00111:
        casez_tmp_345 = ldq_7_bits_uop_is_fencei;
      5'b01000:
        casez_tmp_345 = ldq_8_bits_uop_is_fencei;
      5'b01001:
        casez_tmp_345 = ldq_9_bits_uop_is_fencei;
      5'b01010:
        casez_tmp_345 = ldq_10_bits_uop_is_fencei;
      5'b01011:
        casez_tmp_345 = ldq_11_bits_uop_is_fencei;
      5'b01100:
        casez_tmp_345 = ldq_12_bits_uop_is_fencei;
      5'b01101:
        casez_tmp_345 = ldq_13_bits_uop_is_fencei;
      5'b01110:
        casez_tmp_345 = ldq_14_bits_uop_is_fencei;
      5'b01111:
        casez_tmp_345 = ldq_15_bits_uop_is_fencei;
      5'b10000:
        casez_tmp_345 = ldq_16_bits_uop_is_fencei;
      5'b10001:
        casez_tmp_345 = ldq_17_bits_uop_is_fencei;
      5'b10010:
        casez_tmp_345 = ldq_18_bits_uop_is_fencei;
      5'b10011:
        casez_tmp_345 = ldq_19_bits_uop_is_fencei;
      5'b10100:
        casez_tmp_345 = ldq_20_bits_uop_is_fencei;
      5'b10101:
        casez_tmp_345 = ldq_21_bits_uop_is_fencei;
      5'b10110:
        casez_tmp_345 = ldq_22_bits_uop_is_fencei;
      5'b10111:
        casez_tmp_345 = ldq_23_bits_uop_is_fencei;
      5'b11000:
        casez_tmp_345 = ldq_24_bits_uop_is_fencei;
      5'b11001:
        casez_tmp_345 = ldq_25_bits_uop_is_fencei;
      5'b11010:
        casez_tmp_345 = ldq_26_bits_uop_is_fencei;
      5'b11011:
        casez_tmp_345 = ldq_27_bits_uop_is_fencei;
      5'b11100:
        casez_tmp_345 = ldq_28_bits_uop_is_fencei;
      5'b11101:
        casez_tmp_345 = ldq_29_bits_uop_is_fencei;
      5'b11110:
        casez_tmp_345 = ldq_30_bits_uop_is_fencei;
      default:
        casez_tmp_345 = ldq_31_bits_uop_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_346;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_346 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_346 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_346 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_346 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_346 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_346 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_346 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_346 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_346 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_346 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_346 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_346 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_346 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_346 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_346 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_346 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_346 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_346 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_346 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_346 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_346 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_346 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_346 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_346 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_346 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_346 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_346 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_346 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_346 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_346 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_346 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_346 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_347;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_347 = ldq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_347 = ldq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_347 = ldq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_347 = ldq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_347 = ldq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_347 = ldq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_347 = ldq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_347 = ldq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_347 = ldq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_347 = ldq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_347 = ldq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_347 = ldq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_347 = ldq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_347 = ldq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_347 = ldq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_347 = ldq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_347 = ldq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_347 = ldq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_347 = ldq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_347 = ldq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_347 = ldq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_347 = ldq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_347 = ldq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_347 = ldq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_347 = ldq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_347 = ldq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_347 = ldq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_347 = ldq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_347 = ldq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_347 = ldq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_347 = ldq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_347 = ldq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_348;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_348 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_348 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_348 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_348 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_348 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_348 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_348 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_348 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_348 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_348 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_348 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_348 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_348 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_348 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_348 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_348 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_348 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_348 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_348 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_348 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_348 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_348 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_348 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_348 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_348 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_348 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_348 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_348 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_348 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_348 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_348 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_348 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_349;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_349 = ldq_0_bits_uop_is_sys_pc2epc;
      5'b00001:
        casez_tmp_349 = ldq_1_bits_uop_is_sys_pc2epc;
      5'b00010:
        casez_tmp_349 = ldq_2_bits_uop_is_sys_pc2epc;
      5'b00011:
        casez_tmp_349 = ldq_3_bits_uop_is_sys_pc2epc;
      5'b00100:
        casez_tmp_349 = ldq_4_bits_uop_is_sys_pc2epc;
      5'b00101:
        casez_tmp_349 = ldq_5_bits_uop_is_sys_pc2epc;
      5'b00110:
        casez_tmp_349 = ldq_6_bits_uop_is_sys_pc2epc;
      5'b00111:
        casez_tmp_349 = ldq_7_bits_uop_is_sys_pc2epc;
      5'b01000:
        casez_tmp_349 = ldq_8_bits_uop_is_sys_pc2epc;
      5'b01001:
        casez_tmp_349 = ldq_9_bits_uop_is_sys_pc2epc;
      5'b01010:
        casez_tmp_349 = ldq_10_bits_uop_is_sys_pc2epc;
      5'b01011:
        casez_tmp_349 = ldq_11_bits_uop_is_sys_pc2epc;
      5'b01100:
        casez_tmp_349 = ldq_12_bits_uop_is_sys_pc2epc;
      5'b01101:
        casez_tmp_349 = ldq_13_bits_uop_is_sys_pc2epc;
      5'b01110:
        casez_tmp_349 = ldq_14_bits_uop_is_sys_pc2epc;
      5'b01111:
        casez_tmp_349 = ldq_15_bits_uop_is_sys_pc2epc;
      5'b10000:
        casez_tmp_349 = ldq_16_bits_uop_is_sys_pc2epc;
      5'b10001:
        casez_tmp_349 = ldq_17_bits_uop_is_sys_pc2epc;
      5'b10010:
        casez_tmp_349 = ldq_18_bits_uop_is_sys_pc2epc;
      5'b10011:
        casez_tmp_349 = ldq_19_bits_uop_is_sys_pc2epc;
      5'b10100:
        casez_tmp_349 = ldq_20_bits_uop_is_sys_pc2epc;
      5'b10101:
        casez_tmp_349 = ldq_21_bits_uop_is_sys_pc2epc;
      5'b10110:
        casez_tmp_349 = ldq_22_bits_uop_is_sys_pc2epc;
      5'b10111:
        casez_tmp_349 = ldq_23_bits_uop_is_sys_pc2epc;
      5'b11000:
        casez_tmp_349 = ldq_24_bits_uop_is_sys_pc2epc;
      5'b11001:
        casez_tmp_349 = ldq_25_bits_uop_is_sys_pc2epc;
      5'b11010:
        casez_tmp_349 = ldq_26_bits_uop_is_sys_pc2epc;
      5'b11011:
        casez_tmp_349 = ldq_27_bits_uop_is_sys_pc2epc;
      5'b11100:
        casez_tmp_349 = ldq_28_bits_uop_is_sys_pc2epc;
      5'b11101:
        casez_tmp_349 = ldq_29_bits_uop_is_sys_pc2epc;
      5'b11110:
        casez_tmp_349 = ldq_30_bits_uop_is_sys_pc2epc;
      default:
        casez_tmp_349 = ldq_31_bits_uop_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_350;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_350 = ldq_0_bits_uop_is_unique;
      5'b00001:
        casez_tmp_350 = ldq_1_bits_uop_is_unique;
      5'b00010:
        casez_tmp_350 = ldq_2_bits_uop_is_unique;
      5'b00011:
        casez_tmp_350 = ldq_3_bits_uop_is_unique;
      5'b00100:
        casez_tmp_350 = ldq_4_bits_uop_is_unique;
      5'b00101:
        casez_tmp_350 = ldq_5_bits_uop_is_unique;
      5'b00110:
        casez_tmp_350 = ldq_6_bits_uop_is_unique;
      5'b00111:
        casez_tmp_350 = ldq_7_bits_uop_is_unique;
      5'b01000:
        casez_tmp_350 = ldq_8_bits_uop_is_unique;
      5'b01001:
        casez_tmp_350 = ldq_9_bits_uop_is_unique;
      5'b01010:
        casez_tmp_350 = ldq_10_bits_uop_is_unique;
      5'b01011:
        casez_tmp_350 = ldq_11_bits_uop_is_unique;
      5'b01100:
        casez_tmp_350 = ldq_12_bits_uop_is_unique;
      5'b01101:
        casez_tmp_350 = ldq_13_bits_uop_is_unique;
      5'b01110:
        casez_tmp_350 = ldq_14_bits_uop_is_unique;
      5'b01111:
        casez_tmp_350 = ldq_15_bits_uop_is_unique;
      5'b10000:
        casez_tmp_350 = ldq_16_bits_uop_is_unique;
      5'b10001:
        casez_tmp_350 = ldq_17_bits_uop_is_unique;
      5'b10010:
        casez_tmp_350 = ldq_18_bits_uop_is_unique;
      5'b10011:
        casez_tmp_350 = ldq_19_bits_uop_is_unique;
      5'b10100:
        casez_tmp_350 = ldq_20_bits_uop_is_unique;
      5'b10101:
        casez_tmp_350 = ldq_21_bits_uop_is_unique;
      5'b10110:
        casez_tmp_350 = ldq_22_bits_uop_is_unique;
      5'b10111:
        casez_tmp_350 = ldq_23_bits_uop_is_unique;
      5'b11000:
        casez_tmp_350 = ldq_24_bits_uop_is_unique;
      5'b11001:
        casez_tmp_350 = ldq_25_bits_uop_is_unique;
      5'b11010:
        casez_tmp_350 = ldq_26_bits_uop_is_unique;
      5'b11011:
        casez_tmp_350 = ldq_27_bits_uop_is_unique;
      5'b11100:
        casez_tmp_350 = ldq_28_bits_uop_is_unique;
      5'b11101:
        casez_tmp_350 = ldq_29_bits_uop_is_unique;
      5'b11110:
        casez_tmp_350 = ldq_30_bits_uop_is_unique;
      default:
        casez_tmp_350 = ldq_31_bits_uop_is_unique;
    endcase
  end // always @(*)
  reg         casez_tmp_351;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_351 = ldq_0_bits_uop_flush_on_commit;
      5'b00001:
        casez_tmp_351 = ldq_1_bits_uop_flush_on_commit;
      5'b00010:
        casez_tmp_351 = ldq_2_bits_uop_flush_on_commit;
      5'b00011:
        casez_tmp_351 = ldq_3_bits_uop_flush_on_commit;
      5'b00100:
        casez_tmp_351 = ldq_4_bits_uop_flush_on_commit;
      5'b00101:
        casez_tmp_351 = ldq_5_bits_uop_flush_on_commit;
      5'b00110:
        casez_tmp_351 = ldq_6_bits_uop_flush_on_commit;
      5'b00111:
        casez_tmp_351 = ldq_7_bits_uop_flush_on_commit;
      5'b01000:
        casez_tmp_351 = ldq_8_bits_uop_flush_on_commit;
      5'b01001:
        casez_tmp_351 = ldq_9_bits_uop_flush_on_commit;
      5'b01010:
        casez_tmp_351 = ldq_10_bits_uop_flush_on_commit;
      5'b01011:
        casez_tmp_351 = ldq_11_bits_uop_flush_on_commit;
      5'b01100:
        casez_tmp_351 = ldq_12_bits_uop_flush_on_commit;
      5'b01101:
        casez_tmp_351 = ldq_13_bits_uop_flush_on_commit;
      5'b01110:
        casez_tmp_351 = ldq_14_bits_uop_flush_on_commit;
      5'b01111:
        casez_tmp_351 = ldq_15_bits_uop_flush_on_commit;
      5'b10000:
        casez_tmp_351 = ldq_16_bits_uop_flush_on_commit;
      5'b10001:
        casez_tmp_351 = ldq_17_bits_uop_flush_on_commit;
      5'b10010:
        casez_tmp_351 = ldq_18_bits_uop_flush_on_commit;
      5'b10011:
        casez_tmp_351 = ldq_19_bits_uop_flush_on_commit;
      5'b10100:
        casez_tmp_351 = ldq_20_bits_uop_flush_on_commit;
      5'b10101:
        casez_tmp_351 = ldq_21_bits_uop_flush_on_commit;
      5'b10110:
        casez_tmp_351 = ldq_22_bits_uop_flush_on_commit;
      5'b10111:
        casez_tmp_351 = ldq_23_bits_uop_flush_on_commit;
      5'b11000:
        casez_tmp_351 = ldq_24_bits_uop_flush_on_commit;
      5'b11001:
        casez_tmp_351 = ldq_25_bits_uop_flush_on_commit;
      5'b11010:
        casez_tmp_351 = ldq_26_bits_uop_flush_on_commit;
      5'b11011:
        casez_tmp_351 = ldq_27_bits_uop_flush_on_commit;
      5'b11100:
        casez_tmp_351 = ldq_28_bits_uop_flush_on_commit;
      5'b11101:
        casez_tmp_351 = ldq_29_bits_uop_flush_on_commit;
      5'b11110:
        casez_tmp_351 = ldq_30_bits_uop_flush_on_commit;
      default:
        casez_tmp_351 = ldq_31_bits_uop_flush_on_commit;
    endcase
  end // always @(*)
  reg         casez_tmp_352;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_352 = ldq_0_bits_uop_ldst_is_rs1;
      5'b00001:
        casez_tmp_352 = ldq_1_bits_uop_ldst_is_rs1;
      5'b00010:
        casez_tmp_352 = ldq_2_bits_uop_ldst_is_rs1;
      5'b00011:
        casez_tmp_352 = ldq_3_bits_uop_ldst_is_rs1;
      5'b00100:
        casez_tmp_352 = ldq_4_bits_uop_ldst_is_rs1;
      5'b00101:
        casez_tmp_352 = ldq_5_bits_uop_ldst_is_rs1;
      5'b00110:
        casez_tmp_352 = ldq_6_bits_uop_ldst_is_rs1;
      5'b00111:
        casez_tmp_352 = ldq_7_bits_uop_ldst_is_rs1;
      5'b01000:
        casez_tmp_352 = ldq_8_bits_uop_ldst_is_rs1;
      5'b01001:
        casez_tmp_352 = ldq_9_bits_uop_ldst_is_rs1;
      5'b01010:
        casez_tmp_352 = ldq_10_bits_uop_ldst_is_rs1;
      5'b01011:
        casez_tmp_352 = ldq_11_bits_uop_ldst_is_rs1;
      5'b01100:
        casez_tmp_352 = ldq_12_bits_uop_ldst_is_rs1;
      5'b01101:
        casez_tmp_352 = ldq_13_bits_uop_ldst_is_rs1;
      5'b01110:
        casez_tmp_352 = ldq_14_bits_uop_ldst_is_rs1;
      5'b01111:
        casez_tmp_352 = ldq_15_bits_uop_ldst_is_rs1;
      5'b10000:
        casez_tmp_352 = ldq_16_bits_uop_ldst_is_rs1;
      5'b10001:
        casez_tmp_352 = ldq_17_bits_uop_ldst_is_rs1;
      5'b10010:
        casez_tmp_352 = ldq_18_bits_uop_ldst_is_rs1;
      5'b10011:
        casez_tmp_352 = ldq_19_bits_uop_ldst_is_rs1;
      5'b10100:
        casez_tmp_352 = ldq_20_bits_uop_ldst_is_rs1;
      5'b10101:
        casez_tmp_352 = ldq_21_bits_uop_ldst_is_rs1;
      5'b10110:
        casez_tmp_352 = ldq_22_bits_uop_ldst_is_rs1;
      5'b10111:
        casez_tmp_352 = ldq_23_bits_uop_ldst_is_rs1;
      5'b11000:
        casez_tmp_352 = ldq_24_bits_uop_ldst_is_rs1;
      5'b11001:
        casez_tmp_352 = ldq_25_bits_uop_ldst_is_rs1;
      5'b11010:
        casez_tmp_352 = ldq_26_bits_uop_ldst_is_rs1;
      5'b11011:
        casez_tmp_352 = ldq_27_bits_uop_ldst_is_rs1;
      5'b11100:
        casez_tmp_352 = ldq_28_bits_uop_ldst_is_rs1;
      5'b11101:
        casez_tmp_352 = ldq_29_bits_uop_ldst_is_rs1;
      5'b11110:
        casez_tmp_352 = ldq_30_bits_uop_ldst_is_rs1;
      default:
        casez_tmp_352 = ldq_31_bits_uop_ldst_is_rs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_353;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_353 = ldq_0_bits_uop_ldst;
      5'b00001:
        casez_tmp_353 = ldq_1_bits_uop_ldst;
      5'b00010:
        casez_tmp_353 = ldq_2_bits_uop_ldst;
      5'b00011:
        casez_tmp_353 = ldq_3_bits_uop_ldst;
      5'b00100:
        casez_tmp_353 = ldq_4_bits_uop_ldst;
      5'b00101:
        casez_tmp_353 = ldq_5_bits_uop_ldst;
      5'b00110:
        casez_tmp_353 = ldq_6_bits_uop_ldst;
      5'b00111:
        casez_tmp_353 = ldq_7_bits_uop_ldst;
      5'b01000:
        casez_tmp_353 = ldq_8_bits_uop_ldst;
      5'b01001:
        casez_tmp_353 = ldq_9_bits_uop_ldst;
      5'b01010:
        casez_tmp_353 = ldq_10_bits_uop_ldst;
      5'b01011:
        casez_tmp_353 = ldq_11_bits_uop_ldst;
      5'b01100:
        casez_tmp_353 = ldq_12_bits_uop_ldst;
      5'b01101:
        casez_tmp_353 = ldq_13_bits_uop_ldst;
      5'b01110:
        casez_tmp_353 = ldq_14_bits_uop_ldst;
      5'b01111:
        casez_tmp_353 = ldq_15_bits_uop_ldst;
      5'b10000:
        casez_tmp_353 = ldq_16_bits_uop_ldst;
      5'b10001:
        casez_tmp_353 = ldq_17_bits_uop_ldst;
      5'b10010:
        casez_tmp_353 = ldq_18_bits_uop_ldst;
      5'b10011:
        casez_tmp_353 = ldq_19_bits_uop_ldst;
      5'b10100:
        casez_tmp_353 = ldq_20_bits_uop_ldst;
      5'b10101:
        casez_tmp_353 = ldq_21_bits_uop_ldst;
      5'b10110:
        casez_tmp_353 = ldq_22_bits_uop_ldst;
      5'b10111:
        casez_tmp_353 = ldq_23_bits_uop_ldst;
      5'b11000:
        casez_tmp_353 = ldq_24_bits_uop_ldst;
      5'b11001:
        casez_tmp_353 = ldq_25_bits_uop_ldst;
      5'b11010:
        casez_tmp_353 = ldq_26_bits_uop_ldst;
      5'b11011:
        casez_tmp_353 = ldq_27_bits_uop_ldst;
      5'b11100:
        casez_tmp_353 = ldq_28_bits_uop_ldst;
      5'b11101:
        casez_tmp_353 = ldq_29_bits_uop_ldst;
      5'b11110:
        casez_tmp_353 = ldq_30_bits_uop_ldst;
      default:
        casez_tmp_353 = ldq_31_bits_uop_ldst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_354;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_354 = ldq_0_bits_uop_lrs1;
      5'b00001:
        casez_tmp_354 = ldq_1_bits_uop_lrs1;
      5'b00010:
        casez_tmp_354 = ldq_2_bits_uop_lrs1;
      5'b00011:
        casez_tmp_354 = ldq_3_bits_uop_lrs1;
      5'b00100:
        casez_tmp_354 = ldq_4_bits_uop_lrs1;
      5'b00101:
        casez_tmp_354 = ldq_5_bits_uop_lrs1;
      5'b00110:
        casez_tmp_354 = ldq_6_bits_uop_lrs1;
      5'b00111:
        casez_tmp_354 = ldq_7_bits_uop_lrs1;
      5'b01000:
        casez_tmp_354 = ldq_8_bits_uop_lrs1;
      5'b01001:
        casez_tmp_354 = ldq_9_bits_uop_lrs1;
      5'b01010:
        casez_tmp_354 = ldq_10_bits_uop_lrs1;
      5'b01011:
        casez_tmp_354 = ldq_11_bits_uop_lrs1;
      5'b01100:
        casez_tmp_354 = ldq_12_bits_uop_lrs1;
      5'b01101:
        casez_tmp_354 = ldq_13_bits_uop_lrs1;
      5'b01110:
        casez_tmp_354 = ldq_14_bits_uop_lrs1;
      5'b01111:
        casez_tmp_354 = ldq_15_bits_uop_lrs1;
      5'b10000:
        casez_tmp_354 = ldq_16_bits_uop_lrs1;
      5'b10001:
        casez_tmp_354 = ldq_17_bits_uop_lrs1;
      5'b10010:
        casez_tmp_354 = ldq_18_bits_uop_lrs1;
      5'b10011:
        casez_tmp_354 = ldq_19_bits_uop_lrs1;
      5'b10100:
        casez_tmp_354 = ldq_20_bits_uop_lrs1;
      5'b10101:
        casez_tmp_354 = ldq_21_bits_uop_lrs1;
      5'b10110:
        casez_tmp_354 = ldq_22_bits_uop_lrs1;
      5'b10111:
        casez_tmp_354 = ldq_23_bits_uop_lrs1;
      5'b11000:
        casez_tmp_354 = ldq_24_bits_uop_lrs1;
      5'b11001:
        casez_tmp_354 = ldq_25_bits_uop_lrs1;
      5'b11010:
        casez_tmp_354 = ldq_26_bits_uop_lrs1;
      5'b11011:
        casez_tmp_354 = ldq_27_bits_uop_lrs1;
      5'b11100:
        casez_tmp_354 = ldq_28_bits_uop_lrs1;
      5'b11101:
        casez_tmp_354 = ldq_29_bits_uop_lrs1;
      5'b11110:
        casez_tmp_354 = ldq_30_bits_uop_lrs1;
      default:
        casez_tmp_354 = ldq_31_bits_uop_lrs1;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_355;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_355 = ldq_0_bits_uop_lrs2;
      5'b00001:
        casez_tmp_355 = ldq_1_bits_uop_lrs2;
      5'b00010:
        casez_tmp_355 = ldq_2_bits_uop_lrs2;
      5'b00011:
        casez_tmp_355 = ldq_3_bits_uop_lrs2;
      5'b00100:
        casez_tmp_355 = ldq_4_bits_uop_lrs2;
      5'b00101:
        casez_tmp_355 = ldq_5_bits_uop_lrs2;
      5'b00110:
        casez_tmp_355 = ldq_6_bits_uop_lrs2;
      5'b00111:
        casez_tmp_355 = ldq_7_bits_uop_lrs2;
      5'b01000:
        casez_tmp_355 = ldq_8_bits_uop_lrs2;
      5'b01001:
        casez_tmp_355 = ldq_9_bits_uop_lrs2;
      5'b01010:
        casez_tmp_355 = ldq_10_bits_uop_lrs2;
      5'b01011:
        casez_tmp_355 = ldq_11_bits_uop_lrs2;
      5'b01100:
        casez_tmp_355 = ldq_12_bits_uop_lrs2;
      5'b01101:
        casez_tmp_355 = ldq_13_bits_uop_lrs2;
      5'b01110:
        casez_tmp_355 = ldq_14_bits_uop_lrs2;
      5'b01111:
        casez_tmp_355 = ldq_15_bits_uop_lrs2;
      5'b10000:
        casez_tmp_355 = ldq_16_bits_uop_lrs2;
      5'b10001:
        casez_tmp_355 = ldq_17_bits_uop_lrs2;
      5'b10010:
        casez_tmp_355 = ldq_18_bits_uop_lrs2;
      5'b10011:
        casez_tmp_355 = ldq_19_bits_uop_lrs2;
      5'b10100:
        casez_tmp_355 = ldq_20_bits_uop_lrs2;
      5'b10101:
        casez_tmp_355 = ldq_21_bits_uop_lrs2;
      5'b10110:
        casez_tmp_355 = ldq_22_bits_uop_lrs2;
      5'b10111:
        casez_tmp_355 = ldq_23_bits_uop_lrs2;
      5'b11000:
        casez_tmp_355 = ldq_24_bits_uop_lrs2;
      5'b11001:
        casez_tmp_355 = ldq_25_bits_uop_lrs2;
      5'b11010:
        casez_tmp_355 = ldq_26_bits_uop_lrs2;
      5'b11011:
        casez_tmp_355 = ldq_27_bits_uop_lrs2;
      5'b11100:
        casez_tmp_355 = ldq_28_bits_uop_lrs2;
      5'b11101:
        casez_tmp_355 = ldq_29_bits_uop_lrs2;
      5'b11110:
        casez_tmp_355 = ldq_30_bits_uop_lrs2;
      default:
        casez_tmp_355 = ldq_31_bits_uop_lrs2;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_356;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_356 = ldq_0_bits_uop_lrs3;
      5'b00001:
        casez_tmp_356 = ldq_1_bits_uop_lrs3;
      5'b00010:
        casez_tmp_356 = ldq_2_bits_uop_lrs3;
      5'b00011:
        casez_tmp_356 = ldq_3_bits_uop_lrs3;
      5'b00100:
        casez_tmp_356 = ldq_4_bits_uop_lrs3;
      5'b00101:
        casez_tmp_356 = ldq_5_bits_uop_lrs3;
      5'b00110:
        casez_tmp_356 = ldq_6_bits_uop_lrs3;
      5'b00111:
        casez_tmp_356 = ldq_7_bits_uop_lrs3;
      5'b01000:
        casez_tmp_356 = ldq_8_bits_uop_lrs3;
      5'b01001:
        casez_tmp_356 = ldq_9_bits_uop_lrs3;
      5'b01010:
        casez_tmp_356 = ldq_10_bits_uop_lrs3;
      5'b01011:
        casez_tmp_356 = ldq_11_bits_uop_lrs3;
      5'b01100:
        casez_tmp_356 = ldq_12_bits_uop_lrs3;
      5'b01101:
        casez_tmp_356 = ldq_13_bits_uop_lrs3;
      5'b01110:
        casez_tmp_356 = ldq_14_bits_uop_lrs3;
      5'b01111:
        casez_tmp_356 = ldq_15_bits_uop_lrs3;
      5'b10000:
        casez_tmp_356 = ldq_16_bits_uop_lrs3;
      5'b10001:
        casez_tmp_356 = ldq_17_bits_uop_lrs3;
      5'b10010:
        casez_tmp_356 = ldq_18_bits_uop_lrs3;
      5'b10011:
        casez_tmp_356 = ldq_19_bits_uop_lrs3;
      5'b10100:
        casez_tmp_356 = ldq_20_bits_uop_lrs3;
      5'b10101:
        casez_tmp_356 = ldq_21_bits_uop_lrs3;
      5'b10110:
        casez_tmp_356 = ldq_22_bits_uop_lrs3;
      5'b10111:
        casez_tmp_356 = ldq_23_bits_uop_lrs3;
      5'b11000:
        casez_tmp_356 = ldq_24_bits_uop_lrs3;
      5'b11001:
        casez_tmp_356 = ldq_25_bits_uop_lrs3;
      5'b11010:
        casez_tmp_356 = ldq_26_bits_uop_lrs3;
      5'b11011:
        casez_tmp_356 = ldq_27_bits_uop_lrs3;
      5'b11100:
        casez_tmp_356 = ldq_28_bits_uop_lrs3;
      5'b11101:
        casez_tmp_356 = ldq_29_bits_uop_lrs3;
      5'b11110:
        casez_tmp_356 = ldq_30_bits_uop_lrs3;
      default:
        casez_tmp_356 = ldq_31_bits_uop_lrs3;
    endcase
  end // always @(*)
  reg         casez_tmp_357;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_357 = ldq_0_bits_uop_ldst_val;
      5'b00001:
        casez_tmp_357 = ldq_1_bits_uop_ldst_val;
      5'b00010:
        casez_tmp_357 = ldq_2_bits_uop_ldst_val;
      5'b00011:
        casez_tmp_357 = ldq_3_bits_uop_ldst_val;
      5'b00100:
        casez_tmp_357 = ldq_4_bits_uop_ldst_val;
      5'b00101:
        casez_tmp_357 = ldq_5_bits_uop_ldst_val;
      5'b00110:
        casez_tmp_357 = ldq_6_bits_uop_ldst_val;
      5'b00111:
        casez_tmp_357 = ldq_7_bits_uop_ldst_val;
      5'b01000:
        casez_tmp_357 = ldq_8_bits_uop_ldst_val;
      5'b01001:
        casez_tmp_357 = ldq_9_bits_uop_ldst_val;
      5'b01010:
        casez_tmp_357 = ldq_10_bits_uop_ldst_val;
      5'b01011:
        casez_tmp_357 = ldq_11_bits_uop_ldst_val;
      5'b01100:
        casez_tmp_357 = ldq_12_bits_uop_ldst_val;
      5'b01101:
        casez_tmp_357 = ldq_13_bits_uop_ldst_val;
      5'b01110:
        casez_tmp_357 = ldq_14_bits_uop_ldst_val;
      5'b01111:
        casez_tmp_357 = ldq_15_bits_uop_ldst_val;
      5'b10000:
        casez_tmp_357 = ldq_16_bits_uop_ldst_val;
      5'b10001:
        casez_tmp_357 = ldq_17_bits_uop_ldst_val;
      5'b10010:
        casez_tmp_357 = ldq_18_bits_uop_ldst_val;
      5'b10011:
        casez_tmp_357 = ldq_19_bits_uop_ldst_val;
      5'b10100:
        casez_tmp_357 = ldq_20_bits_uop_ldst_val;
      5'b10101:
        casez_tmp_357 = ldq_21_bits_uop_ldst_val;
      5'b10110:
        casez_tmp_357 = ldq_22_bits_uop_ldst_val;
      5'b10111:
        casez_tmp_357 = ldq_23_bits_uop_ldst_val;
      5'b11000:
        casez_tmp_357 = ldq_24_bits_uop_ldst_val;
      5'b11001:
        casez_tmp_357 = ldq_25_bits_uop_ldst_val;
      5'b11010:
        casez_tmp_357 = ldq_26_bits_uop_ldst_val;
      5'b11011:
        casez_tmp_357 = ldq_27_bits_uop_ldst_val;
      5'b11100:
        casez_tmp_357 = ldq_28_bits_uop_ldst_val;
      5'b11101:
        casez_tmp_357 = ldq_29_bits_uop_ldst_val;
      5'b11110:
        casez_tmp_357 = ldq_30_bits_uop_ldst_val;
      default:
        casez_tmp_357 = ldq_31_bits_uop_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_358;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_358 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_358 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_358 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_358 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_358 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_358 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_358 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_358 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_358 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_358 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_358 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_358 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_358 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_358 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_358 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_358 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_358 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_358 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_358 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_358 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_358 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_358 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_358 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_358 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_358 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_358 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_358 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_358 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_358 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_358 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_358 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_358 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_359;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_359 = ldq_0_bits_uop_lrs1_rtype;
      5'b00001:
        casez_tmp_359 = ldq_1_bits_uop_lrs1_rtype;
      5'b00010:
        casez_tmp_359 = ldq_2_bits_uop_lrs1_rtype;
      5'b00011:
        casez_tmp_359 = ldq_3_bits_uop_lrs1_rtype;
      5'b00100:
        casez_tmp_359 = ldq_4_bits_uop_lrs1_rtype;
      5'b00101:
        casez_tmp_359 = ldq_5_bits_uop_lrs1_rtype;
      5'b00110:
        casez_tmp_359 = ldq_6_bits_uop_lrs1_rtype;
      5'b00111:
        casez_tmp_359 = ldq_7_bits_uop_lrs1_rtype;
      5'b01000:
        casez_tmp_359 = ldq_8_bits_uop_lrs1_rtype;
      5'b01001:
        casez_tmp_359 = ldq_9_bits_uop_lrs1_rtype;
      5'b01010:
        casez_tmp_359 = ldq_10_bits_uop_lrs1_rtype;
      5'b01011:
        casez_tmp_359 = ldq_11_bits_uop_lrs1_rtype;
      5'b01100:
        casez_tmp_359 = ldq_12_bits_uop_lrs1_rtype;
      5'b01101:
        casez_tmp_359 = ldq_13_bits_uop_lrs1_rtype;
      5'b01110:
        casez_tmp_359 = ldq_14_bits_uop_lrs1_rtype;
      5'b01111:
        casez_tmp_359 = ldq_15_bits_uop_lrs1_rtype;
      5'b10000:
        casez_tmp_359 = ldq_16_bits_uop_lrs1_rtype;
      5'b10001:
        casez_tmp_359 = ldq_17_bits_uop_lrs1_rtype;
      5'b10010:
        casez_tmp_359 = ldq_18_bits_uop_lrs1_rtype;
      5'b10011:
        casez_tmp_359 = ldq_19_bits_uop_lrs1_rtype;
      5'b10100:
        casez_tmp_359 = ldq_20_bits_uop_lrs1_rtype;
      5'b10101:
        casez_tmp_359 = ldq_21_bits_uop_lrs1_rtype;
      5'b10110:
        casez_tmp_359 = ldq_22_bits_uop_lrs1_rtype;
      5'b10111:
        casez_tmp_359 = ldq_23_bits_uop_lrs1_rtype;
      5'b11000:
        casez_tmp_359 = ldq_24_bits_uop_lrs1_rtype;
      5'b11001:
        casez_tmp_359 = ldq_25_bits_uop_lrs1_rtype;
      5'b11010:
        casez_tmp_359 = ldq_26_bits_uop_lrs1_rtype;
      5'b11011:
        casez_tmp_359 = ldq_27_bits_uop_lrs1_rtype;
      5'b11100:
        casez_tmp_359 = ldq_28_bits_uop_lrs1_rtype;
      5'b11101:
        casez_tmp_359 = ldq_29_bits_uop_lrs1_rtype;
      5'b11110:
        casez_tmp_359 = ldq_30_bits_uop_lrs1_rtype;
      default:
        casez_tmp_359 = ldq_31_bits_uop_lrs1_rtype;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_360;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_360 = ldq_0_bits_uop_lrs2_rtype;
      5'b00001:
        casez_tmp_360 = ldq_1_bits_uop_lrs2_rtype;
      5'b00010:
        casez_tmp_360 = ldq_2_bits_uop_lrs2_rtype;
      5'b00011:
        casez_tmp_360 = ldq_3_bits_uop_lrs2_rtype;
      5'b00100:
        casez_tmp_360 = ldq_4_bits_uop_lrs2_rtype;
      5'b00101:
        casez_tmp_360 = ldq_5_bits_uop_lrs2_rtype;
      5'b00110:
        casez_tmp_360 = ldq_6_bits_uop_lrs2_rtype;
      5'b00111:
        casez_tmp_360 = ldq_7_bits_uop_lrs2_rtype;
      5'b01000:
        casez_tmp_360 = ldq_8_bits_uop_lrs2_rtype;
      5'b01001:
        casez_tmp_360 = ldq_9_bits_uop_lrs2_rtype;
      5'b01010:
        casez_tmp_360 = ldq_10_bits_uop_lrs2_rtype;
      5'b01011:
        casez_tmp_360 = ldq_11_bits_uop_lrs2_rtype;
      5'b01100:
        casez_tmp_360 = ldq_12_bits_uop_lrs2_rtype;
      5'b01101:
        casez_tmp_360 = ldq_13_bits_uop_lrs2_rtype;
      5'b01110:
        casez_tmp_360 = ldq_14_bits_uop_lrs2_rtype;
      5'b01111:
        casez_tmp_360 = ldq_15_bits_uop_lrs2_rtype;
      5'b10000:
        casez_tmp_360 = ldq_16_bits_uop_lrs2_rtype;
      5'b10001:
        casez_tmp_360 = ldq_17_bits_uop_lrs2_rtype;
      5'b10010:
        casez_tmp_360 = ldq_18_bits_uop_lrs2_rtype;
      5'b10011:
        casez_tmp_360 = ldq_19_bits_uop_lrs2_rtype;
      5'b10100:
        casez_tmp_360 = ldq_20_bits_uop_lrs2_rtype;
      5'b10101:
        casez_tmp_360 = ldq_21_bits_uop_lrs2_rtype;
      5'b10110:
        casez_tmp_360 = ldq_22_bits_uop_lrs2_rtype;
      5'b10111:
        casez_tmp_360 = ldq_23_bits_uop_lrs2_rtype;
      5'b11000:
        casez_tmp_360 = ldq_24_bits_uop_lrs2_rtype;
      5'b11001:
        casez_tmp_360 = ldq_25_bits_uop_lrs2_rtype;
      5'b11010:
        casez_tmp_360 = ldq_26_bits_uop_lrs2_rtype;
      5'b11011:
        casez_tmp_360 = ldq_27_bits_uop_lrs2_rtype;
      5'b11100:
        casez_tmp_360 = ldq_28_bits_uop_lrs2_rtype;
      5'b11101:
        casez_tmp_360 = ldq_29_bits_uop_lrs2_rtype;
      5'b11110:
        casez_tmp_360 = ldq_30_bits_uop_lrs2_rtype;
      default:
        casez_tmp_360 = ldq_31_bits_uop_lrs2_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_361;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_361 = ldq_0_bits_uop_frs3_en;
      5'b00001:
        casez_tmp_361 = ldq_1_bits_uop_frs3_en;
      5'b00010:
        casez_tmp_361 = ldq_2_bits_uop_frs3_en;
      5'b00011:
        casez_tmp_361 = ldq_3_bits_uop_frs3_en;
      5'b00100:
        casez_tmp_361 = ldq_4_bits_uop_frs3_en;
      5'b00101:
        casez_tmp_361 = ldq_5_bits_uop_frs3_en;
      5'b00110:
        casez_tmp_361 = ldq_6_bits_uop_frs3_en;
      5'b00111:
        casez_tmp_361 = ldq_7_bits_uop_frs3_en;
      5'b01000:
        casez_tmp_361 = ldq_8_bits_uop_frs3_en;
      5'b01001:
        casez_tmp_361 = ldq_9_bits_uop_frs3_en;
      5'b01010:
        casez_tmp_361 = ldq_10_bits_uop_frs3_en;
      5'b01011:
        casez_tmp_361 = ldq_11_bits_uop_frs3_en;
      5'b01100:
        casez_tmp_361 = ldq_12_bits_uop_frs3_en;
      5'b01101:
        casez_tmp_361 = ldq_13_bits_uop_frs3_en;
      5'b01110:
        casez_tmp_361 = ldq_14_bits_uop_frs3_en;
      5'b01111:
        casez_tmp_361 = ldq_15_bits_uop_frs3_en;
      5'b10000:
        casez_tmp_361 = ldq_16_bits_uop_frs3_en;
      5'b10001:
        casez_tmp_361 = ldq_17_bits_uop_frs3_en;
      5'b10010:
        casez_tmp_361 = ldq_18_bits_uop_frs3_en;
      5'b10011:
        casez_tmp_361 = ldq_19_bits_uop_frs3_en;
      5'b10100:
        casez_tmp_361 = ldq_20_bits_uop_frs3_en;
      5'b10101:
        casez_tmp_361 = ldq_21_bits_uop_frs3_en;
      5'b10110:
        casez_tmp_361 = ldq_22_bits_uop_frs3_en;
      5'b10111:
        casez_tmp_361 = ldq_23_bits_uop_frs3_en;
      5'b11000:
        casez_tmp_361 = ldq_24_bits_uop_frs3_en;
      5'b11001:
        casez_tmp_361 = ldq_25_bits_uop_frs3_en;
      5'b11010:
        casez_tmp_361 = ldq_26_bits_uop_frs3_en;
      5'b11011:
        casez_tmp_361 = ldq_27_bits_uop_frs3_en;
      5'b11100:
        casez_tmp_361 = ldq_28_bits_uop_frs3_en;
      5'b11101:
        casez_tmp_361 = ldq_29_bits_uop_frs3_en;
      5'b11110:
        casez_tmp_361 = ldq_30_bits_uop_frs3_en;
      default:
        casez_tmp_361 = ldq_31_bits_uop_frs3_en;
    endcase
  end // always @(*)
  reg         casez_tmp_362;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_362 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_362 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_362 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_362 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_362 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_362 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_362 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_362 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_362 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_362 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_362 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_362 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_362 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_362 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_362 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_362 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_362 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_362 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_362 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_362 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_362 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_362 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_362 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_362 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_362 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_362 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_362 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_362 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_362 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_362 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_362 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_362 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  reg         casez_tmp_363;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_363 = ldq_0_bits_uop_fp_single;
      5'b00001:
        casez_tmp_363 = ldq_1_bits_uop_fp_single;
      5'b00010:
        casez_tmp_363 = ldq_2_bits_uop_fp_single;
      5'b00011:
        casez_tmp_363 = ldq_3_bits_uop_fp_single;
      5'b00100:
        casez_tmp_363 = ldq_4_bits_uop_fp_single;
      5'b00101:
        casez_tmp_363 = ldq_5_bits_uop_fp_single;
      5'b00110:
        casez_tmp_363 = ldq_6_bits_uop_fp_single;
      5'b00111:
        casez_tmp_363 = ldq_7_bits_uop_fp_single;
      5'b01000:
        casez_tmp_363 = ldq_8_bits_uop_fp_single;
      5'b01001:
        casez_tmp_363 = ldq_9_bits_uop_fp_single;
      5'b01010:
        casez_tmp_363 = ldq_10_bits_uop_fp_single;
      5'b01011:
        casez_tmp_363 = ldq_11_bits_uop_fp_single;
      5'b01100:
        casez_tmp_363 = ldq_12_bits_uop_fp_single;
      5'b01101:
        casez_tmp_363 = ldq_13_bits_uop_fp_single;
      5'b01110:
        casez_tmp_363 = ldq_14_bits_uop_fp_single;
      5'b01111:
        casez_tmp_363 = ldq_15_bits_uop_fp_single;
      5'b10000:
        casez_tmp_363 = ldq_16_bits_uop_fp_single;
      5'b10001:
        casez_tmp_363 = ldq_17_bits_uop_fp_single;
      5'b10010:
        casez_tmp_363 = ldq_18_bits_uop_fp_single;
      5'b10011:
        casez_tmp_363 = ldq_19_bits_uop_fp_single;
      5'b10100:
        casez_tmp_363 = ldq_20_bits_uop_fp_single;
      5'b10101:
        casez_tmp_363 = ldq_21_bits_uop_fp_single;
      5'b10110:
        casez_tmp_363 = ldq_22_bits_uop_fp_single;
      5'b10111:
        casez_tmp_363 = ldq_23_bits_uop_fp_single;
      5'b11000:
        casez_tmp_363 = ldq_24_bits_uop_fp_single;
      5'b11001:
        casez_tmp_363 = ldq_25_bits_uop_fp_single;
      5'b11010:
        casez_tmp_363 = ldq_26_bits_uop_fp_single;
      5'b11011:
        casez_tmp_363 = ldq_27_bits_uop_fp_single;
      5'b11100:
        casez_tmp_363 = ldq_28_bits_uop_fp_single;
      5'b11101:
        casez_tmp_363 = ldq_29_bits_uop_fp_single;
      5'b11110:
        casez_tmp_363 = ldq_30_bits_uop_fp_single;
      default:
        casez_tmp_363 = ldq_31_bits_uop_fp_single;
    endcase
  end // always @(*)
  reg         casez_tmp_364;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_364 = ldq_0_bits_uop_xcpt_pf_if;
      5'b00001:
        casez_tmp_364 = ldq_1_bits_uop_xcpt_pf_if;
      5'b00010:
        casez_tmp_364 = ldq_2_bits_uop_xcpt_pf_if;
      5'b00011:
        casez_tmp_364 = ldq_3_bits_uop_xcpt_pf_if;
      5'b00100:
        casez_tmp_364 = ldq_4_bits_uop_xcpt_pf_if;
      5'b00101:
        casez_tmp_364 = ldq_5_bits_uop_xcpt_pf_if;
      5'b00110:
        casez_tmp_364 = ldq_6_bits_uop_xcpt_pf_if;
      5'b00111:
        casez_tmp_364 = ldq_7_bits_uop_xcpt_pf_if;
      5'b01000:
        casez_tmp_364 = ldq_8_bits_uop_xcpt_pf_if;
      5'b01001:
        casez_tmp_364 = ldq_9_bits_uop_xcpt_pf_if;
      5'b01010:
        casez_tmp_364 = ldq_10_bits_uop_xcpt_pf_if;
      5'b01011:
        casez_tmp_364 = ldq_11_bits_uop_xcpt_pf_if;
      5'b01100:
        casez_tmp_364 = ldq_12_bits_uop_xcpt_pf_if;
      5'b01101:
        casez_tmp_364 = ldq_13_bits_uop_xcpt_pf_if;
      5'b01110:
        casez_tmp_364 = ldq_14_bits_uop_xcpt_pf_if;
      5'b01111:
        casez_tmp_364 = ldq_15_bits_uop_xcpt_pf_if;
      5'b10000:
        casez_tmp_364 = ldq_16_bits_uop_xcpt_pf_if;
      5'b10001:
        casez_tmp_364 = ldq_17_bits_uop_xcpt_pf_if;
      5'b10010:
        casez_tmp_364 = ldq_18_bits_uop_xcpt_pf_if;
      5'b10011:
        casez_tmp_364 = ldq_19_bits_uop_xcpt_pf_if;
      5'b10100:
        casez_tmp_364 = ldq_20_bits_uop_xcpt_pf_if;
      5'b10101:
        casez_tmp_364 = ldq_21_bits_uop_xcpt_pf_if;
      5'b10110:
        casez_tmp_364 = ldq_22_bits_uop_xcpt_pf_if;
      5'b10111:
        casez_tmp_364 = ldq_23_bits_uop_xcpt_pf_if;
      5'b11000:
        casez_tmp_364 = ldq_24_bits_uop_xcpt_pf_if;
      5'b11001:
        casez_tmp_364 = ldq_25_bits_uop_xcpt_pf_if;
      5'b11010:
        casez_tmp_364 = ldq_26_bits_uop_xcpt_pf_if;
      5'b11011:
        casez_tmp_364 = ldq_27_bits_uop_xcpt_pf_if;
      5'b11100:
        casez_tmp_364 = ldq_28_bits_uop_xcpt_pf_if;
      5'b11101:
        casez_tmp_364 = ldq_29_bits_uop_xcpt_pf_if;
      5'b11110:
        casez_tmp_364 = ldq_30_bits_uop_xcpt_pf_if;
      default:
        casez_tmp_364 = ldq_31_bits_uop_xcpt_pf_if;
    endcase
  end // always @(*)
  reg         casez_tmp_365;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_365 = ldq_0_bits_uop_xcpt_ae_if;
      5'b00001:
        casez_tmp_365 = ldq_1_bits_uop_xcpt_ae_if;
      5'b00010:
        casez_tmp_365 = ldq_2_bits_uop_xcpt_ae_if;
      5'b00011:
        casez_tmp_365 = ldq_3_bits_uop_xcpt_ae_if;
      5'b00100:
        casez_tmp_365 = ldq_4_bits_uop_xcpt_ae_if;
      5'b00101:
        casez_tmp_365 = ldq_5_bits_uop_xcpt_ae_if;
      5'b00110:
        casez_tmp_365 = ldq_6_bits_uop_xcpt_ae_if;
      5'b00111:
        casez_tmp_365 = ldq_7_bits_uop_xcpt_ae_if;
      5'b01000:
        casez_tmp_365 = ldq_8_bits_uop_xcpt_ae_if;
      5'b01001:
        casez_tmp_365 = ldq_9_bits_uop_xcpt_ae_if;
      5'b01010:
        casez_tmp_365 = ldq_10_bits_uop_xcpt_ae_if;
      5'b01011:
        casez_tmp_365 = ldq_11_bits_uop_xcpt_ae_if;
      5'b01100:
        casez_tmp_365 = ldq_12_bits_uop_xcpt_ae_if;
      5'b01101:
        casez_tmp_365 = ldq_13_bits_uop_xcpt_ae_if;
      5'b01110:
        casez_tmp_365 = ldq_14_bits_uop_xcpt_ae_if;
      5'b01111:
        casez_tmp_365 = ldq_15_bits_uop_xcpt_ae_if;
      5'b10000:
        casez_tmp_365 = ldq_16_bits_uop_xcpt_ae_if;
      5'b10001:
        casez_tmp_365 = ldq_17_bits_uop_xcpt_ae_if;
      5'b10010:
        casez_tmp_365 = ldq_18_bits_uop_xcpt_ae_if;
      5'b10011:
        casez_tmp_365 = ldq_19_bits_uop_xcpt_ae_if;
      5'b10100:
        casez_tmp_365 = ldq_20_bits_uop_xcpt_ae_if;
      5'b10101:
        casez_tmp_365 = ldq_21_bits_uop_xcpt_ae_if;
      5'b10110:
        casez_tmp_365 = ldq_22_bits_uop_xcpt_ae_if;
      5'b10111:
        casez_tmp_365 = ldq_23_bits_uop_xcpt_ae_if;
      5'b11000:
        casez_tmp_365 = ldq_24_bits_uop_xcpt_ae_if;
      5'b11001:
        casez_tmp_365 = ldq_25_bits_uop_xcpt_ae_if;
      5'b11010:
        casez_tmp_365 = ldq_26_bits_uop_xcpt_ae_if;
      5'b11011:
        casez_tmp_365 = ldq_27_bits_uop_xcpt_ae_if;
      5'b11100:
        casez_tmp_365 = ldq_28_bits_uop_xcpt_ae_if;
      5'b11101:
        casez_tmp_365 = ldq_29_bits_uop_xcpt_ae_if;
      5'b11110:
        casez_tmp_365 = ldq_30_bits_uop_xcpt_ae_if;
      default:
        casez_tmp_365 = ldq_31_bits_uop_xcpt_ae_if;
    endcase
  end // always @(*)
  reg         casez_tmp_366;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_366 = ldq_0_bits_uop_xcpt_ma_if;
      5'b00001:
        casez_tmp_366 = ldq_1_bits_uop_xcpt_ma_if;
      5'b00010:
        casez_tmp_366 = ldq_2_bits_uop_xcpt_ma_if;
      5'b00011:
        casez_tmp_366 = ldq_3_bits_uop_xcpt_ma_if;
      5'b00100:
        casez_tmp_366 = ldq_4_bits_uop_xcpt_ma_if;
      5'b00101:
        casez_tmp_366 = ldq_5_bits_uop_xcpt_ma_if;
      5'b00110:
        casez_tmp_366 = ldq_6_bits_uop_xcpt_ma_if;
      5'b00111:
        casez_tmp_366 = ldq_7_bits_uop_xcpt_ma_if;
      5'b01000:
        casez_tmp_366 = ldq_8_bits_uop_xcpt_ma_if;
      5'b01001:
        casez_tmp_366 = ldq_9_bits_uop_xcpt_ma_if;
      5'b01010:
        casez_tmp_366 = ldq_10_bits_uop_xcpt_ma_if;
      5'b01011:
        casez_tmp_366 = ldq_11_bits_uop_xcpt_ma_if;
      5'b01100:
        casez_tmp_366 = ldq_12_bits_uop_xcpt_ma_if;
      5'b01101:
        casez_tmp_366 = ldq_13_bits_uop_xcpt_ma_if;
      5'b01110:
        casez_tmp_366 = ldq_14_bits_uop_xcpt_ma_if;
      5'b01111:
        casez_tmp_366 = ldq_15_bits_uop_xcpt_ma_if;
      5'b10000:
        casez_tmp_366 = ldq_16_bits_uop_xcpt_ma_if;
      5'b10001:
        casez_tmp_366 = ldq_17_bits_uop_xcpt_ma_if;
      5'b10010:
        casez_tmp_366 = ldq_18_bits_uop_xcpt_ma_if;
      5'b10011:
        casez_tmp_366 = ldq_19_bits_uop_xcpt_ma_if;
      5'b10100:
        casez_tmp_366 = ldq_20_bits_uop_xcpt_ma_if;
      5'b10101:
        casez_tmp_366 = ldq_21_bits_uop_xcpt_ma_if;
      5'b10110:
        casez_tmp_366 = ldq_22_bits_uop_xcpt_ma_if;
      5'b10111:
        casez_tmp_366 = ldq_23_bits_uop_xcpt_ma_if;
      5'b11000:
        casez_tmp_366 = ldq_24_bits_uop_xcpt_ma_if;
      5'b11001:
        casez_tmp_366 = ldq_25_bits_uop_xcpt_ma_if;
      5'b11010:
        casez_tmp_366 = ldq_26_bits_uop_xcpt_ma_if;
      5'b11011:
        casez_tmp_366 = ldq_27_bits_uop_xcpt_ma_if;
      5'b11100:
        casez_tmp_366 = ldq_28_bits_uop_xcpt_ma_if;
      5'b11101:
        casez_tmp_366 = ldq_29_bits_uop_xcpt_ma_if;
      5'b11110:
        casez_tmp_366 = ldq_30_bits_uop_xcpt_ma_if;
      default:
        casez_tmp_366 = ldq_31_bits_uop_xcpt_ma_if;
    endcase
  end // always @(*)
  reg         casez_tmp_367;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_367 = ldq_0_bits_uop_bp_debug_if;
      5'b00001:
        casez_tmp_367 = ldq_1_bits_uop_bp_debug_if;
      5'b00010:
        casez_tmp_367 = ldq_2_bits_uop_bp_debug_if;
      5'b00011:
        casez_tmp_367 = ldq_3_bits_uop_bp_debug_if;
      5'b00100:
        casez_tmp_367 = ldq_4_bits_uop_bp_debug_if;
      5'b00101:
        casez_tmp_367 = ldq_5_bits_uop_bp_debug_if;
      5'b00110:
        casez_tmp_367 = ldq_6_bits_uop_bp_debug_if;
      5'b00111:
        casez_tmp_367 = ldq_7_bits_uop_bp_debug_if;
      5'b01000:
        casez_tmp_367 = ldq_8_bits_uop_bp_debug_if;
      5'b01001:
        casez_tmp_367 = ldq_9_bits_uop_bp_debug_if;
      5'b01010:
        casez_tmp_367 = ldq_10_bits_uop_bp_debug_if;
      5'b01011:
        casez_tmp_367 = ldq_11_bits_uop_bp_debug_if;
      5'b01100:
        casez_tmp_367 = ldq_12_bits_uop_bp_debug_if;
      5'b01101:
        casez_tmp_367 = ldq_13_bits_uop_bp_debug_if;
      5'b01110:
        casez_tmp_367 = ldq_14_bits_uop_bp_debug_if;
      5'b01111:
        casez_tmp_367 = ldq_15_bits_uop_bp_debug_if;
      5'b10000:
        casez_tmp_367 = ldq_16_bits_uop_bp_debug_if;
      5'b10001:
        casez_tmp_367 = ldq_17_bits_uop_bp_debug_if;
      5'b10010:
        casez_tmp_367 = ldq_18_bits_uop_bp_debug_if;
      5'b10011:
        casez_tmp_367 = ldq_19_bits_uop_bp_debug_if;
      5'b10100:
        casez_tmp_367 = ldq_20_bits_uop_bp_debug_if;
      5'b10101:
        casez_tmp_367 = ldq_21_bits_uop_bp_debug_if;
      5'b10110:
        casez_tmp_367 = ldq_22_bits_uop_bp_debug_if;
      5'b10111:
        casez_tmp_367 = ldq_23_bits_uop_bp_debug_if;
      5'b11000:
        casez_tmp_367 = ldq_24_bits_uop_bp_debug_if;
      5'b11001:
        casez_tmp_367 = ldq_25_bits_uop_bp_debug_if;
      5'b11010:
        casez_tmp_367 = ldq_26_bits_uop_bp_debug_if;
      5'b11011:
        casez_tmp_367 = ldq_27_bits_uop_bp_debug_if;
      5'b11100:
        casez_tmp_367 = ldq_28_bits_uop_bp_debug_if;
      5'b11101:
        casez_tmp_367 = ldq_29_bits_uop_bp_debug_if;
      5'b11110:
        casez_tmp_367 = ldq_30_bits_uop_bp_debug_if;
      default:
        casez_tmp_367 = ldq_31_bits_uop_bp_debug_if;
    endcase
  end // always @(*)
  reg         casez_tmp_368;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_368 = ldq_0_bits_uop_bp_xcpt_if;
      5'b00001:
        casez_tmp_368 = ldq_1_bits_uop_bp_xcpt_if;
      5'b00010:
        casez_tmp_368 = ldq_2_bits_uop_bp_xcpt_if;
      5'b00011:
        casez_tmp_368 = ldq_3_bits_uop_bp_xcpt_if;
      5'b00100:
        casez_tmp_368 = ldq_4_bits_uop_bp_xcpt_if;
      5'b00101:
        casez_tmp_368 = ldq_5_bits_uop_bp_xcpt_if;
      5'b00110:
        casez_tmp_368 = ldq_6_bits_uop_bp_xcpt_if;
      5'b00111:
        casez_tmp_368 = ldq_7_bits_uop_bp_xcpt_if;
      5'b01000:
        casez_tmp_368 = ldq_8_bits_uop_bp_xcpt_if;
      5'b01001:
        casez_tmp_368 = ldq_9_bits_uop_bp_xcpt_if;
      5'b01010:
        casez_tmp_368 = ldq_10_bits_uop_bp_xcpt_if;
      5'b01011:
        casez_tmp_368 = ldq_11_bits_uop_bp_xcpt_if;
      5'b01100:
        casez_tmp_368 = ldq_12_bits_uop_bp_xcpt_if;
      5'b01101:
        casez_tmp_368 = ldq_13_bits_uop_bp_xcpt_if;
      5'b01110:
        casez_tmp_368 = ldq_14_bits_uop_bp_xcpt_if;
      5'b01111:
        casez_tmp_368 = ldq_15_bits_uop_bp_xcpt_if;
      5'b10000:
        casez_tmp_368 = ldq_16_bits_uop_bp_xcpt_if;
      5'b10001:
        casez_tmp_368 = ldq_17_bits_uop_bp_xcpt_if;
      5'b10010:
        casez_tmp_368 = ldq_18_bits_uop_bp_xcpt_if;
      5'b10011:
        casez_tmp_368 = ldq_19_bits_uop_bp_xcpt_if;
      5'b10100:
        casez_tmp_368 = ldq_20_bits_uop_bp_xcpt_if;
      5'b10101:
        casez_tmp_368 = ldq_21_bits_uop_bp_xcpt_if;
      5'b10110:
        casez_tmp_368 = ldq_22_bits_uop_bp_xcpt_if;
      5'b10111:
        casez_tmp_368 = ldq_23_bits_uop_bp_xcpt_if;
      5'b11000:
        casez_tmp_368 = ldq_24_bits_uop_bp_xcpt_if;
      5'b11001:
        casez_tmp_368 = ldq_25_bits_uop_bp_xcpt_if;
      5'b11010:
        casez_tmp_368 = ldq_26_bits_uop_bp_xcpt_if;
      5'b11011:
        casez_tmp_368 = ldq_27_bits_uop_bp_xcpt_if;
      5'b11100:
        casez_tmp_368 = ldq_28_bits_uop_bp_xcpt_if;
      5'b11101:
        casez_tmp_368 = ldq_29_bits_uop_bp_xcpt_if;
      5'b11110:
        casez_tmp_368 = ldq_30_bits_uop_bp_xcpt_if;
      default:
        casez_tmp_368 = ldq_31_bits_uop_bp_xcpt_if;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_369;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_369 = ldq_0_bits_uop_debug_fsrc;
      5'b00001:
        casez_tmp_369 = ldq_1_bits_uop_debug_fsrc;
      5'b00010:
        casez_tmp_369 = ldq_2_bits_uop_debug_fsrc;
      5'b00011:
        casez_tmp_369 = ldq_3_bits_uop_debug_fsrc;
      5'b00100:
        casez_tmp_369 = ldq_4_bits_uop_debug_fsrc;
      5'b00101:
        casez_tmp_369 = ldq_5_bits_uop_debug_fsrc;
      5'b00110:
        casez_tmp_369 = ldq_6_bits_uop_debug_fsrc;
      5'b00111:
        casez_tmp_369 = ldq_7_bits_uop_debug_fsrc;
      5'b01000:
        casez_tmp_369 = ldq_8_bits_uop_debug_fsrc;
      5'b01001:
        casez_tmp_369 = ldq_9_bits_uop_debug_fsrc;
      5'b01010:
        casez_tmp_369 = ldq_10_bits_uop_debug_fsrc;
      5'b01011:
        casez_tmp_369 = ldq_11_bits_uop_debug_fsrc;
      5'b01100:
        casez_tmp_369 = ldq_12_bits_uop_debug_fsrc;
      5'b01101:
        casez_tmp_369 = ldq_13_bits_uop_debug_fsrc;
      5'b01110:
        casez_tmp_369 = ldq_14_bits_uop_debug_fsrc;
      5'b01111:
        casez_tmp_369 = ldq_15_bits_uop_debug_fsrc;
      5'b10000:
        casez_tmp_369 = ldq_16_bits_uop_debug_fsrc;
      5'b10001:
        casez_tmp_369 = ldq_17_bits_uop_debug_fsrc;
      5'b10010:
        casez_tmp_369 = ldq_18_bits_uop_debug_fsrc;
      5'b10011:
        casez_tmp_369 = ldq_19_bits_uop_debug_fsrc;
      5'b10100:
        casez_tmp_369 = ldq_20_bits_uop_debug_fsrc;
      5'b10101:
        casez_tmp_369 = ldq_21_bits_uop_debug_fsrc;
      5'b10110:
        casez_tmp_369 = ldq_22_bits_uop_debug_fsrc;
      5'b10111:
        casez_tmp_369 = ldq_23_bits_uop_debug_fsrc;
      5'b11000:
        casez_tmp_369 = ldq_24_bits_uop_debug_fsrc;
      5'b11001:
        casez_tmp_369 = ldq_25_bits_uop_debug_fsrc;
      5'b11010:
        casez_tmp_369 = ldq_26_bits_uop_debug_fsrc;
      5'b11011:
        casez_tmp_369 = ldq_27_bits_uop_debug_fsrc;
      5'b11100:
        casez_tmp_369 = ldq_28_bits_uop_debug_fsrc;
      5'b11101:
        casez_tmp_369 = ldq_29_bits_uop_debug_fsrc;
      5'b11110:
        casez_tmp_369 = ldq_30_bits_uop_debug_fsrc;
      default:
        casez_tmp_369 = ldq_31_bits_uop_debug_fsrc;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_370;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_370 = ldq_0_bits_uop_debug_tsrc;
      5'b00001:
        casez_tmp_370 = ldq_1_bits_uop_debug_tsrc;
      5'b00010:
        casez_tmp_370 = ldq_2_bits_uop_debug_tsrc;
      5'b00011:
        casez_tmp_370 = ldq_3_bits_uop_debug_tsrc;
      5'b00100:
        casez_tmp_370 = ldq_4_bits_uop_debug_tsrc;
      5'b00101:
        casez_tmp_370 = ldq_5_bits_uop_debug_tsrc;
      5'b00110:
        casez_tmp_370 = ldq_6_bits_uop_debug_tsrc;
      5'b00111:
        casez_tmp_370 = ldq_7_bits_uop_debug_tsrc;
      5'b01000:
        casez_tmp_370 = ldq_8_bits_uop_debug_tsrc;
      5'b01001:
        casez_tmp_370 = ldq_9_bits_uop_debug_tsrc;
      5'b01010:
        casez_tmp_370 = ldq_10_bits_uop_debug_tsrc;
      5'b01011:
        casez_tmp_370 = ldq_11_bits_uop_debug_tsrc;
      5'b01100:
        casez_tmp_370 = ldq_12_bits_uop_debug_tsrc;
      5'b01101:
        casez_tmp_370 = ldq_13_bits_uop_debug_tsrc;
      5'b01110:
        casez_tmp_370 = ldq_14_bits_uop_debug_tsrc;
      5'b01111:
        casez_tmp_370 = ldq_15_bits_uop_debug_tsrc;
      5'b10000:
        casez_tmp_370 = ldq_16_bits_uop_debug_tsrc;
      5'b10001:
        casez_tmp_370 = ldq_17_bits_uop_debug_tsrc;
      5'b10010:
        casez_tmp_370 = ldq_18_bits_uop_debug_tsrc;
      5'b10011:
        casez_tmp_370 = ldq_19_bits_uop_debug_tsrc;
      5'b10100:
        casez_tmp_370 = ldq_20_bits_uop_debug_tsrc;
      5'b10101:
        casez_tmp_370 = ldq_21_bits_uop_debug_tsrc;
      5'b10110:
        casez_tmp_370 = ldq_22_bits_uop_debug_tsrc;
      5'b10111:
        casez_tmp_370 = ldq_23_bits_uop_debug_tsrc;
      5'b11000:
        casez_tmp_370 = ldq_24_bits_uop_debug_tsrc;
      5'b11001:
        casez_tmp_370 = ldq_25_bits_uop_debug_tsrc;
      5'b11010:
        casez_tmp_370 = ldq_26_bits_uop_debug_tsrc;
      5'b11011:
        casez_tmp_370 = ldq_27_bits_uop_debug_tsrc;
      5'b11100:
        casez_tmp_370 = ldq_28_bits_uop_debug_tsrc;
      5'b11101:
        casez_tmp_370 = ldq_29_bits_uop_debug_tsrc;
      5'b11110:
        casez_tmp_370 = ldq_30_bits_uop_debug_tsrc;
      default:
        casez_tmp_370 = ldq_31_bits_uop_debug_tsrc;
    endcase
  end // always @(*)
  reg         casez_tmp_371;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_371 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_371 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_371 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_371 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_371 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_371 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_371 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_371 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_371 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_371 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_371 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_371 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_371 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_371 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_371 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_371 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_371 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_371 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_371 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_371 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_371 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_371 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_371 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_371 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_371 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_371 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_371 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_371 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_371 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_371 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_371 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_371 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg  [39:0] casez_tmp_372;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_372 = ldq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_372 = ldq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_372 = ldq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_372 = ldq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_372 = ldq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_372 = ldq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_372 = ldq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_372 = ldq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_372 = ldq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_372 = ldq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_372 = ldq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_372 = ldq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_372 = ldq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_372 = ldq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_372 = ldq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_372 = ldq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_372 = ldq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_372 = ldq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_372 = ldq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_372 = ldq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_372 = ldq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_372 = ldq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_372 = ldq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_372 = ldq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_372 = ldq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_372 = ldq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_372 = ldq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_372 = ldq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_372 = ldq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_372 = ldq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_372 = ldq_30_bits_addr_bits;
      default:
        casez_tmp_372 = ldq_31_bits_addr_bits;
    endcase
  end // always @(*)
  reg         casez_tmp_373;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_373 = ldq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_373 = ldq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_373 = ldq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_373 = ldq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_373 = ldq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_373 = ldq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_373 = ldq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_373 = ldq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_373 = ldq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_373 = ldq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_373 = ldq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_373 = ldq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_373 = ldq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_373 = ldq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_373 = ldq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_373 = ldq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_373 = ldq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_373 = ldq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_373 = ldq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_373 = ldq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_373 = ldq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_373 = ldq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_373 = ldq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_373 = ldq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_373 = ldq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_373 = ldq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_373 = ldq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_373 = ldq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_373 = ldq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_373 = ldq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_373 = ldq_30_bits_addr_is_virtual;
      default:
        casez_tmp_373 = ldq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         casez_tmp_374;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_374 = ldq_0_bits_addr_is_uncacheable;
      5'b00001:
        casez_tmp_374 = ldq_1_bits_addr_is_uncacheable;
      5'b00010:
        casez_tmp_374 = ldq_2_bits_addr_is_uncacheable;
      5'b00011:
        casez_tmp_374 = ldq_3_bits_addr_is_uncacheable;
      5'b00100:
        casez_tmp_374 = ldq_4_bits_addr_is_uncacheable;
      5'b00101:
        casez_tmp_374 = ldq_5_bits_addr_is_uncacheable;
      5'b00110:
        casez_tmp_374 = ldq_6_bits_addr_is_uncacheable;
      5'b00111:
        casez_tmp_374 = ldq_7_bits_addr_is_uncacheable;
      5'b01000:
        casez_tmp_374 = ldq_8_bits_addr_is_uncacheable;
      5'b01001:
        casez_tmp_374 = ldq_9_bits_addr_is_uncacheable;
      5'b01010:
        casez_tmp_374 = ldq_10_bits_addr_is_uncacheable;
      5'b01011:
        casez_tmp_374 = ldq_11_bits_addr_is_uncacheable;
      5'b01100:
        casez_tmp_374 = ldq_12_bits_addr_is_uncacheable;
      5'b01101:
        casez_tmp_374 = ldq_13_bits_addr_is_uncacheable;
      5'b01110:
        casez_tmp_374 = ldq_14_bits_addr_is_uncacheable;
      5'b01111:
        casez_tmp_374 = ldq_15_bits_addr_is_uncacheable;
      5'b10000:
        casez_tmp_374 = ldq_16_bits_addr_is_uncacheable;
      5'b10001:
        casez_tmp_374 = ldq_17_bits_addr_is_uncacheable;
      5'b10010:
        casez_tmp_374 = ldq_18_bits_addr_is_uncacheable;
      5'b10011:
        casez_tmp_374 = ldq_19_bits_addr_is_uncacheable;
      5'b10100:
        casez_tmp_374 = ldq_20_bits_addr_is_uncacheable;
      5'b10101:
        casez_tmp_374 = ldq_21_bits_addr_is_uncacheable;
      5'b10110:
        casez_tmp_374 = ldq_22_bits_addr_is_uncacheable;
      5'b10111:
        casez_tmp_374 = ldq_23_bits_addr_is_uncacheable;
      5'b11000:
        casez_tmp_374 = ldq_24_bits_addr_is_uncacheable;
      5'b11001:
        casez_tmp_374 = ldq_25_bits_addr_is_uncacheable;
      5'b11010:
        casez_tmp_374 = ldq_26_bits_addr_is_uncacheable;
      5'b11011:
        casez_tmp_374 = ldq_27_bits_addr_is_uncacheable;
      5'b11100:
        casez_tmp_374 = ldq_28_bits_addr_is_uncacheable;
      5'b11101:
        casez_tmp_374 = ldq_29_bits_addr_is_uncacheable;
      5'b11110:
        casez_tmp_374 = ldq_30_bits_addr_is_uncacheable;
      default:
        casez_tmp_374 = ldq_31_bits_addr_is_uncacheable;
    endcase
  end // always @(*)
  reg         casez_tmp_375;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_375 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_375 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_375 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_375 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_375 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_375 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_375 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_375 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_375 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_375 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_375 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_375 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_375 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_375 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_375 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_375 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_375 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_375 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_375 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_375 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_375 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_375 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_375 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_375 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_375 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_375 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_375 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_375 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_375 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_375 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_375 = ldq_30_bits_executed;
      default:
        casez_tmp_375 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg         casez_tmp_376;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_376 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_376 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_376 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_376 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_376 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_376 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_376 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_376 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_376 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_376 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_376 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_376 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_376 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_376 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_376 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_376 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_376 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_376 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_376 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_376 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_376 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_376 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_376 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_376 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_376 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_376 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_376 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_376 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_376 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_376 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_376 = ldq_30_bits_succeeded;
      default:
        casez_tmp_376 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  reg         casez_tmp_377;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_377 = ldq_0_bits_order_fail;
      5'b00001:
        casez_tmp_377 = ldq_1_bits_order_fail;
      5'b00010:
        casez_tmp_377 = ldq_2_bits_order_fail;
      5'b00011:
        casez_tmp_377 = ldq_3_bits_order_fail;
      5'b00100:
        casez_tmp_377 = ldq_4_bits_order_fail;
      5'b00101:
        casez_tmp_377 = ldq_5_bits_order_fail;
      5'b00110:
        casez_tmp_377 = ldq_6_bits_order_fail;
      5'b00111:
        casez_tmp_377 = ldq_7_bits_order_fail;
      5'b01000:
        casez_tmp_377 = ldq_8_bits_order_fail;
      5'b01001:
        casez_tmp_377 = ldq_9_bits_order_fail;
      5'b01010:
        casez_tmp_377 = ldq_10_bits_order_fail;
      5'b01011:
        casez_tmp_377 = ldq_11_bits_order_fail;
      5'b01100:
        casez_tmp_377 = ldq_12_bits_order_fail;
      5'b01101:
        casez_tmp_377 = ldq_13_bits_order_fail;
      5'b01110:
        casez_tmp_377 = ldq_14_bits_order_fail;
      5'b01111:
        casez_tmp_377 = ldq_15_bits_order_fail;
      5'b10000:
        casez_tmp_377 = ldq_16_bits_order_fail;
      5'b10001:
        casez_tmp_377 = ldq_17_bits_order_fail;
      5'b10010:
        casez_tmp_377 = ldq_18_bits_order_fail;
      5'b10011:
        casez_tmp_377 = ldq_19_bits_order_fail;
      5'b10100:
        casez_tmp_377 = ldq_20_bits_order_fail;
      5'b10101:
        casez_tmp_377 = ldq_21_bits_order_fail;
      5'b10110:
        casez_tmp_377 = ldq_22_bits_order_fail;
      5'b10111:
        casez_tmp_377 = ldq_23_bits_order_fail;
      5'b11000:
        casez_tmp_377 = ldq_24_bits_order_fail;
      5'b11001:
        casez_tmp_377 = ldq_25_bits_order_fail;
      5'b11010:
        casez_tmp_377 = ldq_26_bits_order_fail;
      5'b11011:
        casez_tmp_377 = ldq_27_bits_order_fail;
      5'b11100:
        casez_tmp_377 = ldq_28_bits_order_fail;
      5'b11101:
        casez_tmp_377 = ldq_29_bits_order_fail;
      5'b11110:
        casez_tmp_377 = ldq_30_bits_order_fail;
      default:
        casez_tmp_377 = ldq_31_bits_order_fail;
    endcase
  end // always @(*)
  reg  [31:0] casez_tmp_378;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_378 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_378 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_378 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_378 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_378 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_378 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_378 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_378 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_378 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_378 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_378 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_378 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_378 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_378 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_378 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_378 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_378 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_378 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_378 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_378 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_378 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_378 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_378 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_378 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_378 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_378 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_378 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_378 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_378 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_378 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_378 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_378 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  reg         casez_tmp_379;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_379 = p1_block_load_mask_0;
      5'b00001:
        casez_tmp_379 = p1_block_load_mask_1;
      5'b00010:
        casez_tmp_379 = p1_block_load_mask_2;
      5'b00011:
        casez_tmp_379 = p1_block_load_mask_3;
      5'b00100:
        casez_tmp_379 = p1_block_load_mask_4;
      5'b00101:
        casez_tmp_379 = p1_block_load_mask_5;
      5'b00110:
        casez_tmp_379 = p1_block_load_mask_6;
      5'b00111:
        casez_tmp_379 = p1_block_load_mask_7;
      5'b01000:
        casez_tmp_379 = p1_block_load_mask_8;
      5'b01001:
        casez_tmp_379 = p1_block_load_mask_9;
      5'b01010:
        casez_tmp_379 = p1_block_load_mask_10;
      5'b01011:
        casez_tmp_379 = p1_block_load_mask_11;
      5'b01100:
        casez_tmp_379 = p1_block_load_mask_12;
      5'b01101:
        casez_tmp_379 = p1_block_load_mask_13;
      5'b01110:
        casez_tmp_379 = p1_block_load_mask_14;
      5'b01111:
        casez_tmp_379 = p1_block_load_mask_15;
      5'b10000:
        casez_tmp_379 = p1_block_load_mask_16;
      5'b10001:
        casez_tmp_379 = p1_block_load_mask_17;
      5'b10010:
        casez_tmp_379 = p1_block_load_mask_18;
      5'b10011:
        casez_tmp_379 = p1_block_load_mask_19;
      5'b10100:
        casez_tmp_379 = p1_block_load_mask_20;
      5'b10101:
        casez_tmp_379 = p1_block_load_mask_21;
      5'b10110:
        casez_tmp_379 = p1_block_load_mask_22;
      5'b10111:
        casez_tmp_379 = p1_block_load_mask_23;
      5'b11000:
        casez_tmp_379 = p1_block_load_mask_24;
      5'b11001:
        casez_tmp_379 = p1_block_load_mask_25;
      5'b11010:
        casez_tmp_379 = p1_block_load_mask_26;
      5'b11011:
        casez_tmp_379 = p1_block_load_mask_27;
      5'b11100:
        casez_tmp_379 = p1_block_load_mask_28;
      5'b11101:
        casez_tmp_379 = p1_block_load_mask_29;
      5'b11110:
        casez_tmp_379 = p1_block_load_mask_30;
      default:
        casez_tmp_379 = p1_block_load_mask_31;
    endcase
  end // always @(*)
  reg         casez_tmp_380;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_380 = p2_block_load_mask_0;
      5'b00001:
        casez_tmp_380 = p2_block_load_mask_1;
      5'b00010:
        casez_tmp_380 = p2_block_load_mask_2;
      5'b00011:
        casez_tmp_380 = p2_block_load_mask_3;
      5'b00100:
        casez_tmp_380 = p2_block_load_mask_4;
      5'b00101:
        casez_tmp_380 = p2_block_load_mask_5;
      5'b00110:
        casez_tmp_380 = p2_block_load_mask_6;
      5'b00111:
        casez_tmp_380 = p2_block_load_mask_7;
      5'b01000:
        casez_tmp_380 = p2_block_load_mask_8;
      5'b01001:
        casez_tmp_380 = p2_block_load_mask_9;
      5'b01010:
        casez_tmp_380 = p2_block_load_mask_10;
      5'b01011:
        casez_tmp_380 = p2_block_load_mask_11;
      5'b01100:
        casez_tmp_380 = p2_block_load_mask_12;
      5'b01101:
        casez_tmp_380 = p2_block_load_mask_13;
      5'b01110:
        casez_tmp_380 = p2_block_load_mask_14;
      5'b01111:
        casez_tmp_380 = p2_block_load_mask_15;
      5'b10000:
        casez_tmp_380 = p2_block_load_mask_16;
      5'b10001:
        casez_tmp_380 = p2_block_load_mask_17;
      5'b10010:
        casez_tmp_380 = p2_block_load_mask_18;
      5'b10011:
        casez_tmp_380 = p2_block_load_mask_19;
      5'b10100:
        casez_tmp_380 = p2_block_load_mask_20;
      5'b10101:
        casez_tmp_380 = p2_block_load_mask_21;
      5'b10110:
        casez_tmp_380 = p2_block_load_mask_22;
      5'b10111:
        casez_tmp_380 = p2_block_load_mask_23;
      5'b11000:
        casez_tmp_380 = p2_block_load_mask_24;
      5'b11001:
        casez_tmp_380 = p2_block_load_mask_25;
      5'b11010:
        casez_tmp_380 = p2_block_load_mask_26;
      5'b11011:
        casez_tmp_380 = p2_block_load_mask_27;
      5'b11100:
        casez_tmp_380 = p2_block_load_mask_28;
      5'b11101:
        casez_tmp_380 = p2_block_load_mask_29;
      5'b11110:
        casez_tmp_380 = p2_block_load_mask_30;
      default:
        casez_tmp_380 = p2_block_load_mask_31;
    endcase
  end // always @(*)
  wire        will_fire_stad_incoming_0_will_fire = _can_fire_sta_incoming_T & exe_req_0_bits_uop_ctrl_is_std & ~will_fire_load_incoming_0_will_fire & ~will_fire_load_incoming_0_will_fire;
  wire        _will_fire_sta_incoming_0_will_fire_T_2 = ~will_fire_load_incoming_0_will_fire & ~will_fire_stad_incoming_0_will_fire;
  wire        will_fire_sta_incoming_0_will_fire = _can_fire_sta_incoming_T & ~exe_req_0_bits_uop_ctrl_is_std & _will_fire_sta_incoming_0_will_fire_T_2 & ~will_fire_load_incoming_0_will_fire & ~will_fire_stad_incoming_0_will_fire & ~will_fire_stad_incoming_0_will_fire;
  wire        _will_fire_sfence_0_will_fire_T_2 = _will_fire_sta_incoming_0_will_fire_T_2 & ~will_fire_sta_incoming_0_will_fire;
  wire        _will_fire_std_incoming_0_will_fire_T_14 = ~will_fire_stad_incoming_0_will_fire & ~will_fire_sta_incoming_0_will_fire;
  wire        will_fire_std_incoming_0_will_fire = can_fire_std_incoming_0 & _will_fire_std_incoming_0_will_fire_T_14;
  wire        will_fire_sfence_0_will_fire = exe_req_0_valid & exe_req_0_bits_sfence_valid & _will_fire_sfence_0_will_fire_T_2 & _will_fire_std_incoming_0_will_fire_T_14 & ~will_fire_std_incoming_0_will_fire;
  assign _will_fire_store_commit_0_T_2 = _will_fire_sfence_0_will_fire_T_2 & ~will_fire_sfence_0_will_fire & ~will_fire_hella_incoming_0_will_fire & ~will_fire_load_retry_0_will_fire & ~will_fire_sta_retry_0_will_fire;
  wire        will_fire_store_commit_0_will_fire = casez_tmp & ~casez_tmp_52 & ~mem_xcpt_valid & ~casez_tmp_46 & (casez_tmp_84 | casez_tmp_54 & casez_tmp_79 & ~casez_tmp_81 & casez_tmp_82) & ~will_fire_load_incoming_0_will_fire & ~will_fire_hella_incoming_0_will_fire & ~will_fire_hella_wakeup_0_will_fire & ~will_fire_load_retry_0_will_fire & ~will_fire_load_wakeup_0_will_fire;
  wire        _exe_cmd_T = will_fire_load_incoming_0_will_fire | will_fire_stad_incoming_0_will_fire;
  wire        _GEN_18 = _exe_cmd_T | will_fire_sta_incoming_0_will_fire;
  wire        _GEN_19 = ldq_wakeup_idx == 5'h0;
  wire        _GEN_20 = ldq_wakeup_idx == 5'h1;
  wire        _GEN_21 = ldq_wakeup_idx == 5'h2;
  wire        _GEN_22 = ldq_wakeup_idx == 5'h3;
  wire        _GEN_23 = ldq_wakeup_idx == 5'h4;
  wire        _GEN_24 = ldq_wakeup_idx == 5'h5;
  wire        _GEN_25 = ldq_wakeup_idx == 5'h6;
  wire        _GEN_26 = ldq_wakeup_idx == 5'h7;
  wire        _GEN_27 = ldq_wakeup_idx == 5'h8;
  wire        _GEN_28 = ldq_wakeup_idx == 5'h9;
  wire        _GEN_29 = ldq_wakeup_idx == 5'hA;
  wire        _GEN_30 = ldq_wakeup_idx == 5'hB;
  wire        _GEN_31 = ldq_wakeup_idx == 5'hC;
  wire        _GEN_32 = ldq_wakeup_idx == 5'hD;
  wire        _GEN_33 = ldq_wakeup_idx == 5'hE;
  wire        _GEN_34 = ldq_wakeup_idx == 5'hF;
  wire        _GEN_35 = ldq_wakeup_idx == 5'h10;
  wire        _GEN_36 = ldq_wakeup_idx == 5'h11;
  wire        _GEN_37 = ldq_wakeup_idx == 5'h12;
  wire        _GEN_38 = ldq_wakeup_idx == 5'h13;
  wire        _GEN_39 = ldq_wakeup_idx == 5'h14;
  wire        _GEN_40 = ldq_wakeup_idx == 5'h15;
  wire        _GEN_41 = ldq_wakeup_idx == 5'h16;
  wire        _GEN_42 = ldq_wakeup_idx == 5'h17;
  wire        _GEN_43 = ldq_wakeup_idx == 5'h18;
  wire        _GEN_44 = ldq_wakeup_idx == 5'h19;
  wire        _GEN_45 = ldq_wakeup_idx == 5'h1A;
  wire        _GEN_46 = ldq_wakeup_idx == 5'h1B;
  wire        _GEN_47 = ldq_wakeup_idx == 5'h1C;
  wire        _GEN_48 = ldq_wakeup_idx == 5'h1D;
  wire        _GEN_49 = ldq_wakeup_idx == 5'h1E;
  wire        _GEN_50 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h0;
  wire        _GEN_51 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h1;
  wire        _GEN_52 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h2;
  wire        _GEN_53 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h3;
  wire        _GEN_54 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h4;
  wire        _GEN_55 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h5;
  wire        _GEN_56 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h6;
  wire        _GEN_57 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h7;
  wire        _GEN_58 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h8;
  wire        _GEN_59 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h9;
  wire        _GEN_60 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'hA;
  wire        _GEN_61 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'hB;
  wire        _GEN_62 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'hC;
  wire        _GEN_63 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'hD;
  wire        _GEN_64 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'hE;
  wire        _GEN_65 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'hF;
  wire        _GEN_66 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h10;
  wire        _GEN_67 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h11;
  wire        _GEN_68 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h12;
  wire        _GEN_69 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h13;
  wire        _GEN_70 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h14;
  wire        _GEN_71 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h15;
  wire        _GEN_72 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h16;
  wire        _GEN_73 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h17;
  wire        _GEN_74 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h18;
  wire        _GEN_75 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h19;
  wire        _GEN_76 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h1A;
  wire        _GEN_77 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h1B;
  wire        _GEN_78 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h1C;
  wire        _GEN_79 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h1D;
  wire        _GEN_80 = _mem_incoming_uop_WIRE_0_ldq_idx == 5'h1E;
  wire        _GEN_81 = ldq_retry_idx == 5'h0;
  wire        _GEN_82 = will_fire_load_wakeup_0_will_fire ? _GEN_19 : will_fire_load_incoming_0_will_fire ? _GEN_50 : will_fire_load_retry_0_will_fire & _GEN_81;
  wire        _GEN_83 = ldq_retry_idx == 5'h1;
  wire        _GEN_84 = will_fire_load_wakeup_0_will_fire ? _GEN_20 : will_fire_load_incoming_0_will_fire ? _GEN_51 : will_fire_load_retry_0_will_fire & _GEN_83;
  wire        _GEN_85 = ldq_retry_idx == 5'h2;
  wire        _GEN_86 = will_fire_load_wakeup_0_will_fire ? _GEN_21 : will_fire_load_incoming_0_will_fire ? _GEN_52 : will_fire_load_retry_0_will_fire & _GEN_85;
  wire        _GEN_87 = ldq_retry_idx == 5'h3;
  wire        _GEN_88 = will_fire_load_wakeup_0_will_fire ? _GEN_22 : will_fire_load_incoming_0_will_fire ? _GEN_53 : will_fire_load_retry_0_will_fire & _GEN_87;
  wire        _GEN_89 = ldq_retry_idx == 5'h4;
  wire        _GEN_90 = will_fire_load_wakeup_0_will_fire ? _GEN_23 : will_fire_load_incoming_0_will_fire ? _GEN_54 : will_fire_load_retry_0_will_fire & _GEN_89;
  wire        _GEN_91 = ldq_retry_idx == 5'h5;
  wire        _GEN_92 = will_fire_load_wakeup_0_will_fire ? _GEN_24 : will_fire_load_incoming_0_will_fire ? _GEN_55 : will_fire_load_retry_0_will_fire & _GEN_91;
  wire        _GEN_93 = ldq_retry_idx == 5'h6;
  wire        _GEN_94 = will_fire_load_wakeup_0_will_fire ? _GEN_25 : will_fire_load_incoming_0_will_fire ? _GEN_56 : will_fire_load_retry_0_will_fire & _GEN_93;
  wire        _GEN_95 = ldq_retry_idx == 5'h7;
  wire        _GEN_96 = will_fire_load_wakeup_0_will_fire ? _GEN_26 : will_fire_load_incoming_0_will_fire ? _GEN_57 : will_fire_load_retry_0_will_fire & _GEN_95;
  wire        _GEN_97 = ldq_retry_idx == 5'h8;
  wire        _GEN_98 = will_fire_load_wakeup_0_will_fire ? _GEN_27 : will_fire_load_incoming_0_will_fire ? _GEN_58 : will_fire_load_retry_0_will_fire & _GEN_97;
  wire        _GEN_99 = ldq_retry_idx == 5'h9;
  wire        _GEN_100 = will_fire_load_wakeup_0_will_fire ? _GEN_28 : will_fire_load_incoming_0_will_fire ? _GEN_59 : will_fire_load_retry_0_will_fire & _GEN_99;
  wire        _GEN_101 = ldq_retry_idx == 5'hA;
  wire        _GEN_102 = will_fire_load_wakeup_0_will_fire ? _GEN_29 : will_fire_load_incoming_0_will_fire ? _GEN_60 : will_fire_load_retry_0_will_fire & _GEN_101;
  wire        _GEN_103 = ldq_retry_idx == 5'hB;
  wire        _GEN_104 = will_fire_load_wakeup_0_will_fire ? _GEN_30 : will_fire_load_incoming_0_will_fire ? _GEN_61 : will_fire_load_retry_0_will_fire & _GEN_103;
  wire        _GEN_105 = ldq_retry_idx == 5'hC;
  wire        _GEN_106 = will_fire_load_wakeup_0_will_fire ? _GEN_31 : will_fire_load_incoming_0_will_fire ? _GEN_62 : will_fire_load_retry_0_will_fire & _GEN_105;
  wire        _GEN_107 = ldq_retry_idx == 5'hD;
  wire        _GEN_108 = will_fire_load_wakeup_0_will_fire ? _GEN_32 : will_fire_load_incoming_0_will_fire ? _GEN_63 : will_fire_load_retry_0_will_fire & _GEN_107;
  wire        _GEN_109 = ldq_retry_idx == 5'hE;
  wire        _GEN_110 = will_fire_load_wakeup_0_will_fire ? _GEN_33 : will_fire_load_incoming_0_will_fire ? _GEN_64 : will_fire_load_retry_0_will_fire & _GEN_109;
  wire        _GEN_111 = ldq_retry_idx == 5'hF;
  wire        _GEN_112 = will_fire_load_wakeup_0_will_fire ? _GEN_34 : will_fire_load_incoming_0_will_fire ? _GEN_65 : will_fire_load_retry_0_will_fire & _GEN_111;
  wire        _GEN_113 = ldq_retry_idx == 5'h10;
  wire        _GEN_114 = will_fire_load_wakeup_0_will_fire ? _GEN_35 : will_fire_load_incoming_0_will_fire ? _GEN_66 : will_fire_load_retry_0_will_fire & _GEN_113;
  wire        _GEN_115 = ldq_retry_idx == 5'h11;
  wire        _GEN_116 = will_fire_load_wakeup_0_will_fire ? _GEN_36 : will_fire_load_incoming_0_will_fire ? _GEN_67 : will_fire_load_retry_0_will_fire & _GEN_115;
  wire        _GEN_117 = ldq_retry_idx == 5'h12;
  wire        _GEN_118 = will_fire_load_wakeup_0_will_fire ? _GEN_37 : will_fire_load_incoming_0_will_fire ? _GEN_68 : will_fire_load_retry_0_will_fire & _GEN_117;
  wire        _GEN_119 = ldq_retry_idx == 5'h13;
  wire        _GEN_120 = will_fire_load_wakeup_0_will_fire ? _GEN_38 : will_fire_load_incoming_0_will_fire ? _GEN_69 : will_fire_load_retry_0_will_fire & _GEN_119;
  wire        _GEN_121 = ldq_retry_idx == 5'h14;
  wire        _GEN_122 = will_fire_load_wakeup_0_will_fire ? _GEN_39 : will_fire_load_incoming_0_will_fire ? _GEN_70 : will_fire_load_retry_0_will_fire & _GEN_121;
  wire        _GEN_123 = ldq_retry_idx == 5'h15;
  wire        _GEN_124 = will_fire_load_wakeup_0_will_fire ? _GEN_40 : will_fire_load_incoming_0_will_fire ? _GEN_71 : will_fire_load_retry_0_will_fire & _GEN_123;
  wire        _GEN_125 = ldq_retry_idx == 5'h16;
  wire        _GEN_126 = will_fire_load_wakeup_0_will_fire ? _GEN_41 : will_fire_load_incoming_0_will_fire ? _GEN_72 : will_fire_load_retry_0_will_fire & _GEN_125;
  wire        _GEN_127 = ldq_retry_idx == 5'h17;
  wire        _GEN_128 = will_fire_load_wakeup_0_will_fire ? _GEN_42 : will_fire_load_incoming_0_will_fire ? _GEN_73 : will_fire_load_retry_0_will_fire & _GEN_127;
  wire        _GEN_129 = ldq_retry_idx == 5'h18;
  wire        _GEN_130 = will_fire_load_wakeup_0_will_fire ? _GEN_43 : will_fire_load_incoming_0_will_fire ? _GEN_74 : will_fire_load_retry_0_will_fire & _GEN_129;
  wire        _GEN_131 = ldq_retry_idx == 5'h19;
  wire        _GEN_132 = will_fire_load_wakeup_0_will_fire ? _GEN_44 : will_fire_load_incoming_0_will_fire ? _GEN_75 : will_fire_load_retry_0_will_fire & _GEN_131;
  wire        _GEN_133 = ldq_retry_idx == 5'h1A;
  wire        _GEN_134 = will_fire_load_wakeup_0_will_fire ? _GEN_45 : will_fire_load_incoming_0_will_fire ? _GEN_76 : will_fire_load_retry_0_will_fire & _GEN_133;
  wire        _GEN_135 = ldq_retry_idx == 5'h1B;
  wire        _GEN_136 = will_fire_load_wakeup_0_will_fire ? _GEN_46 : will_fire_load_incoming_0_will_fire ? _GEN_77 : will_fire_load_retry_0_will_fire & _GEN_135;
  wire        _GEN_137 = ldq_retry_idx == 5'h1C;
  wire        _GEN_138 = will_fire_load_wakeup_0_will_fire ? _GEN_47 : will_fire_load_incoming_0_will_fire ? _GEN_78 : will_fire_load_retry_0_will_fire & _GEN_137;
  wire        _GEN_139 = ldq_retry_idx == 5'h1D;
  wire        _GEN_140 = will_fire_load_wakeup_0_will_fire ? _GEN_48 : will_fire_load_incoming_0_will_fire ? _GEN_79 : will_fire_load_retry_0_will_fire & _GEN_139;
  wire        _GEN_141 = ldq_retry_idx == 5'h1E;
  wire        _GEN_142 = will_fire_load_wakeup_0_will_fire ? _GEN_49 : will_fire_load_incoming_0_will_fire ? _GEN_80 : will_fire_load_retry_0_will_fire & _GEN_141;
  wire        _GEN_143 = will_fire_load_wakeup_0_will_fire ? (&ldq_wakeup_idx) : will_fire_load_incoming_0_will_fire ? (&_mem_incoming_uop_WIRE_0_ldq_idx) : will_fire_load_retry_0_will_fire & (&ldq_retry_idx);
  wire        will_fire_stad_incoming_1_will_fire = _can_fire_sta_incoming_T_3 & exe_req_1_bits_uop_ctrl_is_std & ~will_fire_load_incoming_1_will_fire & ~will_fire_load_incoming_1_will_fire;
  wire        _will_fire_sta_incoming_1_will_fire_T_2 = ~will_fire_load_incoming_1_will_fire & ~will_fire_stad_incoming_1_will_fire;
  wire        _will_fire_sta_incoming_1_will_fire_T_6 = ~will_fire_load_incoming_1_will_fire & ~will_fire_stad_incoming_1_will_fire;
  wire        will_fire_sta_incoming_1_will_fire = _can_fire_sta_incoming_T_3 & ~exe_req_1_bits_uop_ctrl_is_std & _will_fire_sta_incoming_1_will_fire_T_2 & _will_fire_sta_incoming_1_will_fire_T_6 & ~will_fire_stad_incoming_1_will_fire;
  wire        _will_fire_sfence_1_will_fire_T_2 = _will_fire_sta_incoming_1_will_fire_T_2 & ~will_fire_sta_incoming_1_will_fire;
  wire        _will_fire_release_1_will_fire_T_6 = _will_fire_sta_incoming_1_will_fire_T_6 & ~will_fire_sta_incoming_1_will_fire;
  wire        _will_fire_std_incoming_1_will_fire_T_14 = ~will_fire_stad_incoming_1_will_fire & ~will_fire_sta_incoming_1_will_fire;
  wire        will_fire_std_incoming_1_will_fire = exe_req_1_valid & exe_req_1_bits_uop_ctrl_is_std & ~exe_req_1_bits_uop_ctrl_is_sta & _will_fire_std_incoming_1_will_fire_T_14;
  wire        _will_fire_sfence_1_will_fire_T_14 = _will_fire_std_incoming_1_will_fire_T_14 & ~will_fire_std_incoming_1_will_fire;
  wire        will_fire_sfence_1_will_fire = exe_req_1_valid & exe_req_1_bits_sfence_valid & _will_fire_sfence_1_will_fire_T_2 & _will_fire_sfence_1_will_fire_T_14;
  wire        _will_fire_hella_incoming_1_will_fire_T_2 = _will_fire_sfence_1_will_fire_T_2 & ~will_fire_sfence_1_will_fire;
  assign will_fire_release_1_will_fire = io_dmem_release_valid & _will_fire_release_1_will_fire_T_6;
  wire        _will_fire_load_retry_1_will_fire_T_6 = _will_fire_release_1_will_fire_T_6 & ~will_fire_release_1_will_fire;
  wire        will_fire_hella_incoming_1_will_fire = _GEN_0 & _GEN_2 & _will_fire_hella_incoming_1_will_fire_T_2 & ~will_fire_load_incoming_1_will_fire;
  wire        _will_fire_load_retry_1_will_fire_T_2 = _will_fire_hella_incoming_1_will_fire_T_2 & ~will_fire_hella_incoming_1_will_fire;
  wire        _will_fire_hella_wakeup_1_will_fire_T_10 = ~will_fire_load_incoming_1_will_fire & ~will_fire_hella_incoming_1_will_fire;
  wire        will_fire_hella_wakeup_1_will_fire = _GEN & _GEN_1 & _will_fire_hella_wakeup_1_will_fire_T_10;
  wire        _will_fire_load_retry_1_will_fire_T_10 = _will_fire_hella_wakeup_1_will_fire_T_10 & ~will_fire_hella_wakeup_1_will_fire;
  wire        will_fire_load_retry_1_will_fire = casez_tmp_123 & casez_tmp_201 & casez_tmp_203 & ~casez_tmp_207 & ~casez_tmp_208 & can_fire_load_retry_REG_1 & ~store_needs_order & ~casez_tmp_205 & _will_fire_load_retry_1_will_fire_T_2 & _will_fire_load_retry_1_will_fire_T_6 & _will_fire_load_retry_1_will_fire_T_10;
  wire        _will_fire_sta_retry_1_will_fire_T_2 = _will_fire_load_retry_1_will_fire_T_2 & ~will_fire_load_retry_1_will_fire;
  wire        _will_fire_sta_retry_1_will_fire_T_6 = _will_fire_load_retry_1_will_fire_T_6 & ~will_fire_load_retry_1_will_fire;
  wire        will_fire_sta_retry_1_will_fire = casez_tmp_209 & casez_tmp_289 & casez_tmp_291 & can_fire_sta_retry_REG_1 & ~(can_fire_std_incoming_0 & _mem_incoming_uop_WIRE_0_stq_idx == stq_retry_idx) & _will_fire_sta_retry_1_will_fire_T_2 & _will_fire_sta_retry_1_will_fire_T_6 & _will_fire_sfence_1_will_fire_T_14 & ~will_fire_sfence_1_will_fire;
  assign _will_fire_store_commit_1_T_2 = _will_fire_sta_retry_1_will_fire_T_2 & ~will_fire_sta_retry_1_will_fire;
  wire        will_fire_load_wakeup_1_will_fire = casez_tmp_293 & casez_tmp_371 & ~casez_tmp_376 & ~casez_tmp_373 & ~casez_tmp_375 & ~casez_tmp_377 & ~casez_tmp_379 & ~casez_tmp_380 & ~store_needs_order & (~casez_tmp_374 | io_core_commit_load_at_rob_head & ldq_head == ldq_wakeup_idx & casez_tmp_378 == 32'h0) & _will_fire_sta_retry_1_will_fire_T_6 & ~will_fire_sta_retry_1_will_fire & _will_fire_load_retry_1_will_fire_T_10 & ~will_fire_load_retry_1_will_fire;
  wire        _exe_cmd_T_7 = will_fire_load_incoming_1_will_fire | will_fire_stad_incoming_1_will_fire;
  wire        _GEN_144 = _exe_cmd_T_7 | will_fire_sta_incoming_1_will_fire;
  wire        _GEN_145 = _GEN_19 | _GEN_82;
  wire        _GEN_146 = _GEN_20 | _GEN_84;
  wire        _GEN_147 = _GEN_21 | _GEN_86;
  wire        _GEN_148 = _GEN_22 | _GEN_88;
  wire        _GEN_149 = _GEN_23 | _GEN_90;
  wire        _GEN_150 = _GEN_24 | _GEN_92;
  wire        _GEN_151 = _GEN_25 | _GEN_94;
  wire        _GEN_152 = _GEN_26 | _GEN_96;
  wire        _GEN_153 = _GEN_27 | _GEN_98;
  wire        _GEN_154 = _GEN_28 | _GEN_100;
  wire        _GEN_155 = _GEN_29 | _GEN_102;
  wire        _GEN_156 = _GEN_30 | _GEN_104;
  wire        _GEN_157 = _GEN_31 | _GEN_106;
  wire        _GEN_158 = _GEN_32 | _GEN_108;
  wire        _GEN_159 = _GEN_33 | _GEN_110;
  wire        _GEN_160 = _GEN_34 | _GEN_112;
  wire        _GEN_161 = _GEN_35 | _GEN_114;
  wire        _GEN_162 = _GEN_36 | _GEN_116;
  wire        _GEN_163 = _GEN_37 | _GEN_118;
  wire        _GEN_164 = _GEN_38 | _GEN_120;
  wire        _GEN_165 = _GEN_39 | _GEN_122;
  wire        _GEN_166 = _GEN_40 | _GEN_124;
  wire        _GEN_167 = _GEN_41 | _GEN_126;
  wire        _GEN_168 = _GEN_42 | _GEN_128;
  wire        _GEN_169 = _GEN_43 | _GEN_130;
  wire        _GEN_170 = _GEN_44 | _GEN_132;
  wire        _GEN_171 = _GEN_45 | _GEN_134;
  wire        _GEN_172 = _GEN_46 | _GEN_136;
  wire        _GEN_173 = _GEN_47 | _GEN_138;
  wire        _GEN_174 = _GEN_48 | _GEN_140;
  wire        _GEN_175 = _GEN_49 | _GEN_142;
  wire        _GEN_176 = (&ldq_wakeup_idx) | _GEN_143;
  wire        _GEN_177 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h0;
  wire        _GEN_178 = _GEN_177 | _GEN_82;
  wire        _GEN_179 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h1;
  wire        _GEN_180 = _GEN_179 | _GEN_84;
  wire        _GEN_181 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h2;
  wire        _GEN_182 = _GEN_181 | _GEN_86;
  wire        _GEN_183 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h3;
  wire        _GEN_184 = _GEN_183 | _GEN_88;
  wire        _GEN_185 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h4;
  wire        _GEN_186 = _GEN_185 | _GEN_90;
  wire        _GEN_187 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h5;
  wire        _GEN_188 = _GEN_187 | _GEN_92;
  wire        _GEN_189 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h6;
  wire        _GEN_190 = _GEN_189 | _GEN_94;
  wire        _GEN_191 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h7;
  wire        _GEN_192 = _GEN_191 | _GEN_96;
  wire        _GEN_193 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h8;
  wire        _GEN_194 = _GEN_193 | _GEN_98;
  wire        _GEN_195 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h9;
  wire        _GEN_196 = _GEN_195 | _GEN_100;
  wire        _GEN_197 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'hA;
  wire        _GEN_198 = _GEN_197 | _GEN_102;
  wire        _GEN_199 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'hB;
  wire        _GEN_200 = _GEN_199 | _GEN_104;
  wire        _GEN_201 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'hC;
  wire        _GEN_202 = _GEN_201 | _GEN_106;
  wire        _GEN_203 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'hD;
  wire        _GEN_204 = _GEN_203 | _GEN_108;
  wire        _GEN_205 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'hE;
  wire        _GEN_206 = _GEN_205 | _GEN_110;
  wire        _GEN_207 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'hF;
  wire        _GEN_208 = _GEN_207 | _GEN_112;
  wire        _GEN_209 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h10;
  wire        _GEN_210 = _GEN_209 | _GEN_114;
  wire        _GEN_211 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h11;
  wire        _GEN_212 = _GEN_211 | _GEN_116;
  wire        _GEN_213 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h12;
  wire        _GEN_214 = _GEN_213 | _GEN_118;
  wire        _GEN_215 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h13;
  wire        _GEN_216 = _GEN_215 | _GEN_120;
  wire        _GEN_217 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h14;
  wire        _GEN_218 = _GEN_217 | _GEN_122;
  wire        _GEN_219 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h15;
  wire        _GEN_220 = _GEN_219 | _GEN_124;
  wire        _GEN_221 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h16;
  wire        _GEN_222 = _GEN_221 | _GEN_126;
  wire        _GEN_223 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h17;
  wire        _GEN_224 = _GEN_223 | _GEN_128;
  wire        _GEN_225 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h18;
  wire        _GEN_226 = _GEN_225 | _GEN_130;
  wire        _GEN_227 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h19;
  wire        _GEN_228 = _GEN_227 | _GEN_132;
  wire        _GEN_229 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h1A;
  wire        _GEN_230 = _GEN_229 | _GEN_134;
  wire        _GEN_231 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h1B;
  wire        _GEN_232 = _GEN_231 | _GEN_136;
  wire        _GEN_233 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h1C;
  wire        _GEN_234 = _GEN_233 | _GEN_138;
  wire        _GEN_235 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h1D;
  wire        _GEN_236 = _GEN_235 | _GEN_140;
  wire        _GEN_237 = _mem_incoming_uop_WIRE_1_ldq_idx == 5'h1E;
  wire        _GEN_238 = _GEN_237 | _GEN_142;
  wire        _GEN_239 = (&_mem_incoming_uop_WIRE_1_ldq_idx) | _GEN_143;
  wire        _GEN_240 = will_fire_load_retry_1_will_fire & _GEN_81 | _GEN_82;
  wire        _GEN_241 = will_fire_load_retry_1_will_fire & _GEN_83 | _GEN_84;
  wire        _GEN_242 = will_fire_load_retry_1_will_fire & _GEN_85 | _GEN_86;
  wire        _GEN_243 = will_fire_load_retry_1_will_fire & _GEN_87 | _GEN_88;
  wire        _GEN_244 = will_fire_load_retry_1_will_fire & _GEN_89 | _GEN_90;
  wire        _GEN_245 = will_fire_load_retry_1_will_fire & _GEN_91 | _GEN_92;
  wire        _GEN_246 = will_fire_load_retry_1_will_fire & _GEN_93 | _GEN_94;
  wire        _GEN_247 = will_fire_load_retry_1_will_fire & _GEN_95 | _GEN_96;
  wire        _GEN_248 = will_fire_load_retry_1_will_fire & _GEN_97 | _GEN_98;
  wire        _GEN_249 = will_fire_load_retry_1_will_fire & _GEN_99 | _GEN_100;
  wire        _GEN_250 = will_fire_load_retry_1_will_fire & _GEN_101 | _GEN_102;
  wire        _GEN_251 = will_fire_load_retry_1_will_fire & _GEN_103 | _GEN_104;
  wire        _GEN_252 = will_fire_load_retry_1_will_fire & _GEN_105 | _GEN_106;
  wire        _GEN_253 = will_fire_load_retry_1_will_fire & _GEN_107 | _GEN_108;
  wire        _GEN_254 = will_fire_load_retry_1_will_fire & _GEN_109 | _GEN_110;
  wire        _GEN_255 = will_fire_load_retry_1_will_fire & _GEN_111 | _GEN_112;
  wire        _GEN_256 = will_fire_load_retry_1_will_fire & _GEN_113 | _GEN_114;
  wire        _GEN_257 = will_fire_load_retry_1_will_fire & _GEN_115 | _GEN_116;
  wire        _GEN_258 = will_fire_load_retry_1_will_fire & _GEN_117 | _GEN_118;
  wire        _GEN_259 = will_fire_load_retry_1_will_fire & _GEN_119 | _GEN_120;
  wire        _GEN_260 = will_fire_load_retry_1_will_fire & _GEN_121 | _GEN_122;
  wire        _GEN_261 = will_fire_load_retry_1_will_fire & _GEN_123 | _GEN_124;
  wire        _GEN_262 = will_fire_load_retry_1_will_fire & _GEN_125 | _GEN_126;
  wire        _GEN_263 = will_fire_load_retry_1_will_fire & _GEN_127 | _GEN_128;
  wire        _GEN_264 = will_fire_load_retry_1_will_fire & _GEN_129 | _GEN_130;
  wire        _GEN_265 = will_fire_load_retry_1_will_fire & _GEN_131 | _GEN_132;
  wire        _GEN_266 = will_fire_load_retry_1_will_fire & _GEN_133 | _GEN_134;
  wire        _GEN_267 = will_fire_load_retry_1_will_fire & _GEN_135 | _GEN_136;
  wire        _GEN_268 = will_fire_load_retry_1_will_fire & _GEN_137 | _GEN_138;
  wire        _GEN_269 = will_fire_load_retry_1_will_fire & _GEN_139 | _GEN_140;
  wire        _GEN_270 = will_fire_load_retry_1_will_fire & _GEN_141 | _GEN_142;
  wire        _GEN_271 = will_fire_load_retry_1_will_fire & (&ldq_retry_idx) | _GEN_143;
  wire        _exe_tlb_uop_T_2 = _exe_cmd_T | will_fire_sta_incoming_0_will_fire | will_fire_sfence_0_will_fire;
  wire [6:0]  _exe_tlb_uop_T_4_pdst = will_fire_sta_retry_0_will_fire ? casez_tmp_246 : 7'h0;
  wire        exe_tlb_uop_0_ctrl_is_load = _exe_tlb_uop_T_2 ? exe_req_0_bits_uop_ctrl_is_load : will_fire_load_retry_0_will_fire ? casez_tmp_138 : will_fire_sta_retry_0_will_fire & casez_tmp_224;
  wire        exe_tlb_uop_0_ctrl_is_sta = _exe_tlb_uop_T_2 ? exe_req_0_bits_uop_ctrl_is_sta : will_fire_load_retry_0_will_fire ? casez_tmp_139 : will_fire_sta_retry_0_will_fire & casez_tmp_225;
  wire [19:0] exe_tlb_uop_0_br_mask = _exe_tlb_uop_T_2 ? exe_req_0_bits_uop_br_mask : will_fire_load_retry_0_will_fire ? casez_tmp_148 : will_fire_sta_retry_0_will_fire ? casez_tmp_234 : 20'h0;
  wire [6:0]  _mem_xcpt_uops_WIRE_0_rob_idx = _exe_tlb_uop_T_2 ? _mem_incoming_uop_WIRE_0_rob_idx : will_fire_load_retry_0_will_fire ? casez_tmp_156 : will_fire_sta_retry_0_will_fire ? casez_tmp_242 : 7'h0;
  wire [4:0]  _mem_xcpt_uops_WIRE_0_ldq_idx = _exe_tlb_uop_T_2 ? _mem_incoming_uop_WIRE_0_ldq_idx : will_fire_load_retry_0_will_fire ? casez_tmp_157 : will_fire_sta_retry_0_will_fire ? casez_tmp_243 : 5'h0;
  wire [4:0]  _mem_xcpt_uops_WIRE_0_stq_idx = _exe_tlb_uop_T_2 ? _mem_incoming_uop_WIRE_0_stq_idx : will_fire_load_retry_0_will_fire ? casez_tmp_158 : will_fire_sta_retry_0_will_fire ? casez_tmp_244 : 5'h0;
  wire [4:0]  exe_tlb_uop_0_mem_cmd = _exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_mem_cmd : io_core_exe_0_req_bits_uop_mem_cmd) : will_fire_load_retry_0_will_fire ? casez_tmp_171 : will_fire_sta_retry_0_will_fire ? casez_tmp_259 : 5'h0;
  wire [1:0]  exe_tlb_uop_0_mem_size = _exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_mem_size : io_core_exe_0_req_bits_uop_mem_size) : will_fire_load_retry_0_will_fire ? casez_tmp_172 : will_fire_sta_retry_0_will_fire ? casez_tmp_260 : 2'h0;
  wire        exe_tlb_uop_0_is_fence = _exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_fence : io_core_exe_0_req_bits_uop_is_fence) : will_fire_load_retry_0_will_fire ? casez_tmp_174 : will_fire_sta_retry_0_will_fire & casez_tmp_262;
  wire        _mem_xcpt_uops_WIRE_0_uses_ldq = _exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_uses_ldq : io_core_exe_0_req_bits_uop_uses_ldq) : will_fire_load_retry_0_will_fire ? casez_tmp_177 : will_fire_sta_retry_0_will_fire & casez_tmp_265;
  wire        _mem_xcpt_uops_WIRE_0_uses_stq = _exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_uses_stq : io_core_exe_0_req_bits_uop_uses_stq) : will_fire_load_retry_0_will_fire ? casez_tmp_178 : will_fire_sta_retry_0_will_fire & casez_tmp_266;
  wire        _exe_tlb_uop_T_9 = _exe_cmd_T_7 | will_fire_sta_incoming_1_will_fire | will_fire_sfence_1_will_fire;
  wire [6:0]  _exe_tlb_uop_T_11_pdst = will_fire_sta_retry_1_will_fire ? casez_tmp_246 : 7'h0;
  wire        exe_tlb_uop_1_ctrl_is_load = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_ctrl_is_load : will_fire_load_retry_1_will_fire ? casez_tmp_138 : will_fire_sta_retry_1_will_fire & casez_tmp_224;
  wire        exe_tlb_uop_1_ctrl_is_sta = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_ctrl_is_sta : will_fire_load_retry_1_will_fire ? casez_tmp_139 : will_fire_sta_retry_1_will_fire & casez_tmp_225;
  wire [19:0] exe_tlb_uop_1_br_mask = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_br_mask : will_fire_load_retry_1_will_fire ? casez_tmp_148 : will_fire_sta_retry_1_will_fire ? casez_tmp_234 : 20'h0;
  wire [6:0]  _mem_xcpt_uops_WIRE_1_rob_idx = _exe_tlb_uop_T_9 ? _mem_incoming_uop_WIRE_1_rob_idx : will_fire_load_retry_1_will_fire ? casez_tmp_156 : will_fire_sta_retry_1_will_fire ? casez_tmp_242 : 7'h0;
  wire [4:0]  _mem_xcpt_uops_WIRE_1_ldq_idx = _exe_tlb_uop_T_9 ? _mem_incoming_uop_WIRE_1_ldq_idx : will_fire_load_retry_1_will_fire ? casez_tmp_157 : will_fire_sta_retry_1_will_fire ? casez_tmp_243 : 5'h0;
  wire [4:0]  _mem_xcpt_uops_WIRE_1_stq_idx = _exe_tlb_uop_T_9 ? _mem_incoming_uop_WIRE_1_stq_idx : will_fire_load_retry_1_will_fire ? casez_tmp_158 : will_fire_sta_retry_1_will_fire ? casez_tmp_244 : 5'h0;
  wire [4:0]  exe_tlb_uop_1_mem_cmd = _exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_mem_cmd : io_core_exe_0_req_bits_uop_mem_cmd) : will_fire_load_retry_1_will_fire ? casez_tmp_171 : will_fire_sta_retry_1_will_fire ? casez_tmp_259 : 5'h0;
  wire [1:0]  exe_tlb_uop_1_mem_size = _exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_mem_size : io_core_exe_0_req_bits_uop_mem_size) : will_fire_load_retry_1_will_fire ? casez_tmp_172 : will_fire_sta_retry_1_will_fire ? casez_tmp_260 : 2'h0;
  wire        exe_tlb_uop_1_is_fence = _exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_fence : io_core_exe_0_req_bits_uop_is_fence) : will_fire_load_retry_1_will_fire ? casez_tmp_174 : will_fire_sta_retry_1_will_fire & casez_tmp_262;
  wire        _mem_xcpt_uops_WIRE_1_uses_ldq = _exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_uses_ldq : io_core_exe_0_req_bits_uop_uses_ldq) : will_fire_load_retry_1_will_fire ? casez_tmp_177 : will_fire_sta_retry_1_will_fire & casez_tmp_265;
  wire        _mem_xcpt_uops_WIRE_1_uses_stq = _exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_uses_stq : io_core_exe_0_req_bits_uop_uses_stq) : will_fire_load_retry_1_will_fire ? casez_tmp_178 : will_fire_sta_retry_1_will_fire & casez_tmp_266;
  wire        _exe_tlb_vaddr_T_1 = _exe_cmd_T | will_fire_sta_incoming_0_will_fire;
  wire [39:0] _exe_tlb_vaddr_T_2 = will_fire_hella_incoming_0_will_fire ? hella_req_addr : 40'h0;
  wire [39:0] _exe_tlb_vaddr_T_3 = will_fire_sta_retry_0_will_fire ? casez_tmp_290 : _exe_tlb_vaddr_T_2;
  wire [39:0] _GEN_272 = {1'h0, exe_req_0_bits_sfence_bits_addr};
  wire [39:0] exe_tlb_vaddr_0 = _exe_tlb_vaddr_T_1 ? exe_req_0_bits_addr : will_fire_sfence_0_will_fire ? _GEN_272 : will_fire_load_retry_0_will_fire ? casez_tmp_202 : _exe_tlb_vaddr_T_3;
  wire        _exe_tlb_vaddr_T_8 = _exe_cmd_T_7 | will_fire_sta_incoming_1_will_fire;
  wire [39:0] _exe_tlb_vaddr_T_9 = will_fire_hella_incoming_1_will_fire ? hella_req_addr : 40'h0;
  wire [39:0] _exe_tlb_vaddr_T_10 = will_fire_sta_retry_1_will_fire ? casez_tmp_290 : _exe_tlb_vaddr_T_9;
  wire [39:0] _GEN_273 = {1'h0, exe_req_1_bits_sfence_bits_addr};
  wire [39:0] exe_tlb_vaddr_1 = _exe_tlb_vaddr_T_8 ? exe_req_1_bits_addr : will_fire_sfence_1_will_fire ? _GEN_273 : will_fire_load_retry_1_will_fire ? casez_tmp_202 : _exe_tlb_vaddr_T_10;
  wire        _stq_idx_T = will_fire_sta_incoming_0_will_fire | will_fire_stad_incoming_0_will_fire;
  wire        _stq_idx_T_1 = will_fire_sta_incoming_1_will_fire | will_fire_stad_incoming_1_will_fire;
  reg         mem_xcpt_valids_0;
  reg         mem_xcpt_valids_1;
  reg  [19:0] mem_xcpt_uops_0_br_mask;
  reg  [6:0]  mem_xcpt_uops_0_rob_idx;
  reg  [4:0]  mem_xcpt_uops_0_ldq_idx;
  reg  [4:0]  mem_xcpt_uops_0_stq_idx;
  reg         mem_xcpt_uops_0_uses_ldq;
  reg         mem_xcpt_uops_0_uses_stq;
  reg  [19:0] mem_xcpt_uops_1_br_mask;
  reg  [6:0]  mem_xcpt_uops_1_rob_idx;
  reg  [4:0]  mem_xcpt_uops_1_ldq_idx;
  reg  [4:0]  mem_xcpt_uops_1_stq_idx;
  reg         mem_xcpt_uops_1_uses_ldq;
  reg         mem_xcpt_uops_1_uses_stq;
  reg  [3:0]  mem_xcpt_causes_0;
  reg  [3:0]  mem_xcpt_causes_1;
  reg  [39:0] mem_xcpt_vaddrs_0;
  reg  [39:0] mem_xcpt_vaddrs_1;
  assign mem_xcpt_valid = mem_xcpt_valids_0 | mem_xcpt_valids_1;
  wire        exe_tlb_miss_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_miss;
  wire        exe_tlb_miss_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_miss;
  wire [32:0] exe_tlb_paddr_0 = {_dtlb_io_resp_0_paddr[32:12], exe_tlb_vaddr_0[11:0]};
  wire [32:0] exe_tlb_paddr_1 = {_dtlb_io_resp_1_paddr[32:12], exe_tlb_vaddr_1[11:0]};
  reg         REG;
  reg         REG_1;
  wire        _io_dmem_req_valid_output = dmem_req_0_valid | dmem_req_1_valid;
  wire        _dmem_req_fire_T_2 = io_dmem_req_ready & _io_dmem_req_valid_output;
  wire        dmem_req_fire_1 = dmem_req_1_valid & _dmem_req_fire_T_2;
  wire [39:0] _GEN_274 = {7'h0, _dtlb_io_resp_0_paddr[32:12], exe_tlb_vaddr_0[11:0]};
  wire        _GEN_275 = will_fire_load_incoming_0_will_fire | will_fire_load_retry_0_will_fire;
  assign _GEN_2 = hella_state == 3'h1;
  wire        _GEN_276 = will_fire_store_commit_0_will_fire | will_fire_load_wakeup_0_will_fire;
  assign _GEN_1 = hella_state == 3'h5;
  assign dmem_req_0_valid = will_fire_load_incoming_0_will_fire ? ~exe_tlb_miss_0 & _dtlb_io_resp_0_cacheable : will_fire_load_retry_0_will_fire ? ~exe_tlb_miss_0 & _dtlb_io_resp_0_cacheable : _GEN_276 | (will_fire_hella_incoming_0_will_fire ? ~io_hellacache_s1_kill : will_fire_hella_wakeup_0_will_fire);
  wire [39:0] _GEN_277 = {7'h0, hella_paddr};
  wire [39:0] _mem_paddr_WIRE_0 = will_fire_load_incoming_0_will_fire | will_fire_load_retry_0_will_fire ? _GEN_274 : will_fire_store_commit_0_will_fire ? casez_tmp_80 : will_fire_load_wakeup_0_will_fire ? casez_tmp_372 : will_fire_hella_incoming_0_will_fire ? _GEN_274 : will_fire_hella_wakeup_0_will_fire ? _GEN_277 : 40'h0;
  wire        _GEN_278 = _stq_idx_T | will_fire_sta_retry_0_will_fire;
  wire        _io_core_fp_stdata_ready_output = ~will_fire_std_incoming_0_will_fire & ~will_fire_stad_incoming_0_will_fire;
  wire        fp_stdata_fire = _io_core_fp_stdata_ready_output & io_core_fp_stdata_valid;
  wire        _stq_bits_data_bits_T = will_fire_std_incoming_0_will_fire | will_fire_stad_incoming_0_will_fire;
  wire        _GEN_279 = _stq_bits_data_bits_T | fp_stdata_fire;
  wire [4:0]  sidx = _stq_bits_data_bits_T ? _mem_incoming_uop_WIRE_0_stq_idx : io_core_fp_stdata_bits_uop_stq_idx;
  reg         casez_tmp_381;
  always @(*) begin
    casez (sidx)
      5'b00000:
        casez_tmp_381 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_381 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_381 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_381 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_381 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_381 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_381 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_381 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_381 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_381 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_381 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_381 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_381 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_381 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_381 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_381 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_381 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_381 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_381 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_381 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_381 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_381 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_381 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_381 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_381 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_381 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_381 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_381 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_381 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_381 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_381 = stq_30_bits_data_valid;
      default:
        casez_tmp_381 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  wire [39:0] _GEN_280 = {7'h0, _dtlb_io_resp_1_paddr[32:12], exe_tlb_vaddr_1[11:0]};
  wire        _GEN_281 = will_fire_load_incoming_1_will_fire | will_fire_load_retry_1_will_fire;
  wire        _GEN_282 = will_fire_store_commit_1_will_fire | will_fire_load_wakeup_1_will_fire;
  assign dmem_req_1_valid = will_fire_load_incoming_1_will_fire ? ~exe_tlb_miss_1 & _dtlb_io_resp_1_cacheable : will_fire_load_retry_1_will_fire ? ~exe_tlb_miss_1 & _dtlb_io_resp_1_cacheable : _GEN_282 | (will_fire_hella_incoming_1_will_fire ? ~io_hellacache_s1_kill : will_fire_hella_wakeup_1_will_fire);
  wire [39:0] _mem_paddr_WIRE_1 = will_fire_load_incoming_1_will_fire | will_fire_load_retry_1_will_fire ? _GEN_280 : will_fire_store_commit_1_will_fire ? casez_tmp_80 : will_fire_load_wakeup_1_will_fire ? casez_tmp_372 : will_fire_hella_incoming_1_will_fire ? _GEN_280 : will_fire_hella_wakeup_1_will_fire ? _GEN_277 : 40'h0;
  wire        _GEN_283 = _stq_idx_T_1 | will_fire_sta_retry_1_will_fire;
  wire        _stq_bits_data_bits_T_2 = will_fire_std_incoming_1_will_fire | will_fire_stad_incoming_1_will_fire;
  wire [4:0]  sidx_1 = _stq_bits_data_bits_T_2 ? _mem_incoming_uop_WIRE_1_stq_idx : io_core_fp_stdata_bits_uop_stq_idx;
  reg         casez_tmp_382;
  always @(*) begin
    casez (sidx_1)
      5'b00000:
        casez_tmp_382 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_382 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_382 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_382 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_382 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_382 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_382 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_382 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_382 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_382 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_382 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_382 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_382 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_382 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_382 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_382 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_382 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_382 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_382 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_382 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_382 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_382 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_382 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_382 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_382 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_382 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_382 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_382 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_382 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_382 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_382 = stq_30_bits_data_valid;
      default:
        casez_tmp_382 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg         fired_load_incoming_REG;
  reg         fired_load_incoming_REG_1;
  reg         fired_stad_incoming_REG;
  reg         fired_stad_incoming_REG_1;
  reg         fired_sta_incoming_REG;
  reg         fired_sta_incoming_REG_1;
  reg         fired_std_incoming_REG;
  reg         fired_std_incoming_REG_1;
  reg         fired_stdf_incoming;
  reg         fired_sfence_0;
  reg         fired_sfence_1;
  reg         fired_release_0;
  reg         fired_release_1;
  reg         fired_load_retry_REG;
  reg         fired_load_retry_REG_1;
  reg         fired_sta_retry_REG;
  reg         fired_sta_retry_REG_1;
  reg         fired_load_wakeup_REG;
  reg         fired_load_wakeup_REG_1;
  reg  [19:0] mem_incoming_uop_0_br_mask;
  reg  [6:0]  mem_incoming_uop_0_rob_idx;
  reg  [4:0]  mem_incoming_uop_0_ldq_idx;
  reg  [4:0]  mem_incoming_uop_0_stq_idx;
  reg  [6:0]  mem_incoming_uop_0_pdst;
  reg         mem_incoming_uop_0_fp_val;
  reg  [19:0] mem_incoming_uop_1_br_mask;
  reg  [6:0]  mem_incoming_uop_1_rob_idx;
  reg  [4:0]  mem_incoming_uop_1_ldq_idx;
  reg  [4:0]  mem_incoming_uop_1_stq_idx;
  reg  [6:0]  mem_incoming_uop_1_pdst;
  reg         mem_incoming_uop_1_fp_val;
  reg  [19:0] mem_ldq_incoming_e_0_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_incoming_e_0_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_incoming_e_0_bits_uop_mem_size;
  reg  [31:0] mem_ldq_incoming_e_0_bits_st_dep_mask;
  reg  [19:0] mem_ldq_incoming_e_1_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_incoming_e_1_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_incoming_e_1_bits_uop_mem_size;
  reg  [31:0] mem_ldq_incoming_e_1_bits_st_dep_mask;
  reg         mem_stq_incoming_e_0_valid;
  reg  [19:0] mem_stq_incoming_e_0_bits_uop_br_mask;
  reg  [6:0]  mem_stq_incoming_e_0_bits_uop_rob_idx;
  reg  [4:0]  mem_stq_incoming_e_0_bits_uop_stq_idx;
  reg  [1:0]  mem_stq_incoming_e_0_bits_uop_mem_size;
  reg         mem_stq_incoming_e_0_bits_uop_is_amo;
  reg         mem_stq_incoming_e_0_bits_addr_valid;
  reg         mem_stq_incoming_e_0_bits_addr_is_virtual;
  reg         mem_stq_incoming_e_0_bits_data_valid;
  reg         mem_stq_incoming_e_1_valid;
  reg  [19:0] mem_stq_incoming_e_1_bits_uop_br_mask;
  reg  [6:0]  mem_stq_incoming_e_1_bits_uop_rob_idx;
  reg  [4:0]  mem_stq_incoming_e_1_bits_uop_stq_idx;
  reg  [1:0]  mem_stq_incoming_e_1_bits_uop_mem_size;
  reg         mem_stq_incoming_e_1_bits_uop_is_amo;
  reg         mem_stq_incoming_e_1_bits_addr_valid;
  reg         mem_stq_incoming_e_1_bits_addr_is_virtual;
  reg         mem_stq_incoming_e_1_bits_data_valid;
  reg  [19:0] mem_ldq_wakeup_e_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_wakeup_e_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_wakeup_e_bits_uop_mem_size;
  reg  [31:0] mem_ldq_wakeup_e_bits_st_dep_mask;
  reg  [19:0] mem_ldq_retry_e_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_retry_e_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_retry_e_bits_uop_mem_size;
  reg  [31:0] mem_ldq_retry_e_bits_st_dep_mask;
  reg         mem_stq_retry_e_valid;
  reg  [19:0] mem_stq_retry_e_bits_uop_br_mask;
  reg  [6:0]  mem_stq_retry_e_bits_uop_rob_idx;
  reg  [4:0]  mem_stq_retry_e_bits_uop_stq_idx;
  reg  [1:0]  mem_stq_retry_e_bits_uop_mem_size;
  reg         mem_stq_retry_e_bits_uop_is_amo;
  reg         mem_stq_retry_e_bits_data_valid;
  wire [31:0] lcam_st_dep_mask_0 = fired_load_incoming_REG ? mem_ldq_incoming_e_0_bits_st_dep_mask : fired_load_retry_REG ? mem_ldq_retry_e_bits_st_dep_mask : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_st_dep_mask : 32'h0;
  wire [31:0] lcam_st_dep_mask_1 = fired_load_incoming_REG_1 ? mem_ldq_incoming_e_1_bits_st_dep_mask : fired_load_retry_REG_1 ? mem_ldq_retry_e_bits_st_dep_mask : fired_load_wakeup_REG_1 ? mem_ldq_wakeup_e_bits_st_dep_mask : 32'h0;
  wire        _lcam_stq_idx_T = fired_stad_incoming_REG | fired_sta_incoming_REG;
  wire        _lcam_stq_idx_T_3 = fired_stad_incoming_REG_1 | fired_sta_incoming_REG_1;
  reg  [19:0] mem_stdf_uop_br_mask;
  reg  [6:0]  mem_stdf_uop_rob_idx;
  reg  [4:0]  mem_stdf_uop_stq_idx;
  reg         mem_tlb_miss_0;
  reg         mem_tlb_miss_1;
  reg         mem_tlb_uncacheable_0;
  reg         mem_tlb_uncacheable_1;
  reg  [39:0] mem_paddr_0;
  reg  [39:0] mem_paddr_1;
  reg         clr_bsy_valid_0;
  reg         clr_bsy_valid_1;
  reg  [6:0]  clr_bsy_rob_idx_0;
  reg  [6:0]  clr_bsy_rob_idx_1;
  reg  [19:0] clr_bsy_brmask_0;
  reg  [19:0] clr_bsy_brmask_1;
  reg         io_core_clr_bsy_0_valid_REG;
  reg         io_core_clr_bsy_0_valid_REG_1;
  reg         io_core_clr_bsy_0_valid_REG_2;
  reg         io_core_clr_bsy_1_valid_REG;
  reg         io_core_clr_bsy_1_valid_REG_1;
  reg         io_core_clr_bsy_1_valid_REG_2;
  reg         stdf_clr_bsy_valid;
  reg  [6:0]  stdf_clr_bsy_rob_idx;
  reg  [19:0] stdf_clr_bsy_brmask;
  reg         casez_tmp_383;
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_383 = stq_0_valid;
      5'b00001:
        casez_tmp_383 = stq_1_valid;
      5'b00010:
        casez_tmp_383 = stq_2_valid;
      5'b00011:
        casez_tmp_383 = stq_3_valid;
      5'b00100:
        casez_tmp_383 = stq_4_valid;
      5'b00101:
        casez_tmp_383 = stq_5_valid;
      5'b00110:
        casez_tmp_383 = stq_6_valid;
      5'b00111:
        casez_tmp_383 = stq_7_valid;
      5'b01000:
        casez_tmp_383 = stq_8_valid;
      5'b01001:
        casez_tmp_383 = stq_9_valid;
      5'b01010:
        casez_tmp_383 = stq_10_valid;
      5'b01011:
        casez_tmp_383 = stq_11_valid;
      5'b01100:
        casez_tmp_383 = stq_12_valid;
      5'b01101:
        casez_tmp_383 = stq_13_valid;
      5'b01110:
        casez_tmp_383 = stq_14_valid;
      5'b01111:
        casez_tmp_383 = stq_15_valid;
      5'b10000:
        casez_tmp_383 = stq_16_valid;
      5'b10001:
        casez_tmp_383 = stq_17_valid;
      5'b10010:
        casez_tmp_383 = stq_18_valid;
      5'b10011:
        casez_tmp_383 = stq_19_valid;
      5'b10100:
        casez_tmp_383 = stq_20_valid;
      5'b10101:
        casez_tmp_383 = stq_21_valid;
      5'b10110:
        casez_tmp_383 = stq_22_valid;
      5'b10111:
        casez_tmp_383 = stq_23_valid;
      5'b11000:
        casez_tmp_383 = stq_24_valid;
      5'b11001:
        casez_tmp_383 = stq_25_valid;
      5'b11010:
        casez_tmp_383 = stq_26_valid;
      5'b11011:
        casez_tmp_383 = stq_27_valid;
      5'b11100:
        casez_tmp_383 = stq_28_valid;
      5'b11101:
        casez_tmp_383 = stq_29_valid;
      5'b11110:
        casez_tmp_383 = stq_30_valid;
      default:
        casez_tmp_383 = stq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_384;
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_384 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_384 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_384 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_384 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_384 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_384 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_384 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_384 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_384 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_384 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_384 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_384 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_384 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_384 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_384 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_384 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_384 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_384 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_384 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_384 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_384 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_384 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_384 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_384 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_384 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_384 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_384 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_384 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_384 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_384 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_384 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_384 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_385;
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_385 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_385 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_385 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_385 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_385 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_385 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_385 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_385 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_385 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_385 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_385 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_385 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_385 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_385 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_385 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_385 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_385 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_385 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_385 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_385 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_385 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_385 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_385 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_385 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_385 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_385 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_385 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_385 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_385 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_385 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_385 = stq_30_bits_addr_valid;
      default:
        casez_tmp_385 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_386;
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_386 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_386 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_386 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_386 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_386 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_386 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_386 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_386 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_386 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_386 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_386 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_386 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_386 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_386 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_386 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_386 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_386 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_386 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_386 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_386 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_386 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_386 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_386 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_386 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_386 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_386 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_386 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_386 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_386 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_386 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_386 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_386 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         io_core_clr_bsy_2_valid_REG;
  reg         io_core_clr_bsy_2_valid_REG_1;
  reg         io_core_clr_bsy_2_valid_REG_2;
  wire        do_st_search_0 = (_lcam_stq_idx_T | fired_sta_retry_REG) & ~mem_tlb_miss_0;
  wire        do_st_search_1 = (_lcam_stq_idx_T_3 | fired_sta_retry_REG_1) & ~mem_tlb_miss_1;
  wire        _can_forward_T = fired_load_incoming_REG | fired_load_retry_REG;
  wire        do_ld_search_0 = _can_forward_T & ~mem_tlb_miss_0 | fired_load_wakeup_REG;
  wire        _can_forward_T_6 = fired_load_incoming_REG_1 | fired_load_retry_REG_1;
  wire        do_ld_search_1 = _can_forward_T_6 & ~mem_tlb_miss_1 | fired_load_wakeup_REG_1;
  reg  [32:0] lcam_addr_REG;
  reg  [32:0] lcam_addr_REG_1;
  wire [39:0] lcam_addr_0 = _lcam_stq_idx_T | fired_sta_retry_REG ? {7'h0, lcam_addr_REG} : fired_release_0 ? {7'h0, lcam_addr_REG_1} : mem_paddr_0;
  reg  [32:0] lcam_addr_REG_2;
  reg  [32:0] lcam_addr_REG_3;
  wire [39:0] lcam_addr_1 = _lcam_stq_idx_T_3 | fired_sta_retry_REG_1 ? {7'h0, lcam_addr_REG_2} : fired_release_1 ? {7'h0, lcam_addr_REG_3} : mem_paddr_1;
  reg  [7:0]  casez_tmp_387;
  wire [14:0] _lcam_mask_mask_T_2 = 15'h1 << lcam_addr_0[2:0];
  wire [14:0] _lcam_mask_mask_T_6 = 15'h3 << {12'h0, lcam_addr_0[2:1], 1'h0};
  always @(*) begin
    casez (do_st_search_0 ? (_lcam_stq_idx_T ? mem_stq_incoming_e_0_bits_uop_mem_size : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_mem_size : 2'h0) : do_ld_search_0 ? (fired_load_incoming_REG ? mem_ldq_incoming_e_0_bits_uop_mem_size : fired_load_retry_REG ? mem_ldq_retry_e_bits_uop_mem_size : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_uop_mem_size : 2'h0) : 2'h0)
      2'b00:
        casez_tmp_387 = _lcam_mask_mask_T_2[7:0];
      2'b01:
        casez_tmp_387 = _lcam_mask_mask_T_6[7:0];
      2'b10:
        casez_tmp_387 = lcam_addr_0[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_387 = 8'hFF;
    endcase
  end // always @(*)
  reg  [7:0]  casez_tmp_388;
  wire [14:0] _lcam_mask_mask_T_17 = 15'h1 << lcam_addr_1[2:0];
  wire [14:0] _lcam_mask_mask_T_21 = 15'h3 << {12'h0, lcam_addr_1[2:1], 1'h0};
  always @(*) begin
    casez (do_st_search_1 ? (_lcam_stq_idx_T_3 ? mem_stq_incoming_e_1_bits_uop_mem_size : fired_sta_retry_REG_1 ? mem_stq_retry_e_bits_uop_mem_size : 2'h0) : do_ld_search_1 ? (fired_load_incoming_REG_1 ? mem_ldq_incoming_e_1_bits_uop_mem_size : fired_load_retry_REG_1 ? mem_ldq_retry_e_bits_uop_mem_size : fired_load_wakeup_REG_1 ? mem_ldq_wakeup_e_bits_uop_mem_size : 2'h0) : 2'h0)
      2'b00:
        casez_tmp_388 = _lcam_mask_mask_T_17[7:0];
      2'b01:
        casez_tmp_388 = _lcam_mask_mask_T_21[7:0];
      2'b10:
        casez_tmp_388 = lcam_addr_1[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_388 = 8'hFF;
    endcase
  end // always @(*)
  reg  [4:0]  lcam_ldq_idx_REG;
  reg  [4:0]  lcam_ldq_idx_REG_1;
  wire [4:0]  lcam_ldq_idx_0 = fired_load_incoming_REG ? mem_incoming_uop_0_ldq_idx : fired_load_wakeup_REG ? lcam_ldq_idx_REG : fired_load_retry_REG ? lcam_ldq_idx_REG_1 : 5'h0;
  reg  [4:0]  lcam_ldq_idx_REG_2;
  reg  [4:0]  lcam_ldq_idx_REG_3;
  wire [4:0]  lcam_ldq_idx_1 = fired_load_incoming_REG_1 ? mem_incoming_uop_1_ldq_idx : fired_load_wakeup_REG_1 ? lcam_ldq_idx_REG_2 : fired_load_retry_REG_1 ? lcam_ldq_idx_REG_3 : 5'h0;
  reg  [4:0]  lcam_stq_idx_REG;
  wire [4:0]  lcam_stq_idx_0 = _lcam_stq_idx_T ? mem_incoming_uop_0_stq_idx : fired_sta_retry_REG ? lcam_stq_idx_REG : 5'h0;
  reg  [4:0]  lcam_stq_idx_REG_1;
  wire [4:0]  lcam_stq_idx_1 = _lcam_stq_idx_T_3 ? mem_incoming_uop_1_stq_idx : fired_sta_retry_REG_1 ? lcam_stq_idx_REG_1 : 5'h0;
  reg         casez_tmp_389;
  always @(*) begin
    casez (lcam_ldq_idx_0)
      5'b00000:
        casez_tmp_389 = ldq_0_bits_addr_is_uncacheable;
      5'b00001:
        casez_tmp_389 = ldq_1_bits_addr_is_uncacheable;
      5'b00010:
        casez_tmp_389 = ldq_2_bits_addr_is_uncacheable;
      5'b00011:
        casez_tmp_389 = ldq_3_bits_addr_is_uncacheable;
      5'b00100:
        casez_tmp_389 = ldq_4_bits_addr_is_uncacheable;
      5'b00101:
        casez_tmp_389 = ldq_5_bits_addr_is_uncacheable;
      5'b00110:
        casez_tmp_389 = ldq_6_bits_addr_is_uncacheable;
      5'b00111:
        casez_tmp_389 = ldq_7_bits_addr_is_uncacheable;
      5'b01000:
        casez_tmp_389 = ldq_8_bits_addr_is_uncacheable;
      5'b01001:
        casez_tmp_389 = ldq_9_bits_addr_is_uncacheable;
      5'b01010:
        casez_tmp_389 = ldq_10_bits_addr_is_uncacheable;
      5'b01011:
        casez_tmp_389 = ldq_11_bits_addr_is_uncacheable;
      5'b01100:
        casez_tmp_389 = ldq_12_bits_addr_is_uncacheable;
      5'b01101:
        casez_tmp_389 = ldq_13_bits_addr_is_uncacheable;
      5'b01110:
        casez_tmp_389 = ldq_14_bits_addr_is_uncacheable;
      5'b01111:
        casez_tmp_389 = ldq_15_bits_addr_is_uncacheable;
      5'b10000:
        casez_tmp_389 = ldq_16_bits_addr_is_uncacheable;
      5'b10001:
        casez_tmp_389 = ldq_17_bits_addr_is_uncacheable;
      5'b10010:
        casez_tmp_389 = ldq_18_bits_addr_is_uncacheable;
      5'b10011:
        casez_tmp_389 = ldq_19_bits_addr_is_uncacheable;
      5'b10100:
        casez_tmp_389 = ldq_20_bits_addr_is_uncacheable;
      5'b10101:
        casez_tmp_389 = ldq_21_bits_addr_is_uncacheable;
      5'b10110:
        casez_tmp_389 = ldq_22_bits_addr_is_uncacheable;
      5'b10111:
        casez_tmp_389 = ldq_23_bits_addr_is_uncacheable;
      5'b11000:
        casez_tmp_389 = ldq_24_bits_addr_is_uncacheable;
      5'b11001:
        casez_tmp_389 = ldq_25_bits_addr_is_uncacheable;
      5'b11010:
        casez_tmp_389 = ldq_26_bits_addr_is_uncacheable;
      5'b11011:
        casez_tmp_389 = ldq_27_bits_addr_is_uncacheable;
      5'b11100:
        casez_tmp_389 = ldq_28_bits_addr_is_uncacheable;
      5'b11101:
        casez_tmp_389 = ldq_29_bits_addr_is_uncacheable;
      5'b11110:
        casez_tmp_389 = ldq_30_bits_addr_is_uncacheable;
      default:
        casez_tmp_389 = ldq_31_bits_addr_is_uncacheable;
    endcase
  end // always @(*)
  reg         casez_tmp_390;
  always @(*) begin
    casez (lcam_ldq_idx_1)
      5'b00000:
        casez_tmp_390 = ldq_0_bits_addr_is_uncacheable;
      5'b00001:
        casez_tmp_390 = ldq_1_bits_addr_is_uncacheable;
      5'b00010:
        casez_tmp_390 = ldq_2_bits_addr_is_uncacheable;
      5'b00011:
        casez_tmp_390 = ldq_3_bits_addr_is_uncacheable;
      5'b00100:
        casez_tmp_390 = ldq_4_bits_addr_is_uncacheable;
      5'b00101:
        casez_tmp_390 = ldq_5_bits_addr_is_uncacheable;
      5'b00110:
        casez_tmp_390 = ldq_6_bits_addr_is_uncacheable;
      5'b00111:
        casez_tmp_390 = ldq_7_bits_addr_is_uncacheable;
      5'b01000:
        casez_tmp_390 = ldq_8_bits_addr_is_uncacheable;
      5'b01001:
        casez_tmp_390 = ldq_9_bits_addr_is_uncacheable;
      5'b01010:
        casez_tmp_390 = ldq_10_bits_addr_is_uncacheable;
      5'b01011:
        casez_tmp_390 = ldq_11_bits_addr_is_uncacheable;
      5'b01100:
        casez_tmp_390 = ldq_12_bits_addr_is_uncacheable;
      5'b01101:
        casez_tmp_390 = ldq_13_bits_addr_is_uncacheable;
      5'b01110:
        casez_tmp_390 = ldq_14_bits_addr_is_uncacheable;
      5'b01111:
        casez_tmp_390 = ldq_15_bits_addr_is_uncacheable;
      5'b10000:
        casez_tmp_390 = ldq_16_bits_addr_is_uncacheable;
      5'b10001:
        casez_tmp_390 = ldq_17_bits_addr_is_uncacheable;
      5'b10010:
        casez_tmp_390 = ldq_18_bits_addr_is_uncacheable;
      5'b10011:
        casez_tmp_390 = ldq_19_bits_addr_is_uncacheable;
      5'b10100:
        casez_tmp_390 = ldq_20_bits_addr_is_uncacheable;
      5'b10101:
        casez_tmp_390 = ldq_21_bits_addr_is_uncacheable;
      5'b10110:
        casez_tmp_390 = ldq_22_bits_addr_is_uncacheable;
      5'b10111:
        casez_tmp_390 = ldq_23_bits_addr_is_uncacheable;
      5'b11000:
        casez_tmp_390 = ldq_24_bits_addr_is_uncacheable;
      5'b11001:
        casez_tmp_390 = ldq_25_bits_addr_is_uncacheable;
      5'b11010:
        casez_tmp_390 = ldq_26_bits_addr_is_uncacheable;
      5'b11011:
        casez_tmp_390 = ldq_27_bits_addr_is_uncacheable;
      5'b11100:
        casez_tmp_390 = ldq_28_bits_addr_is_uncacheable;
      5'b11101:
        casez_tmp_390 = ldq_29_bits_addr_is_uncacheable;
      5'b11110:
        casez_tmp_390 = ldq_30_bits_addr_is_uncacheable;
      default:
        casez_tmp_390 = ldq_31_bits_addr_is_uncacheable;
    endcase
  end // always @(*)
  reg         s1_executing_loads_0;
  reg         s1_executing_loads_1;
  reg         s1_executing_loads_2;
  reg         s1_executing_loads_3;
  reg         s1_executing_loads_4;
  reg         s1_executing_loads_5;
  reg         s1_executing_loads_6;
  reg         s1_executing_loads_7;
  reg         s1_executing_loads_8;
  reg         s1_executing_loads_9;
  reg         s1_executing_loads_10;
  reg         s1_executing_loads_11;
  reg         s1_executing_loads_12;
  reg         s1_executing_loads_13;
  reg         s1_executing_loads_14;
  reg         s1_executing_loads_15;
  reg         s1_executing_loads_16;
  reg         s1_executing_loads_17;
  reg         s1_executing_loads_18;
  reg         s1_executing_loads_19;
  reg         s1_executing_loads_20;
  reg         s1_executing_loads_21;
  reg         s1_executing_loads_22;
  reg         s1_executing_loads_23;
  reg         s1_executing_loads_24;
  reg         s1_executing_loads_25;
  reg         s1_executing_loads_26;
  reg         s1_executing_loads_27;
  reg         s1_executing_loads_28;
  reg         s1_executing_loads_29;
  reg         s1_executing_loads_30;
  reg         s1_executing_loads_31;
  reg         wb_forward_valid_0;
  reg         wb_forward_valid_1;
  reg  [4:0]  wb_forward_ldq_idx_0;
  reg  [4:0]  wb_forward_ldq_idx_1;
  reg  [39:0] wb_forward_ld_addr_0;
  reg  [39:0] wb_forward_ld_addr_1;
  reg  [4:0]  wb_forward_stq_idx_0;
  reg  [4:0]  wb_forward_stq_idx_1;
  reg  [7:0]  casez_tmp_391;
  wire [14:0] _l_mask_mask_T_2 = 15'h1 << ldq_0_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_6 = 15'h3 << {12'h0, ldq_0_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_0_bits_uop_mem_size)
      2'b00:
        casez_tmp_391 = _l_mask_mask_T_2[7:0];
      2'b01:
        casez_tmp_391 = _l_mask_mask_T_6[7:0];
      2'b10:
        casez_tmp_391 = ldq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_391 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_0 = wb_forward_valid_0 & ~(|wb_forward_ldq_idx_0);
  wire        l_forwarders_1 = wb_forward_valid_1 & ~(|wb_forward_ldq_idx_1);
  wire        l_is_forwarding = l_forwarders_0 | l_forwarders_1;
  wire [4:0]  l_forward_stq_idx = l_is_forwarding ? (l_forwarders_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_0_bits_forward_stq_idx;
  wire        block_addr_matches_0 = lcam_addr_0[39:6] == ldq_0_bits_addr_bits[39:6];
  wire        block_addr_matches_1 = lcam_addr_1[39:6] == ldq_0_bits_addr_bits[39:6];
  wire        dword_addr_matches_0 = block_addr_matches_0 & lcam_addr_0[5:3] == ldq_0_bits_addr_bits[5:3];
  wire        dword_addr_matches_1 = block_addr_matches_1 & lcam_addr_1[5:3] == ldq_0_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T = casez_tmp_391 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_2 = casez_tmp_391 & casez_tmp_388;
  wire        _GEN_284 = fired_release_0 & ldq_0_valid & ldq_0_bits_addr_valid & block_addr_matches_0;
  wire        _GEN_285 = ldq_0_bits_executed | ldq_0_bits_succeeded;
  wire        _GEN_286 = _GEN_285 | l_is_forwarding;
  wire [31:0] _GEN_287 = {27'h0, lcam_stq_idx_0};
  wire [31:0] _GEN_288 = ldq_0_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_289 = do_st_search_0 & ldq_0_valid & ldq_0_bits_addr_valid & _GEN_286 & ~ldq_0_bits_addr_is_virtual & _GEN_288[0] & dword_addr_matches_0 & (|_mask_overlap_T);
  wire        _GEN_290 = ~ldq_0_bits_forward_std_val | l_forward_stq_idx != lcam_stq_idx_0 & (l_forward_stq_idx < lcam_stq_idx_0 ^ l_forward_stq_idx < ldq_0_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_0_bits_youngest_stq_idx);
  wire        _GEN_291 = do_ld_search_0 & ldq_0_valid & ldq_0_bits_addr_valid & ~ldq_0_bits_addr_is_virtual & dword_addr_matches_0 & (|_mask_overlap_T);
  wire        searcher_is_older = lcam_ldq_idx_0 < ldq_head ^ (|ldq_head);
  wire        _GEN_292 = _GEN_286 & ~s1_executing_loads_0 & ldq_0_bits_observed;
  wire        _GEN_293 = ~_GEN_284 & (_GEN_289 ? _GEN_290 : _GEN_291 & searcher_is_older & _GEN_292);
  reg         older_nacked_REG;
  wire        _GEN_294 = ~_GEN_285 | nacking_loads_0 | older_nacked_REG;
  wire        _GEN_295 = _GEN_284 | _GEN_289;
  wire        _GEN_296 = lcam_ldq_idx_0 == 5'h1;
  wire        _GEN_297 = lcam_ldq_idx_0 == 5'h2;
  wire        _GEN_298 = lcam_ldq_idx_0 == 5'h3;
  wire        _GEN_299 = lcam_ldq_idx_0 == 5'h4;
  wire        _GEN_300 = lcam_ldq_idx_0 == 5'h5;
  wire        _GEN_301 = lcam_ldq_idx_0 == 5'h6;
  wire        _GEN_302 = lcam_ldq_idx_0 == 5'h7;
  wire        _GEN_303 = lcam_ldq_idx_0 == 5'h8;
  wire        _GEN_304 = lcam_ldq_idx_0 == 5'h9;
  wire        _GEN_305 = lcam_ldq_idx_0 == 5'hA;
  wire        _GEN_306 = lcam_ldq_idx_0 == 5'hB;
  wire        _GEN_307 = lcam_ldq_idx_0 == 5'hC;
  wire        _GEN_308 = lcam_ldq_idx_0 == 5'hD;
  wire        _GEN_309 = lcam_ldq_idx_0 == 5'hE;
  wire        _GEN_310 = lcam_ldq_idx_0 == 5'hF;
  wire        _GEN_311 = lcam_ldq_idx_0 == 5'h10;
  wire        _GEN_312 = lcam_ldq_idx_0 == 5'h11;
  wire        _GEN_313 = lcam_ldq_idx_0 == 5'h12;
  wire        _GEN_314 = lcam_ldq_idx_0 == 5'h13;
  wire        _GEN_315 = lcam_ldq_idx_0 == 5'h14;
  wire        _GEN_316 = lcam_ldq_idx_0 == 5'h15;
  wire        _GEN_317 = lcam_ldq_idx_0 == 5'h16;
  wire        _GEN_318 = lcam_ldq_idx_0 == 5'h17;
  wire        _GEN_319 = lcam_ldq_idx_0 == 5'h18;
  wire        _GEN_320 = lcam_ldq_idx_0 == 5'h19;
  wire        _GEN_321 = lcam_ldq_idx_0 == 5'h1A;
  wire        _GEN_322 = lcam_ldq_idx_0 == 5'h1B;
  wire        _GEN_323 = lcam_ldq_idx_0 == 5'h1C;
  wire        _GEN_324 = lcam_ldq_idx_0 == 5'h1D;
  wire        _GEN_325 = lcam_ldq_idx_0 == 5'h1E;
  reg         io_dmem_s1_kill_0_REG;
  wire        _GEN_326 = (|lcam_ldq_idx_0) & _GEN_294;
  wire        _GEN_327 = fired_release_1 & ldq_0_valid & ldq_0_bits_addr_valid & block_addr_matches_1;
  wire [31:0] _GEN_328 = {27'h0, lcam_stq_idx_1};
  wire [31:0] _GEN_329 = ldq_0_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_330 = do_st_search_1 & ldq_0_valid & ldq_0_bits_addr_valid & _GEN_286 & ~ldq_0_bits_addr_is_virtual & _GEN_329[0] & dword_addr_matches_1 & (|_mask_overlap_T_2);
  wire        _GEN_331 = ~ldq_0_bits_forward_std_val | l_forward_stq_idx != lcam_stq_idx_1 & (l_forward_stq_idx < lcam_stq_idx_1 ^ l_forward_stq_idx < ldq_0_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_0_bits_youngest_stq_idx);
  wire        _GEN_332 = do_ld_search_1 & ldq_0_valid & ldq_0_bits_addr_valid & ~ldq_0_bits_addr_is_virtual & dword_addr_matches_1 & (|_mask_overlap_T_2);
  wire        searcher_is_older_1 = lcam_ldq_idx_1 < ldq_head ^ (|ldq_head);
  wire        _GEN_333 = _GEN_332 & searcher_is_older_1 & _GEN_292;
  wire        _temp_bits_WIRE_1_32 = _GEN_327 ? _GEN_293 : _GEN_330 ? _GEN_331 | _GEN_293 : _GEN_333 | _GEN_293;
  reg         older_nacked_REG_1;
  wire        _GEN_334 = ~_GEN_285 | nacking_loads_0 | older_nacked_REG_1;
  wire        _GEN_335 = _GEN_327 | _GEN_330;
  wire        _GEN_336 = lcam_ldq_idx_1 == 5'h1;
  wire        _GEN_337 = lcam_ldq_idx_1 == 5'h2;
  wire        _GEN_338 = lcam_ldq_idx_1 == 5'h3;
  wire        _GEN_339 = lcam_ldq_idx_1 == 5'h4;
  wire        _GEN_340 = lcam_ldq_idx_1 == 5'h5;
  wire        _GEN_341 = lcam_ldq_idx_1 == 5'h6;
  wire        _GEN_342 = lcam_ldq_idx_1 == 5'h7;
  wire        _GEN_343 = lcam_ldq_idx_1 == 5'h8;
  wire        _GEN_344 = lcam_ldq_idx_1 == 5'h9;
  wire        _GEN_345 = lcam_ldq_idx_1 == 5'hA;
  wire        _GEN_346 = lcam_ldq_idx_1 == 5'hB;
  wire        _GEN_347 = lcam_ldq_idx_1 == 5'hC;
  wire        _GEN_348 = lcam_ldq_idx_1 == 5'hD;
  wire        _GEN_349 = lcam_ldq_idx_1 == 5'hE;
  wire        _GEN_350 = lcam_ldq_idx_1 == 5'hF;
  wire        _GEN_351 = lcam_ldq_idx_1 == 5'h10;
  wire        _GEN_352 = lcam_ldq_idx_1 == 5'h11;
  wire        _GEN_353 = lcam_ldq_idx_1 == 5'h12;
  wire        _GEN_354 = lcam_ldq_idx_1 == 5'h13;
  wire        _GEN_355 = lcam_ldq_idx_1 == 5'h14;
  wire        _GEN_356 = lcam_ldq_idx_1 == 5'h15;
  wire        _GEN_357 = lcam_ldq_idx_1 == 5'h16;
  wire        _GEN_358 = lcam_ldq_idx_1 == 5'h17;
  wire        _GEN_359 = lcam_ldq_idx_1 == 5'h18;
  wire        _GEN_360 = lcam_ldq_idx_1 == 5'h19;
  wire        _GEN_361 = lcam_ldq_idx_1 == 5'h1A;
  wire        _GEN_362 = lcam_ldq_idx_1 == 5'h1B;
  wire        _GEN_363 = lcam_ldq_idx_1 == 5'h1C;
  wire        _GEN_364 = lcam_ldq_idx_1 == 5'h1D;
  wire        _GEN_365 = lcam_ldq_idx_1 == 5'h1E;
  reg         io_dmem_s1_kill_1_REG;
  wire        _GEN_366 = (|lcam_ldq_idx_1) & _GEN_334;
  reg  [7:0]  casez_tmp_392;
  wire [14:0] _l_mask_mask_T_17 = 15'h1 << ldq_1_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_21 = 15'h3 << {12'h0, ldq_1_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_1_bits_uop_mem_size)
      2'b00:
        casez_tmp_392 = _l_mask_mask_T_17[7:0];
      2'b01:
        casez_tmp_392 = _l_mask_mask_T_21[7:0];
      2'b10:
        casez_tmp_392 = ldq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_392 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_1_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1;
  wire        l_forwarders_1_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1;
  wire        l_is_forwarding_1 = l_forwarders_1_0 | l_forwarders_1_1;
  wire [4:0]  l_forward_stq_idx_1 = l_is_forwarding_1 ? (l_forwarders_1_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_1_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_1_bits_forward_stq_idx;
  wire        block_addr_matches_1_0 = lcam_addr_0[39:6] == ldq_1_bits_addr_bits[39:6];
  wire        block_addr_matches_1_1 = lcam_addr_1[39:6] == ldq_1_bits_addr_bits[39:6];
  wire        dword_addr_matches_1_0 = block_addr_matches_1_0 & lcam_addr_0[5:3] == ldq_1_bits_addr_bits[5:3];
  wire        dword_addr_matches_1_1 = block_addr_matches_1_1 & lcam_addr_1[5:3] == ldq_1_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_4 = casez_tmp_392 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_6 = casez_tmp_392 & casez_tmp_388;
  wire        _GEN_367 = fired_release_0 & ldq_1_valid & ldq_1_bits_addr_valid & block_addr_matches_1_0;
  wire        _GEN_368 = ldq_1_bits_executed | ldq_1_bits_succeeded;
  wire        _GEN_369 = _GEN_368 | l_is_forwarding_1;
  wire [31:0] _GEN_370 = ldq_1_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_371 = do_st_search_0 & ldq_1_valid & ldq_1_bits_addr_valid & _GEN_369 & ~ldq_1_bits_addr_is_virtual & _GEN_370[0] & dword_addr_matches_1_0 & (|_mask_overlap_T_4);
  wire        _GEN_372 = ~ldq_1_bits_forward_std_val | l_forward_stq_idx_1 != lcam_stq_idx_0 & (l_forward_stq_idx_1 < lcam_stq_idx_0 ^ l_forward_stq_idx_1 < ldq_1_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_1_bits_youngest_stq_idx);
  wire        _GEN_373 = do_ld_search_0 & ldq_1_valid & ldq_1_bits_addr_valid & ~ldq_1_bits_addr_is_virtual & dword_addr_matches_1_0 & (|_mask_overlap_T_4);
  wire        searcher_is_older_2 = lcam_ldq_idx_0 == 5'h0 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[4:1]));
  wire        _GEN_374 = _GEN_369 & ~s1_executing_loads_1 & ldq_1_bits_observed;
  wire        _GEN_375 = ~_GEN_367 & (_GEN_371 ? _GEN_372 : _GEN_373 & searcher_is_older_2 & _GEN_374);
  reg         older_nacked_REG_2;
  wire        _GEN_376 = ~_GEN_368 | nacking_loads_1 | older_nacked_REG_2;
  wire        _GEN_377 = searcher_is_older_2 | _GEN_296;
  wire        _GEN_378 = _GEN_367 | _GEN_371;
  reg         io_dmem_s1_kill_0_REG_1;
  wire        _GEN_379 = _GEN_378 | ~_GEN_373 | _GEN_377 | ~_GEN_376;
  wire        _GEN_380 = fired_release_1 & ldq_1_valid & ldq_1_bits_addr_valid & block_addr_matches_1_1;
  wire [31:0] _GEN_381 = ldq_1_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_382 = do_st_search_1 & ldq_1_valid & ldq_1_bits_addr_valid & _GEN_369 & ~ldq_1_bits_addr_is_virtual & _GEN_381[0] & dword_addr_matches_1_1 & (|_mask_overlap_T_6);
  wire        _GEN_383 = ~ldq_1_bits_forward_std_val | l_forward_stq_idx_1 != lcam_stq_idx_1 & (l_forward_stq_idx_1 < lcam_stq_idx_1 ^ l_forward_stq_idx_1 < ldq_1_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_1_bits_youngest_stq_idx);
  wire        _GEN_384 = do_ld_search_1 & ldq_1_valid & ldq_1_bits_addr_valid & ~ldq_1_bits_addr_is_virtual & dword_addr_matches_1_1 & (|_mask_overlap_T_6);
  wire        searcher_is_older_3 = lcam_ldq_idx_1 == 5'h0 ^ lcam_ldq_idx_1 < ldq_head ^ (|(ldq_head[4:1]));
  wire        _GEN_385 = _GEN_384 & searcher_is_older_3 & _GEN_374;
  wire        _temp_bits_WIRE_1_33 = _GEN_380 ? _GEN_375 : _GEN_382 ? _GEN_383 | _GEN_375 : _GEN_385 | _GEN_375;
  reg         older_nacked_REG_3;
  wire        _GEN_386 = ~_GEN_368 | nacking_loads_1 | older_nacked_REG_3;
  wire        _GEN_387 = searcher_is_older_3 | _GEN_336;
  wire        _GEN_388 = _GEN_380 | _GEN_382;
  reg         io_dmem_s1_kill_1_REG_1;
  wire        _GEN_389 = _GEN_388 | ~_GEN_384 | _GEN_387 | ~_GEN_386;
  reg  [7:0]  casez_tmp_393;
  wire [14:0] _l_mask_mask_T_32 = 15'h1 << ldq_2_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_36 = 15'h3 << {12'h0, ldq_2_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_2_bits_uop_mem_size)
      2'b00:
        casez_tmp_393 = _l_mask_mask_T_32[7:0];
      2'b01:
        casez_tmp_393 = _l_mask_mask_T_36[7:0];
      2'b10:
        casez_tmp_393 = ldq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_393 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_2_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h2;
  wire        l_forwarders_2_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h2;
  wire        l_is_forwarding_2 = l_forwarders_2_0 | l_forwarders_2_1;
  wire [4:0]  l_forward_stq_idx_2 = l_is_forwarding_2 ? (l_forwarders_2_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_2_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_2_bits_forward_stq_idx;
  wire        block_addr_matches_2_0 = lcam_addr_0[39:6] == ldq_2_bits_addr_bits[39:6];
  wire        block_addr_matches_2_1 = lcam_addr_1[39:6] == ldq_2_bits_addr_bits[39:6];
  wire        dword_addr_matches_2_0 = block_addr_matches_2_0 & lcam_addr_0[5:3] == ldq_2_bits_addr_bits[5:3];
  wire        dword_addr_matches_2_1 = block_addr_matches_2_1 & lcam_addr_1[5:3] == ldq_2_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_8 = casez_tmp_393 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_10 = casez_tmp_393 & casez_tmp_388;
  wire        _GEN_390 = fired_release_0 & ldq_2_valid & ldq_2_bits_addr_valid & block_addr_matches_2_0;
  wire        _GEN_391 = ldq_2_bits_executed | ldq_2_bits_succeeded;
  wire        _GEN_392 = _GEN_391 | l_is_forwarding_2;
  wire [31:0] _GEN_393 = ldq_2_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_394 = do_st_search_0 & ldq_2_valid & ldq_2_bits_addr_valid & _GEN_392 & ~ldq_2_bits_addr_is_virtual & _GEN_393[0] & dword_addr_matches_2_0 & (|_mask_overlap_T_8);
  wire        _GEN_395 = ~ldq_2_bits_forward_std_val | l_forward_stq_idx_2 != lcam_stq_idx_0 & (l_forward_stq_idx_2 < lcam_stq_idx_0 ^ l_forward_stq_idx_2 < ldq_2_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_2_bits_youngest_stq_idx);
  wire        _GEN_396 = do_ld_search_0 & ldq_2_valid & ldq_2_bits_addr_valid & ~ldq_2_bits_addr_is_virtual & dword_addr_matches_2_0 & (|_mask_overlap_T_8);
  wire        searcher_is_older_4 = lcam_ldq_idx_0 < 5'h2 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h2;
  wire        _GEN_397 = _GEN_392 & ~s1_executing_loads_2 & ldq_2_bits_observed;
  wire        _GEN_398 = ~_GEN_390 & (_GEN_394 ? _GEN_395 : _GEN_396 & searcher_is_older_4 & _GEN_397);
  reg         older_nacked_REG_4;
  wire        _GEN_399 = ~_GEN_391 | nacking_loads_2 | older_nacked_REG_4;
  wire        _GEN_400 = searcher_is_older_4 | _GEN_297;
  wire        _GEN_401 = _GEN_390 | _GEN_394;
  reg         io_dmem_s1_kill_0_REG_2;
  wire        _GEN_402 = _GEN_401 | ~_GEN_396 | _GEN_400 | ~_GEN_399;
  wire        _GEN_403 = fired_release_1 & ldq_2_valid & ldq_2_bits_addr_valid & block_addr_matches_2_1;
  wire [31:0] _GEN_404 = ldq_2_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_405 = do_st_search_1 & ldq_2_valid & ldq_2_bits_addr_valid & _GEN_392 & ~ldq_2_bits_addr_is_virtual & _GEN_404[0] & dword_addr_matches_2_1 & (|_mask_overlap_T_10);
  wire        _GEN_406 = ~ldq_2_bits_forward_std_val | l_forward_stq_idx_2 != lcam_stq_idx_1 & (l_forward_stq_idx_2 < lcam_stq_idx_1 ^ l_forward_stq_idx_2 < ldq_2_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_2_bits_youngest_stq_idx);
  wire        _GEN_407 = do_ld_search_1 & ldq_2_valid & ldq_2_bits_addr_valid & ~ldq_2_bits_addr_is_virtual & dword_addr_matches_2_1 & (|_mask_overlap_T_10);
  wire        searcher_is_older_5 = lcam_ldq_idx_1 < 5'h2 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h2;
  wire        _GEN_408 = _GEN_407 & searcher_is_older_5 & _GEN_397;
  wire        _temp_bits_WIRE_1_34 = _GEN_403 ? _GEN_398 : _GEN_405 ? _GEN_406 | _GEN_398 : _GEN_408 | _GEN_398;
  reg         older_nacked_REG_5;
  wire        _GEN_409 = ~_GEN_391 | nacking_loads_2 | older_nacked_REG_5;
  wire        _GEN_410 = searcher_is_older_5 | _GEN_337;
  wire        _GEN_411 = _GEN_403 | _GEN_405;
  reg         io_dmem_s1_kill_1_REG_2;
  wire        _GEN_412 = _GEN_411 | ~_GEN_407 | _GEN_410 | ~_GEN_409;
  reg  [7:0]  casez_tmp_394;
  wire [14:0] _l_mask_mask_T_47 = 15'h1 << ldq_3_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_51 = 15'h3 << {12'h0, ldq_3_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_3_bits_uop_mem_size)
      2'b00:
        casez_tmp_394 = _l_mask_mask_T_47[7:0];
      2'b01:
        casez_tmp_394 = _l_mask_mask_T_51[7:0];
      2'b10:
        casez_tmp_394 = ldq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_394 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_3_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h3;
  wire        l_forwarders_3_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h3;
  wire        l_is_forwarding_3 = l_forwarders_3_0 | l_forwarders_3_1;
  wire [4:0]  l_forward_stq_idx_3 = l_is_forwarding_3 ? (l_forwarders_3_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_3_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_3_bits_forward_stq_idx;
  wire        block_addr_matches_3_0 = lcam_addr_0[39:6] == ldq_3_bits_addr_bits[39:6];
  wire        block_addr_matches_3_1 = lcam_addr_1[39:6] == ldq_3_bits_addr_bits[39:6];
  wire        dword_addr_matches_3_0 = block_addr_matches_3_0 & lcam_addr_0[5:3] == ldq_3_bits_addr_bits[5:3];
  wire        dword_addr_matches_3_1 = block_addr_matches_3_1 & lcam_addr_1[5:3] == ldq_3_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_12 = casez_tmp_394 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_14 = casez_tmp_394 & casez_tmp_388;
  wire        _GEN_413 = fired_release_0 & ldq_3_valid & ldq_3_bits_addr_valid & block_addr_matches_3_0;
  wire        _GEN_414 = ldq_3_bits_executed | ldq_3_bits_succeeded;
  wire        _GEN_415 = _GEN_414 | l_is_forwarding_3;
  wire [31:0] _GEN_416 = ldq_3_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_417 = do_st_search_0 & ldq_3_valid & ldq_3_bits_addr_valid & _GEN_415 & ~ldq_3_bits_addr_is_virtual & _GEN_416[0] & dword_addr_matches_3_0 & (|_mask_overlap_T_12);
  wire        _GEN_418 = ~ldq_3_bits_forward_std_val | l_forward_stq_idx_3 != lcam_stq_idx_0 & (l_forward_stq_idx_3 < lcam_stq_idx_0 ^ l_forward_stq_idx_3 < ldq_3_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_3_bits_youngest_stq_idx);
  wire        _GEN_419 = do_ld_search_0 & ldq_3_valid & ldq_3_bits_addr_valid & ~ldq_3_bits_addr_is_virtual & dword_addr_matches_3_0 & (|_mask_overlap_T_12);
  wire        searcher_is_older_6 = lcam_ldq_idx_0 < 5'h3 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[4:2]));
  wire        _GEN_420 = _GEN_415 & ~s1_executing_loads_3 & ldq_3_bits_observed;
  wire        _GEN_421 = ~_GEN_413 & (_GEN_417 ? _GEN_418 : _GEN_419 & searcher_is_older_6 & _GEN_420);
  reg         older_nacked_REG_6;
  wire        _GEN_422 = ~_GEN_414 | nacking_loads_3 | older_nacked_REG_6;
  wire        _GEN_423 = searcher_is_older_6 | _GEN_298;
  wire        _GEN_424 = _GEN_413 | _GEN_417;
  reg         io_dmem_s1_kill_0_REG_3;
  wire        _GEN_425 = _GEN_424 | ~_GEN_419 | _GEN_423 | ~_GEN_422;
  wire        _GEN_426 = fired_release_1 & ldq_3_valid & ldq_3_bits_addr_valid & block_addr_matches_3_1;
  wire [31:0] _GEN_427 = ldq_3_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_428 = do_st_search_1 & ldq_3_valid & ldq_3_bits_addr_valid & _GEN_415 & ~ldq_3_bits_addr_is_virtual & _GEN_427[0] & dword_addr_matches_3_1 & (|_mask_overlap_T_14);
  wire        _GEN_429 = ~ldq_3_bits_forward_std_val | l_forward_stq_idx_3 != lcam_stq_idx_1 & (l_forward_stq_idx_3 < lcam_stq_idx_1 ^ l_forward_stq_idx_3 < ldq_3_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_3_bits_youngest_stq_idx);
  wire        _GEN_430 = do_ld_search_1 & ldq_3_valid & ldq_3_bits_addr_valid & ~ldq_3_bits_addr_is_virtual & dword_addr_matches_3_1 & (|_mask_overlap_T_14);
  wire        searcher_is_older_7 = lcam_ldq_idx_1 < 5'h3 ^ lcam_ldq_idx_1 < ldq_head ^ (|(ldq_head[4:2]));
  wire        _GEN_431 = _GEN_430 & searcher_is_older_7 & _GEN_420;
  wire        _temp_bits_WIRE_1_35 = _GEN_426 ? _GEN_421 : _GEN_428 ? _GEN_429 | _GEN_421 : _GEN_431 | _GEN_421;
  reg         older_nacked_REG_7;
  wire        _GEN_432 = ~_GEN_414 | nacking_loads_3 | older_nacked_REG_7;
  wire        _GEN_433 = searcher_is_older_7 | _GEN_338;
  wire        _GEN_434 = _GEN_426 | _GEN_428;
  reg         io_dmem_s1_kill_1_REG_3;
  wire        _GEN_435 = _GEN_434 | ~_GEN_430 | _GEN_433 | ~_GEN_432;
  reg  [7:0]  casez_tmp_395;
  wire [14:0] _l_mask_mask_T_62 = 15'h1 << ldq_4_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_66 = 15'h3 << {12'h0, ldq_4_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_4_bits_uop_mem_size)
      2'b00:
        casez_tmp_395 = _l_mask_mask_T_62[7:0];
      2'b01:
        casez_tmp_395 = _l_mask_mask_T_66[7:0];
      2'b10:
        casez_tmp_395 = ldq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_395 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_4_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h4;
  wire        l_forwarders_4_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h4;
  wire        l_is_forwarding_4 = l_forwarders_4_0 | l_forwarders_4_1;
  wire [4:0]  l_forward_stq_idx_4 = l_is_forwarding_4 ? (l_forwarders_4_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_4_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_4_bits_forward_stq_idx;
  wire        block_addr_matches_4_0 = lcam_addr_0[39:6] == ldq_4_bits_addr_bits[39:6];
  wire        block_addr_matches_4_1 = lcam_addr_1[39:6] == ldq_4_bits_addr_bits[39:6];
  wire        dword_addr_matches_4_0 = block_addr_matches_4_0 & lcam_addr_0[5:3] == ldq_4_bits_addr_bits[5:3];
  wire        dword_addr_matches_4_1 = block_addr_matches_4_1 & lcam_addr_1[5:3] == ldq_4_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_16 = casez_tmp_395 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_18 = casez_tmp_395 & casez_tmp_388;
  wire        _GEN_436 = fired_release_0 & ldq_4_valid & ldq_4_bits_addr_valid & block_addr_matches_4_0;
  wire        _GEN_437 = ldq_4_bits_executed | ldq_4_bits_succeeded;
  wire        _GEN_438 = _GEN_437 | l_is_forwarding_4;
  wire [31:0] _GEN_439 = ldq_4_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_440 = do_st_search_0 & ldq_4_valid & ldq_4_bits_addr_valid & _GEN_438 & ~ldq_4_bits_addr_is_virtual & _GEN_439[0] & dword_addr_matches_4_0 & (|_mask_overlap_T_16);
  wire        _GEN_441 = ~ldq_4_bits_forward_std_val | l_forward_stq_idx_4 != lcam_stq_idx_0 & (l_forward_stq_idx_4 < lcam_stq_idx_0 ^ l_forward_stq_idx_4 < ldq_4_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_4_bits_youngest_stq_idx);
  wire        _GEN_442 = do_ld_search_0 & ldq_4_valid & ldq_4_bits_addr_valid & ~ldq_4_bits_addr_is_virtual & dword_addr_matches_4_0 & (|_mask_overlap_T_16);
  wire        searcher_is_older_8 = lcam_ldq_idx_0 < 5'h4 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h4;
  wire        _GEN_443 = _GEN_438 & ~s1_executing_loads_4 & ldq_4_bits_observed;
  wire        _GEN_444 = ~_GEN_436 & (_GEN_440 ? _GEN_441 : _GEN_442 & searcher_is_older_8 & _GEN_443);
  reg         older_nacked_REG_8;
  wire        _GEN_445 = ~_GEN_437 | nacking_loads_4 | older_nacked_REG_8;
  wire        _GEN_446 = searcher_is_older_8 | _GEN_299;
  wire        _GEN_447 = _GEN_436 | _GEN_440;
  reg         io_dmem_s1_kill_0_REG_4;
  wire        _GEN_448 = _GEN_447 | ~_GEN_442 | _GEN_446 | ~_GEN_445;
  wire        _GEN_449 = fired_release_1 & ldq_4_valid & ldq_4_bits_addr_valid & block_addr_matches_4_1;
  wire [31:0] _GEN_450 = ldq_4_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_451 = do_st_search_1 & ldq_4_valid & ldq_4_bits_addr_valid & _GEN_438 & ~ldq_4_bits_addr_is_virtual & _GEN_450[0] & dword_addr_matches_4_1 & (|_mask_overlap_T_18);
  wire        _GEN_452 = ~ldq_4_bits_forward_std_val | l_forward_stq_idx_4 != lcam_stq_idx_1 & (l_forward_stq_idx_4 < lcam_stq_idx_1 ^ l_forward_stq_idx_4 < ldq_4_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_4_bits_youngest_stq_idx);
  wire        _GEN_453 = do_ld_search_1 & ldq_4_valid & ldq_4_bits_addr_valid & ~ldq_4_bits_addr_is_virtual & dword_addr_matches_4_1 & (|_mask_overlap_T_18);
  wire        searcher_is_older_9 = lcam_ldq_idx_1 < 5'h4 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h4;
  wire        _GEN_454 = _GEN_453 & searcher_is_older_9 & _GEN_443;
  wire        _temp_bits_WIRE_1_36 = _GEN_449 ? _GEN_444 : _GEN_451 ? _GEN_452 | _GEN_444 : _GEN_454 | _GEN_444;
  reg         older_nacked_REG_9;
  wire        _GEN_455 = ~_GEN_437 | nacking_loads_4 | older_nacked_REG_9;
  wire        _GEN_456 = searcher_is_older_9 | _GEN_339;
  wire        _GEN_457 = _GEN_449 | _GEN_451;
  reg         io_dmem_s1_kill_1_REG_4;
  wire        _GEN_458 = _GEN_457 | ~_GEN_453 | _GEN_456 | ~_GEN_455;
  reg  [7:0]  casez_tmp_396;
  wire [14:0] _l_mask_mask_T_77 = 15'h1 << ldq_5_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_81 = 15'h3 << {12'h0, ldq_5_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_5_bits_uop_mem_size)
      2'b00:
        casez_tmp_396 = _l_mask_mask_T_77[7:0];
      2'b01:
        casez_tmp_396 = _l_mask_mask_T_81[7:0];
      2'b10:
        casez_tmp_396 = ldq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_396 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_5_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h5;
  wire        l_forwarders_5_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h5;
  wire        l_is_forwarding_5 = l_forwarders_5_0 | l_forwarders_5_1;
  wire [4:0]  l_forward_stq_idx_5 = l_is_forwarding_5 ? (l_forwarders_5_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_5_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_5_bits_forward_stq_idx;
  wire        block_addr_matches_5_0 = lcam_addr_0[39:6] == ldq_5_bits_addr_bits[39:6];
  wire        block_addr_matches_5_1 = lcam_addr_1[39:6] == ldq_5_bits_addr_bits[39:6];
  wire        dword_addr_matches_5_0 = block_addr_matches_5_0 & lcam_addr_0[5:3] == ldq_5_bits_addr_bits[5:3];
  wire        dword_addr_matches_5_1 = block_addr_matches_5_1 & lcam_addr_1[5:3] == ldq_5_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_20 = casez_tmp_396 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_22 = casez_tmp_396 & casez_tmp_388;
  wire        _GEN_459 = fired_release_0 & ldq_5_valid & ldq_5_bits_addr_valid & block_addr_matches_5_0;
  wire        _GEN_460 = ldq_5_bits_executed | ldq_5_bits_succeeded;
  wire        _GEN_461 = _GEN_460 | l_is_forwarding_5;
  wire [31:0] _GEN_462 = ldq_5_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_463 = do_st_search_0 & ldq_5_valid & ldq_5_bits_addr_valid & _GEN_461 & ~ldq_5_bits_addr_is_virtual & _GEN_462[0] & dword_addr_matches_5_0 & (|_mask_overlap_T_20);
  wire        _GEN_464 = ~ldq_5_bits_forward_std_val | l_forward_stq_idx_5 != lcam_stq_idx_0 & (l_forward_stq_idx_5 < lcam_stq_idx_0 ^ l_forward_stq_idx_5 < ldq_5_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_5_bits_youngest_stq_idx);
  wire        _GEN_465 = do_ld_search_0 & ldq_5_valid & ldq_5_bits_addr_valid & ~ldq_5_bits_addr_is_virtual & dword_addr_matches_5_0 & (|_mask_overlap_T_20);
  wire        searcher_is_older_10 = lcam_ldq_idx_0 < 5'h5 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h5;
  wire        _GEN_466 = _GEN_461 & ~s1_executing_loads_5 & ldq_5_bits_observed;
  wire        _GEN_467 = ~_GEN_459 & (_GEN_463 ? _GEN_464 : _GEN_465 & searcher_is_older_10 & _GEN_466);
  reg         older_nacked_REG_10;
  wire        _GEN_468 = ~_GEN_460 | nacking_loads_5 | older_nacked_REG_10;
  wire        _GEN_469 = searcher_is_older_10 | _GEN_300;
  wire        _GEN_470 = _GEN_459 | _GEN_463;
  reg         io_dmem_s1_kill_0_REG_5;
  wire        _GEN_471 = _GEN_470 | ~_GEN_465 | _GEN_469 | ~_GEN_468;
  wire        _GEN_472 = fired_release_1 & ldq_5_valid & ldq_5_bits_addr_valid & block_addr_matches_5_1;
  wire [31:0] _GEN_473 = ldq_5_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_474 = do_st_search_1 & ldq_5_valid & ldq_5_bits_addr_valid & _GEN_461 & ~ldq_5_bits_addr_is_virtual & _GEN_473[0] & dword_addr_matches_5_1 & (|_mask_overlap_T_22);
  wire        _GEN_475 = ~ldq_5_bits_forward_std_val | l_forward_stq_idx_5 != lcam_stq_idx_1 & (l_forward_stq_idx_5 < lcam_stq_idx_1 ^ l_forward_stq_idx_5 < ldq_5_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_5_bits_youngest_stq_idx);
  wire        _GEN_476 = do_ld_search_1 & ldq_5_valid & ldq_5_bits_addr_valid & ~ldq_5_bits_addr_is_virtual & dword_addr_matches_5_1 & (|_mask_overlap_T_22);
  wire        searcher_is_older_11 = lcam_ldq_idx_1 < 5'h5 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h5;
  wire        _GEN_477 = _GEN_476 & searcher_is_older_11 & _GEN_466;
  wire        _temp_bits_WIRE_1_37 = _GEN_472 ? _GEN_467 : _GEN_474 ? _GEN_475 | _GEN_467 : _GEN_477 | _GEN_467;
  reg         older_nacked_REG_11;
  wire        _GEN_478 = ~_GEN_460 | nacking_loads_5 | older_nacked_REG_11;
  wire        _GEN_479 = searcher_is_older_11 | _GEN_340;
  wire        _GEN_480 = _GEN_472 | _GEN_474;
  reg         io_dmem_s1_kill_1_REG_5;
  wire        _GEN_481 = _GEN_480 | ~_GEN_476 | _GEN_479 | ~_GEN_478;
  reg  [7:0]  casez_tmp_397;
  wire [14:0] _l_mask_mask_T_92 = 15'h1 << ldq_6_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_96 = 15'h3 << {12'h0, ldq_6_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_6_bits_uop_mem_size)
      2'b00:
        casez_tmp_397 = _l_mask_mask_T_92[7:0];
      2'b01:
        casez_tmp_397 = _l_mask_mask_T_96[7:0];
      2'b10:
        casez_tmp_397 = ldq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_397 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_6_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h6;
  wire        l_forwarders_6_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h6;
  wire        l_is_forwarding_6 = l_forwarders_6_0 | l_forwarders_6_1;
  wire [4:0]  l_forward_stq_idx_6 = l_is_forwarding_6 ? (l_forwarders_6_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_6_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_6_bits_forward_stq_idx;
  wire        block_addr_matches_6_0 = lcam_addr_0[39:6] == ldq_6_bits_addr_bits[39:6];
  wire        block_addr_matches_6_1 = lcam_addr_1[39:6] == ldq_6_bits_addr_bits[39:6];
  wire        dword_addr_matches_6_0 = block_addr_matches_6_0 & lcam_addr_0[5:3] == ldq_6_bits_addr_bits[5:3];
  wire        dword_addr_matches_6_1 = block_addr_matches_6_1 & lcam_addr_1[5:3] == ldq_6_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_24 = casez_tmp_397 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_26 = casez_tmp_397 & casez_tmp_388;
  wire        _GEN_482 = fired_release_0 & ldq_6_valid & ldq_6_bits_addr_valid & block_addr_matches_6_0;
  wire        _GEN_483 = ldq_6_bits_executed | ldq_6_bits_succeeded;
  wire        _GEN_484 = _GEN_483 | l_is_forwarding_6;
  wire [31:0] _GEN_485 = ldq_6_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_486 = do_st_search_0 & ldq_6_valid & ldq_6_bits_addr_valid & _GEN_484 & ~ldq_6_bits_addr_is_virtual & _GEN_485[0] & dword_addr_matches_6_0 & (|_mask_overlap_T_24);
  wire        _GEN_487 = ~ldq_6_bits_forward_std_val | l_forward_stq_idx_6 != lcam_stq_idx_0 & (l_forward_stq_idx_6 < lcam_stq_idx_0 ^ l_forward_stq_idx_6 < ldq_6_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_6_bits_youngest_stq_idx);
  wire        _GEN_488 = do_ld_search_0 & ldq_6_valid & ldq_6_bits_addr_valid & ~ldq_6_bits_addr_is_virtual & dword_addr_matches_6_0 & (|_mask_overlap_T_24);
  wire        searcher_is_older_12 = lcam_ldq_idx_0 < 5'h6 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h6;
  wire        _GEN_489 = _GEN_484 & ~s1_executing_loads_6 & ldq_6_bits_observed;
  wire        _GEN_490 = ~_GEN_482 & (_GEN_486 ? _GEN_487 : _GEN_488 & searcher_is_older_12 & _GEN_489);
  reg         older_nacked_REG_12;
  wire        _GEN_491 = ~_GEN_483 | nacking_loads_6 | older_nacked_REG_12;
  wire        _GEN_492 = searcher_is_older_12 | _GEN_301;
  wire        _GEN_493 = _GEN_482 | _GEN_486;
  reg         io_dmem_s1_kill_0_REG_6;
  wire        _GEN_494 = _GEN_493 | ~_GEN_488 | _GEN_492 | ~_GEN_491;
  wire        _GEN_495 = fired_release_1 & ldq_6_valid & ldq_6_bits_addr_valid & block_addr_matches_6_1;
  wire [31:0] _GEN_496 = ldq_6_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_497 = do_st_search_1 & ldq_6_valid & ldq_6_bits_addr_valid & _GEN_484 & ~ldq_6_bits_addr_is_virtual & _GEN_496[0] & dword_addr_matches_6_1 & (|_mask_overlap_T_26);
  wire        _GEN_498 = ~ldq_6_bits_forward_std_val | l_forward_stq_idx_6 != lcam_stq_idx_1 & (l_forward_stq_idx_6 < lcam_stq_idx_1 ^ l_forward_stq_idx_6 < ldq_6_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_6_bits_youngest_stq_idx);
  wire        _GEN_499 = do_ld_search_1 & ldq_6_valid & ldq_6_bits_addr_valid & ~ldq_6_bits_addr_is_virtual & dword_addr_matches_6_1 & (|_mask_overlap_T_26);
  wire        searcher_is_older_13 = lcam_ldq_idx_1 < 5'h6 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h6;
  wire        _GEN_500 = _GEN_499 & searcher_is_older_13 & _GEN_489;
  wire        _temp_bits_WIRE_1_38 = _GEN_495 ? _GEN_490 : _GEN_497 ? _GEN_498 | _GEN_490 : _GEN_500 | _GEN_490;
  reg         older_nacked_REG_13;
  wire        _GEN_501 = ~_GEN_483 | nacking_loads_6 | older_nacked_REG_13;
  wire        _GEN_502 = searcher_is_older_13 | _GEN_341;
  wire        _GEN_503 = _GEN_495 | _GEN_497;
  reg         io_dmem_s1_kill_1_REG_6;
  wire        _GEN_504 = _GEN_503 | ~_GEN_499 | _GEN_502 | ~_GEN_501;
  reg  [7:0]  casez_tmp_398;
  wire [14:0] _l_mask_mask_T_107 = 15'h1 << ldq_7_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_111 = 15'h3 << {12'h0, ldq_7_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_7_bits_uop_mem_size)
      2'b00:
        casez_tmp_398 = _l_mask_mask_T_107[7:0];
      2'b01:
        casez_tmp_398 = _l_mask_mask_T_111[7:0];
      2'b10:
        casez_tmp_398 = ldq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_398 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_7_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h7;
  wire        l_forwarders_7_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h7;
  wire        l_is_forwarding_7 = l_forwarders_7_0 | l_forwarders_7_1;
  wire [4:0]  l_forward_stq_idx_7 = l_is_forwarding_7 ? (l_forwarders_7_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_7_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_7_bits_forward_stq_idx;
  wire        block_addr_matches_7_0 = lcam_addr_0[39:6] == ldq_7_bits_addr_bits[39:6];
  wire        block_addr_matches_7_1 = lcam_addr_1[39:6] == ldq_7_bits_addr_bits[39:6];
  wire        dword_addr_matches_7_0 = block_addr_matches_7_0 & lcam_addr_0[5:3] == ldq_7_bits_addr_bits[5:3];
  wire        dword_addr_matches_7_1 = block_addr_matches_7_1 & lcam_addr_1[5:3] == ldq_7_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_28 = casez_tmp_398 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_30 = casez_tmp_398 & casez_tmp_388;
  wire        _GEN_505 = fired_release_0 & ldq_7_valid & ldq_7_bits_addr_valid & block_addr_matches_7_0;
  wire        _GEN_506 = ldq_7_bits_executed | ldq_7_bits_succeeded;
  wire        _GEN_507 = _GEN_506 | l_is_forwarding_7;
  wire [31:0] _GEN_508 = ldq_7_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_509 = do_st_search_0 & ldq_7_valid & ldq_7_bits_addr_valid & _GEN_507 & ~ldq_7_bits_addr_is_virtual & _GEN_508[0] & dword_addr_matches_7_0 & (|_mask_overlap_T_28);
  wire        _GEN_510 = ~ldq_7_bits_forward_std_val | l_forward_stq_idx_7 != lcam_stq_idx_0 & (l_forward_stq_idx_7 < lcam_stq_idx_0 ^ l_forward_stq_idx_7 < ldq_7_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_7_bits_youngest_stq_idx);
  wire        _GEN_511 = do_ld_search_0 & ldq_7_valid & ldq_7_bits_addr_valid & ~ldq_7_bits_addr_is_virtual & dword_addr_matches_7_0 & (|_mask_overlap_T_28);
  wire        searcher_is_older_14 = lcam_ldq_idx_0 < 5'h7 ^ lcam_ldq_idx_0 < ldq_head ^ (|(ldq_head[4:3]));
  wire        _GEN_512 = _GEN_507 & ~s1_executing_loads_7 & ldq_7_bits_observed;
  wire        _GEN_513 = ~_GEN_505 & (_GEN_509 ? _GEN_510 : _GEN_511 & searcher_is_older_14 & _GEN_512);
  reg         older_nacked_REG_14;
  wire        _GEN_514 = ~_GEN_506 | nacking_loads_7 | older_nacked_REG_14;
  wire        _GEN_515 = searcher_is_older_14 | _GEN_302;
  wire        _GEN_516 = _GEN_505 | _GEN_509;
  reg         io_dmem_s1_kill_0_REG_7;
  wire        _GEN_517 = _GEN_516 | ~_GEN_511 | _GEN_515 | ~_GEN_514;
  wire        _GEN_518 = fired_release_1 & ldq_7_valid & ldq_7_bits_addr_valid & block_addr_matches_7_1;
  wire [31:0] _GEN_519 = ldq_7_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_520 = do_st_search_1 & ldq_7_valid & ldq_7_bits_addr_valid & _GEN_507 & ~ldq_7_bits_addr_is_virtual & _GEN_519[0] & dword_addr_matches_7_1 & (|_mask_overlap_T_30);
  wire        _GEN_521 = ~ldq_7_bits_forward_std_val | l_forward_stq_idx_7 != lcam_stq_idx_1 & (l_forward_stq_idx_7 < lcam_stq_idx_1 ^ l_forward_stq_idx_7 < ldq_7_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_7_bits_youngest_stq_idx);
  wire        _GEN_522 = do_ld_search_1 & ldq_7_valid & ldq_7_bits_addr_valid & ~ldq_7_bits_addr_is_virtual & dword_addr_matches_7_1 & (|_mask_overlap_T_30);
  wire        searcher_is_older_15 = lcam_ldq_idx_1 < 5'h7 ^ lcam_ldq_idx_1 < ldq_head ^ (|(ldq_head[4:3]));
  wire        _GEN_523 = _GEN_522 & searcher_is_older_15 & _GEN_512;
  wire        _temp_bits_WIRE_1_39 = _GEN_518 ? _GEN_513 : _GEN_520 ? _GEN_521 | _GEN_513 : _GEN_523 | _GEN_513;
  reg         older_nacked_REG_15;
  wire        _GEN_524 = ~_GEN_506 | nacking_loads_7 | older_nacked_REG_15;
  wire        _GEN_525 = searcher_is_older_15 | _GEN_342;
  wire        _GEN_526 = _GEN_518 | _GEN_520;
  reg         io_dmem_s1_kill_1_REG_7;
  wire        _GEN_527 = _GEN_526 | ~_GEN_522 | _GEN_525 | ~_GEN_524;
  reg  [7:0]  casez_tmp_399;
  wire [14:0] _l_mask_mask_T_122 = 15'h1 << ldq_8_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_126 = 15'h3 << {12'h0, ldq_8_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_8_bits_uop_mem_size)
      2'b00:
        casez_tmp_399 = _l_mask_mask_T_122[7:0];
      2'b01:
        casez_tmp_399 = _l_mask_mask_T_126[7:0];
      2'b10:
        casez_tmp_399 = ldq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_399 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_8_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h8;
  wire        l_forwarders_8_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h8;
  wire        l_is_forwarding_8 = l_forwarders_8_0 | l_forwarders_8_1;
  wire [4:0]  l_forward_stq_idx_8 = l_is_forwarding_8 ? (l_forwarders_8_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_8_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_8_bits_forward_stq_idx;
  wire        block_addr_matches_8_0 = lcam_addr_0[39:6] == ldq_8_bits_addr_bits[39:6];
  wire        block_addr_matches_8_1 = lcam_addr_1[39:6] == ldq_8_bits_addr_bits[39:6];
  wire        dword_addr_matches_8_0 = block_addr_matches_8_0 & lcam_addr_0[5:3] == ldq_8_bits_addr_bits[5:3];
  wire        dword_addr_matches_8_1 = block_addr_matches_8_1 & lcam_addr_1[5:3] == ldq_8_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_32 = casez_tmp_399 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_34 = casez_tmp_399 & casez_tmp_388;
  wire        _GEN_528 = fired_release_0 & ldq_8_valid & ldq_8_bits_addr_valid & block_addr_matches_8_0;
  wire        _GEN_529 = ldq_8_bits_executed | ldq_8_bits_succeeded;
  wire        _GEN_530 = _GEN_529 | l_is_forwarding_8;
  wire [31:0] _GEN_531 = ldq_8_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_532 = do_st_search_0 & ldq_8_valid & ldq_8_bits_addr_valid & _GEN_530 & ~ldq_8_bits_addr_is_virtual & _GEN_531[0] & dword_addr_matches_8_0 & (|_mask_overlap_T_32);
  wire        _GEN_533 = ~ldq_8_bits_forward_std_val | l_forward_stq_idx_8 != lcam_stq_idx_0 & (l_forward_stq_idx_8 < lcam_stq_idx_0 ^ l_forward_stq_idx_8 < ldq_8_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_8_bits_youngest_stq_idx);
  wire        _GEN_534 = do_ld_search_0 & ldq_8_valid & ldq_8_bits_addr_valid & ~ldq_8_bits_addr_is_virtual & dword_addr_matches_8_0 & (|_mask_overlap_T_32);
  wire        searcher_is_older_16 = lcam_ldq_idx_0 < 5'h8 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h8;
  wire        _GEN_535 = _GEN_530 & ~s1_executing_loads_8 & ldq_8_bits_observed;
  wire        _GEN_536 = ~_GEN_528 & (_GEN_532 ? _GEN_533 : _GEN_534 & searcher_is_older_16 & _GEN_535);
  reg         older_nacked_REG_16;
  wire        _GEN_537 = ~_GEN_529 | nacking_loads_8 | older_nacked_REG_16;
  wire        _GEN_538 = searcher_is_older_16 | _GEN_303;
  wire        _GEN_539 = _GEN_528 | _GEN_532;
  reg         io_dmem_s1_kill_0_REG_8;
  wire        _GEN_540 = _GEN_539 | ~_GEN_534 | _GEN_538 | ~_GEN_537;
  wire        _GEN_541 = fired_release_1 & ldq_8_valid & ldq_8_bits_addr_valid & block_addr_matches_8_1;
  wire [31:0] _GEN_542 = ldq_8_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_543 = do_st_search_1 & ldq_8_valid & ldq_8_bits_addr_valid & _GEN_530 & ~ldq_8_bits_addr_is_virtual & _GEN_542[0] & dword_addr_matches_8_1 & (|_mask_overlap_T_34);
  wire        _GEN_544 = ~ldq_8_bits_forward_std_val | l_forward_stq_idx_8 != lcam_stq_idx_1 & (l_forward_stq_idx_8 < lcam_stq_idx_1 ^ l_forward_stq_idx_8 < ldq_8_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_8_bits_youngest_stq_idx);
  wire        _GEN_545 = do_ld_search_1 & ldq_8_valid & ldq_8_bits_addr_valid & ~ldq_8_bits_addr_is_virtual & dword_addr_matches_8_1 & (|_mask_overlap_T_34);
  wire        searcher_is_older_17 = lcam_ldq_idx_1 < 5'h8 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h8;
  wire        _GEN_546 = _GEN_545 & searcher_is_older_17 & _GEN_535;
  wire        _temp_bits_WIRE_1_40 = _GEN_541 ? _GEN_536 : _GEN_543 ? _GEN_544 | _GEN_536 : _GEN_546 | _GEN_536;
  reg         older_nacked_REG_17;
  wire        _GEN_547 = ~_GEN_529 | nacking_loads_8 | older_nacked_REG_17;
  wire        _GEN_548 = searcher_is_older_17 | _GEN_343;
  wire        _GEN_549 = _GEN_541 | _GEN_543;
  reg         io_dmem_s1_kill_1_REG_8;
  wire        _GEN_550 = _GEN_549 | ~_GEN_545 | _GEN_548 | ~_GEN_547;
  reg  [7:0]  casez_tmp_400;
  wire [14:0] _l_mask_mask_T_137 = 15'h1 << ldq_9_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_141 = 15'h3 << {12'h0, ldq_9_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_9_bits_uop_mem_size)
      2'b00:
        casez_tmp_400 = _l_mask_mask_T_137[7:0];
      2'b01:
        casez_tmp_400 = _l_mask_mask_T_141[7:0];
      2'b10:
        casez_tmp_400 = ldq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_400 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_9_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h9;
  wire        l_forwarders_9_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h9;
  wire        l_is_forwarding_9 = l_forwarders_9_0 | l_forwarders_9_1;
  wire [4:0]  l_forward_stq_idx_9 = l_is_forwarding_9 ? (l_forwarders_9_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_9_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_9_bits_forward_stq_idx;
  wire        block_addr_matches_9_0 = lcam_addr_0[39:6] == ldq_9_bits_addr_bits[39:6];
  wire        block_addr_matches_9_1 = lcam_addr_1[39:6] == ldq_9_bits_addr_bits[39:6];
  wire        dword_addr_matches_9_0 = block_addr_matches_9_0 & lcam_addr_0[5:3] == ldq_9_bits_addr_bits[5:3];
  wire        dword_addr_matches_9_1 = block_addr_matches_9_1 & lcam_addr_1[5:3] == ldq_9_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_36 = casez_tmp_400 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_38 = casez_tmp_400 & casez_tmp_388;
  wire        _GEN_551 = fired_release_0 & ldq_9_valid & ldq_9_bits_addr_valid & block_addr_matches_9_0;
  wire        _GEN_552 = ldq_9_bits_executed | ldq_9_bits_succeeded;
  wire        _GEN_553 = _GEN_552 | l_is_forwarding_9;
  wire [31:0] _GEN_554 = ldq_9_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_555 = do_st_search_0 & ldq_9_valid & ldq_9_bits_addr_valid & _GEN_553 & ~ldq_9_bits_addr_is_virtual & _GEN_554[0] & dword_addr_matches_9_0 & (|_mask_overlap_T_36);
  wire        _GEN_556 = ~ldq_9_bits_forward_std_val | l_forward_stq_idx_9 != lcam_stq_idx_0 & (l_forward_stq_idx_9 < lcam_stq_idx_0 ^ l_forward_stq_idx_9 < ldq_9_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_9_bits_youngest_stq_idx);
  wire        _GEN_557 = do_ld_search_0 & ldq_9_valid & ldq_9_bits_addr_valid & ~ldq_9_bits_addr_is_virtual & dword_addr_matches_9_0 & (|_mask_overlap_T_36);
  wire        searcher_is_older_18 = lcam_ldq_idx_0 < 5'h9 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h9;
  wire        _GEN_558 = _GEN_553 & ~s1_executing_loads_9 & ldq_9_bits_observed;
  wire        _GEN_559 = ~_GEN_551 & (_GEN_555 ? _GEN_556 : _GEN_557 & searcher_is_older_18 & _GEN_558);
  reg         older_nacked_REG_18;
  wire        _GEN_560 = ~_GEN_552 | nacking_loads_9 | older_nacked_REG_18;
  wire        _GEN_561 = searcher_is_older_18 | _GEN_304;
  wire        _GEN_562 = _GEN_551 | _GEN_555;
  reg         io_dmem_s1_kill_0_REG_9;
  wire        _GEN_563 = _GEN_562 | ~_GEN_557 | _GEN_561 | ~_GEN_560;
  wire        _GEN_564 = fired_release_1 & ldq_9_valid & ldq_9_bits_addr_valid & block_addr_matches_9_1;
  wire [31:0] _GEN_565 = ldq_9_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_566 = do_st_search_1 & ldq_9_valid & ldq_9_bits_addr_valid & _GEN_553 & ~ldq_9_bits_addr_is_virtual & _GEN_565[0] & dword_addr_matches_9_1 & (|_mask_overlap_T_38);
  wire        _GEN_567 = ~ldq_9_bits_forward_std_val | l_forward_stq_idx_9 != lcam_stq_idx_1 & (l_forward_stq_idx_9 < lcam_stq_idx_1 ^ l_forward_stq_idx_9 < ldq_9_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_9_bits_youngest_stq_idx);
  wire        _GEN_568 = do_ld_search_1 & ldq_9_valid & ldq_9_bits_addr_valid & ~ldq_9_bits_addr_is_virtual & dword_addr_matches_9_1 & (|_mask_overlap_T_38);
  wire        searcher_is_older_19 = lcam_ldq_idx_1 < 5'h9 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h9;
  wire        _GEN_569 = _GEN_568 & searcher_is_older_19 & _GEN_558;
  wire        _temp_bits_WIRE_1_41 = _GEN_564 ? _GEN_559 : _GEN_566 ? _GEN_567 | _GEN_559 : _GEN_569 | _GEN_559;
  reg         older_nacked_REG_19;
  wire        _GEN_570 = ~_GEN_552 | nacking_loads_9 | older_nacked_REG_19;
  wire        _GEN_571 = searcher_is_older_19 | _GEN_344;
  wire        _GEN_572 = _GEN_564 | _GEN_566;
  reg         io_dmem_s1_kill_1_REG_9;
  wire        _GEN_573 = _GEN_572 | ~_GEN_568 | _GEN_571 | ~_GEN_570;
  reg  [7:0]  casez_tmp_401;
  wire [14:0] _l_mask_mask_T_152 = 15'h1 << ldq_10_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_156 = 15'h3 << {12'h0, ldq_10_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_10_bits_uop_mem_size)
      2'b00:
        casez_tmp_401 = _l_mask_mask_T_152[7:0];
      2'b01:
        casez_tmp_401 = _l_mask_mask_T_156[7:0];
      2'b10:
        casez_tmp_401 = ldq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_401 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_10_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hA;
  wire        l_forwarders_10_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hA;
  wire        l_is_forwarding_10 = l_forwarders_10_0 | l_forwarders_10_1;
  wire [4:0]  l_forward_stq_idx_10 = l_is_forwarding_10 ? (l_forwarders_10_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_10_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_10_bits_forward_stq_idx;
  wire        block_addr_matches_10_0 = lcam_addr_0[39:6] == ldq_10_bits_addr_bits[39:6];
  wire        block_addr_matches_10_1 = lcam_addr_1[39:6] == ldq_10_bits_addr_bits[39:6];
  wire        dword_addr_matches_10_0 = block_addr_matches_10_0 & lcam_addr_0[5:3] == ldq_10_bits_addr_bits[5:3];
  wire        dword_addr_matches_10_1 = block_addr_matches_10_1 & lcam_addr_1[5:3] == ldq_10_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_40 = casez_tmp_401 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_42 = casez_tmp_401 & casez_tmp_388;
  wire        _GEN_574 = fired_release_0 & ldq_10_valid & ldq_10_bits_addr_valid & block_addr_matches_10_0;
  wire        _GEN_575 = ldq_10_bits_executed | ldq_10_bits_succeeded;
  wire        _GEN_576 = _GEN_575 | l_is_forwarding_10;
  wire [31:0] _GEN_577 = ldq_10_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_578 = do_st_search_0 & ldq_10_valid & ldq_10_bits_addr_valid & _GEN_576 & ~ldq_10_bits_addr_is_virtual & _GEN_577[0] & dword_addr_matches_10_0 & (|_mask_overlap_T_40);
  wire        _GEN_579 = ~ldq_10_bits_forward_std_val | l_forward_stq_idx_10 != lcam_stq_idx_0 & (l_forward_stq_idx_10 < lcam_stq_idx_0 ^ l_forward_stq_idx_10 < ldq_10_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_10_bits_youngest_stq_idx);
  wire        _GEN_580 = do_ld_search_0 & ldq_10_valid & ldq_10_bits_addr_valid & ~ldq_10_bits_addr_is_virtual & dword_addr_matches_10_0 & (|_mask_overlap_T_40);
  wire        searcher_is_older_20 = lcam_ldq_idx_0 < 5'hA ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hA;
  wire        _GEN_581 = _GEN_576 & ~s1_executing_loads_10 & ldq_10_bits_observed;
  wire        _GEN_582 = ~_GEN_574 & (_GEN_578 ? _GEN_579 : _GEN_580 & searcher_is_older_20 & _GEN_581);
  reg         older_nacked_REG_20;
  wire        _GEN_583 = ~_GEN_575 | nacking_loads_10 | older_nacked_REG_20;
  wire        _GEN_584 = searcher_is_older_20 | _GEN_305;
  wire        _GEN_585 = _GEN_574 | _GEN_578;
  reg         io_dmem_s1_kill_0_REG_10;
  wire        _GEN_586 = _GEN_585 | ~_GEN_580 | _GEN_584 | ~_GEN_583;
  wire        _GEN_587 = fired_release_1 & ldq_10_valid & ldq_10_bits_addr_valid & block_addr_matches_10_1;
  wire [31:0] _GEN_588 = ldq_10_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_589 = do_st_search_1 & ldq_10_valid & ldq_10_bits_addr_valid & _GEN_576 & ~ldq_10_bits_addr_is_virtual & _GEN_588[0] & dword_addr_matches_10_1 & (|_mask_overlap_T_42);
  wire        _GEN_590 = ~ldq_10_bits_forward_std_val | l_forward_stq_idx_10 != lcam_stq_idx_1 & (l_forward_stq_idx_10 < lcam_stq_idx_1 ^ l_forward_stq_idx_10 < ldq_10_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_10_bits_youngest_stq_idx);
  wire        _GEN_591 = do_ld_search_1 & ldq_10_valid & ldq_10_bits_addr_valid & ~ldq_10_bits_addr_is_virtual & dword_addr_matches_10_1 & (|_mask_overlap_T_42);
  wire        searcher_is_older_21 = lcam_ldq_idx_1 < 5'hA ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'hA;
  wire        _GEN_592 = _GEN_591 & searcher_is_older_21 & _GEN_581;
  wire        _temp_bits_WIRE_1_42 = _GEN_587 ? _GEN_582 : _GEN_589 ? _GEN_590 | _GEN_582 : _GEN_592 | _GEN_582;
  reg         older_nacked_REG_21;
  wire        _GEN_593 = ~_GEN_575 | nacking_loads_10 | older_nacked_REG_21;
  wire        _GEN_594 = searcher_is_older_21 | _GEN_345;
  wire        _GEN_595 = _GEN_587 | _GEN_589;
  reg         io_dmem_s1_kill_1_REG_10;
  wire        _GEN_596 = _GEN_595 | ~_GEN_591 | _GEN_594 | ~_GEN_593;
  reg  [7:0]  casez_tmp_402;
  wire [14:0] _l_mask_mask_T_167 = 15'h1 << ldq_11_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_171 = 15'h3 << {12'h0, ldq_11_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_11_bits_uop_mem_size)
      2'b00:
        casez_tmp_402 = _l_mask_mask_T_167[7:0];
      2'b01:
        casez_tmp_402 = _l_mask_mask_T_171[7:0];
      2'b10:
        casez_tmp_402 = ldq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_402 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_11_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hB;
  wire        l_forwarders_11_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hB;
  wire        l_is_forwarding_11 = l_forwarders_11_0 | l_forwarders_11_1;
  wire [4:0]  l_forward_stq_idx_11 = l_is_forwarding_11 ? (l_forwarders_11_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_11_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_11_bits_forward_stq_idx;
  wire        block_addr_matches_11_0 = lcam_addr_0[39:6] == ldq_11_bits_addr_bits[39:6];
  wire        block_addr_matches_11_1 = lcam_addr_1[39:6] == ldq_11_bits_addr_bits[39:6];
  wire        dword_addr_matches_11_0 = block_addr_matches_11_0 & lcam_addr_0[5:3] == ldq_11_bits_addr_bits[5:3];
  wire        dword_addr_matches_11_1 = block_addr_matches_11_1 & lcam_addr_1[5:3] == ldq_11_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_44 = casez_tmp_402 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_46 = casez_tmp_402 & casez_tmp_388;
  wire        _GEN_597 = fired_release_0 & ldq_11_valid & ldq_11_bits_addr_valid & block_addr_matches_11_0;
  wire        _GEN_598 = ldq_11_bits_executed | ldq_11_bits_succeeded;
  wire        _GEN_599 = _GEN_598 | l_is_forwarding_11;
  wire [31:0] _GEN_600 = ldq_11_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_601 = do_st_search_0 & ldq_11_valid & ldq_11_bits_addr_valid & _GEN_599 & ~ldq_11_bits_addr_is_virtual & _GEN_600[0] & dword_addr_matches_11_0 & (|_mask_overlap_T_44);
  wire        _GEN_602 = ~ldq_11_bits_forward_std_val | l_forward_stq_idx_11 != lcam_stq_idx_0 & (l_forward_stq_idx_11 < lcam_stq_idx_0 ^ l_forward_stq_idx_11 < ldq_11_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_11_bits_youngest_stq_idx);
  wire        _GEN_603 = do_ld_search_0 & ldq_11_valid & ldq_11_bits_addr_valid & ~ldq_11_bits_addr_is_virtual & dword_addr_matches_11_0 & (|_mask_overlap_T_44);
  wire        searcher_is_older_22 = lcam_ldq_idx_0 < 5'hB ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hB;
  wire        _GEN_604 = _GEN_599 & ~s1_executing_loads_11 & ldq_11_bits_observed;
  wire        _GEN_605 = ~_GEN_597 & (_GEN_601 ? _GEN_602 : _GEN_603 & searcher_is_older_22 & _GEN_604);
  reg         older_nacked_REG_22;
  wire        _GEN_606 = ~_GEN_598 | nacking_loads_11 | older_nacked_REG_22;
  wire        _GEN_607 = searcher_is_older_22 | _GEN_306;
  wire        _GEN_608 = _GEN_597 | _GEN_601;
  reg         io_dmem_s1_kill_0_REG_11;
  wire        _GEN_609 = _GEN_608 | ~_GEN_603 | _GEN_607 | ~_GEN_606;
  wire        _GEN_610 = fired_release_1 & ldq_11_valid & ldq_11_bits_addr_valid & block_addr_matches_11_1;
  wire [31:0] _GEN_611 = ldq_11_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_612 = do_st_search_1 & ldq_11_valid & ldq_11_bits_addr_valid & _GEN_599 & ~ldq_11_bits_addr_is_virtual & _GEN_611[0] & dword_addr_matches_11_1 & (|_mask_overlap_T_46);
  wire        _GEN_613 = ~ldq_11_bits_forward_std_val | l_forward_stq_idx_11 != lcam_stq_idx_1 & (l_forward_stq_idx_11 < lcam_stq_idx_1 ^ l_forward_stq_idx_11 < ldq_11_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_11_bits_youngest_stq_idx);
  wire        _GEN_614 = do_ld_search_1 & ldq_11_valid & ldq_11_bits_addr_valid & ~ldq_11_bits_addr_is_virtual & dword_addr_matches_11_1 & (|_mask_overlap_T_46);
  wire        searcher_is_older_23 = lcam_ldq_idx_1 < 5'hB ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'hB;
  wire        _GEN_615 = _GEN_614 & searcher_is_older_23 & _GEN_604;
  wire        _temp_bits_WIRE_1_43 = _GEN_610 ? _GEN_605 : _GEN_612 ? _GEN_613 | _GEN_605 : _GEN_615 | _GEN_605;
  reg         older_nacked_REG_23;
  wire        _GEN_616 = ~_GEN_598 | nacking_loads_11 | older_nacked_REG_23;
  wire        _GEN_617 = searcher_is_older_23 | _GEN_346;
  wire        _GEN_618 = _GEN_610 | _GEN_612;
  reg         io_dmem_s1_kill_1_REG_11;
  wire        _GEN_619 = _GEN_618 | ~_GEN_614 | _GEN_617 | ~_GEN_616;
  reg  [7:0]  casez_tmp_403;
  wire [14:0] _l_mask_mask_T_182 = 15'h1 << ldq_12_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_186 = 15'h3 << {12'h0, ldq_12_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_12_bits_uop_mem_size)
      2'b00:
        casez_tmp_403 = _l_mask_mask_T_182[7:0];
      2'b01:
        casez_tmp_403 = _l_mask_mask_T_186[7:0];
      2'b10:
        casez_tmp_403 = ldq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_403 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_12_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hC;
  wire        l_forwarders_12_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hC;
  wire        l_is_forwarding_12 = l_forwarders_12_0 | l_forwarders_12_1;
  wire [4:0]  l_forward_stq_idx_12 = l_is_forwarding_12 ? (l_forwarders_12_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_12_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_12_bits_forward_stq_idx;
  wire        block_addr_matches_12_0 = lcam_addr_0[39:6] == ldq_12_bits_addr_bits[39:6];
  wire        block_addr_matches_12_1 = lcam_addr_1[39:6] == ldq_12_bits_addr_bits[39:6];
  wire        dword_addr_matches_12_0 = block_addr_matches_12_0 & lcam_addr_0[5:3] == ldq_12_bits_addr_bits[5:3];
  wire        dword_addr_matches_12_1 = block_addr_matches_12_1 & lcam_addr_1[5:3] == ldq_12_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_48 = casez_tmp_403 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_50 = casez_tmp_403 & casez_tmp_388;
  wire        _GEN_620 = fired_release_0 & ldq_12_valid & ldq_12_bits_addr_valid & block_addr_matches_12_0;
  wire        _GEN_621 = ldq_12_bits_executed | ldq_12_bits_succeeded;
  wire        _GEN_622 = _GEN_621 | l_is_forwarding_12;
  wire [31:0] _GEN_623 = ldq_12_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_624 = do_st_search_0 & ldq_12_valid & ldq_12_bits_addr_valid & _GEN_622 & ~ldq_12_bits_addr_is_virtual & _GEN_623[0] & dword_addr_matches_12_0 & (|_mask_overlap_T_48);
  wire        _GEN_625 = ~ldq_12_bits_forward_std_val | l_forward_stq_idx_12 != lcam_stq_idx_0 & (l_forward_stq_idx_12 < lcam_stq_idx_0 ^ l_forward_stq_idx_12 < ldq_12_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_12_bits_youngest_stq_idx);
  wire        _GEN_626 = do_ld_search_0 & ldq_12_valid & ldq_12_bits_addr_valid & ~ldq_12_bits_addr_is_virtual & dword_addr_matches_12_0 & (|_mask_overlap_T_48);
  wire        searcher_is_older_24 = lcam_ldq_idx_0 < 5'hC ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hC;
  wire        _GEN_627 = _GEN_622 & ~s1_executing_loads_12 & ldq_12_bits_observed;
  wire        _GEN_628 = ~_GEN_620 & (_GEN_624 ? _GEN_625 : _GEN_626 & searcher_is_older_24 & _GEN_627);
  reg         older_nacked_REG_24;
  wire        _GEN_629 = ~_GEN_621 | nacking_loads_12 | older_nacked_REG_24;
  wire        _GEN_630 = searcher_is_older_24 | _GEN_307;
  wire        _GEN_631 = _GEN_620 | _GEN_624;
  reg         io_dmem_s1_kill_0_REG_12;
  wire        _GEN_632 = _GEN_631 | ~_GEN_626 | _GEN_630 | ~_GEN_629;
  wire        _GEN_633 = fired_release_1 & ldq_12_valid & ldq_12_bits_addr_valid & block_addr_matches_12_1;
  wire [31:0] _GEN_634 = ldq_12_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_635 = do_st_search_1 & ldq_12_valid & ldq_12_bits_addr_valid & _GEN_622 & ~ldq_12_bits_addr_is_virtual & _GEN_634[0] & dword_addr_matches_12_1 & (|_mask_overlap_T_50);
  wire        _GEN_636 = ~ldq_12_bits_forward_std_val | l_forward_stq_idx_12 != lcam_stq_idx_1 & (l_forward_stq_idx_12 < lcam_stq_idx_1 ^ l_forward_stq_idx_12 < ldq_12_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_12_bits_youngest_stq_idx);
  wire        _GEN_637 = do_ld_search_1 & ldq_12_valid & ldq_12_bits_addr_valid & ~ldq_12_bits_addr_is_virtual & dword_addr_matches_12_1 & (|_mask_overlap_T_50);
  wire        searcher_is_older_25 = lcam_ldq_idx_1 < 5'hC ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'hC;
  wire        _GEN_638 = _GEN_637 & searcher_is_older_25 & _GEN_627;
  wire        _temp_bits_WIRE_1_44 = _GEN_633 ? _GEN_628 : _GEN_635 ? _GEN_636 | _GEN_628 : _GEN_638 | _GEN_628;
  reg         older_nacked_REG_25;
  wire        _GEN_639 = ~_GEN_621 | nacking_loads_12 | older_nacked_REG_25;
  wire        _GEN_640 = searcher_is_older_25 | _GEN_347;
  wire        _GEN_641 = _GEN_633 | _GEN_635;
  reg         io_dmem_s1_kill_1_REG_12;
  wire        _GEN_642 = _GEN_641 | ~_GEN_637 | _GEN_640 | ~_GEN_639;
  reg  [7:0]  casez_tmp_404;
  wire [14:0] _l_mask_mask_T_197 = 15'h1 << ldq_13_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_201 = 15'h3 << {12'h0, ldq_13_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_13_bits_uop_mem_size)
      2'b00:
        casez_tmp_404 = _l_mask_mask_T_197[7:0];
      2'b01:
        casez_tmp_404 = _l_mask_mask_T_201[7:0];
      2'b10:
        casez_tmp_404 = ldq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_404 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_13_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hD;
  wire        l_forwarders_13_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hD;
  wire        l_is_forwarding_13 = l_forwarders_13_0 | l_forwarders_13_1;
  wire [4:0]  l_forward_stq_idx_13 = l_is_forwarding_13 ? (l_forwarders_13_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_13_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_13_bits_forward_stq_idx;
  wire        block_addr_matches_13_0 = lcam_addr_0[39:6] == ldq_13_bits_addr_bits[39:6];
  wire        block_addr_matches_13_1 = lcam_addr_1[39:6] == ldq_13_bits_addr_bits[39:6];
  wire        dword_addr_matches_13_0 = block_addr_matches_13_0 & lcam_addr_0[5:3] == ldq_13_bits_addr_bits[5:3];
  wire        dword_addr_matches_13_1 = block_addr_matches_13_1 & lcam_addr_1[5:3] == ldq_13_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_52 = casez_tmp_404 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_54 = casez_tmp_404 & casez_tmp_388;
  wire        _GEN_643 = fired_release_0 & ldq_13_valid & ldq_13_bits_addr_valid & block_addr_matches_13_0;
  wire        _GEN_644 = ldq_13_bits_executed | ldq_13_bits_succeeded;
  wire        _GEN_645 = _GEN_644 | l_is_forwarding_13;
  wire [31:0] _GEN_646 = ldq_13_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_647 = do_st_search_0 & ldq_13_valid & ldq_13_bits_addr_valid & _GEN_645 & ~ldq_13_bits_addr_is_virtual & _GEN_646[0] & dword_addr_matches_13_0 & (|_mask_overlap_T_52);
  wire        _GEN_648 = ~ldq_13_bits_forward_std_val | l_forward_stq_idx_13 != lcam_stq_idx_0 & (l_forward_stq_idx_13 < lcam_stq_idx_0 ^ l_forward_stq_idx_13 < ldq_13_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_13_bits_youngest_stq_idx);
  wire        _GEN_649 = do_ld_search_0 & ldq_13_valid & ldq_13_bits_addr_valid & ~ldq_13_bits_addr_is_virtual & dword_addr_matches_13_0 & (|_mask_overlap_T_52);
  wire        searcher_is_older_26 = lcam_ldq_idx_0 < 5'hD ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hD;
  wire        _GEN_650 = _GEN_645 & ~s1_executing_loads_13 & ldq_13_bits_observed;
  wire        _GEN_651 = ~_GEN_643 & (_GEN_647 ? _GEN_648 : _GEN_649 & searcher_is_older_26 & _GEN_650);
  reg         older_nacked_REG_26;
  wire        _GEN_652 = ~_GEN_644 | nacking_loads_13 | older_nacked_REG_26;
  wire        _GEN_653 = searcher_is_older_26 | _GEN_308;
  wire        _GEN_654 = _GEN_643 | _GEN_647;
  reg         io_dmem_s1_kill_0_REG_13;
  wire        _GEN_655 = _GEN_654 | ~_GEN_649 | _GEN_653 | ~_GEN_652;
  wire        _GEN_656 = fired_release_1 & ldq_13_valid & ldq_13_bits_addr_valid & block_addr_matches_13_1;
  wire [31:0] _GEN_657 = ldq_13_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_658 = do_st_search_1 & ldq_13_valid & ldq_13_bits_addr_valid & _GEN_645 & ~ldq_13_bits_addr_is_virtual & _GEN_657[0] & dword_addr_matches_13_1 & (|_mask_overlap_T_54);
  wire        _GEN_659 = ~ldq_13_bits_forward_std_val | l_forward_stq_idx_13 != lcam_stq_idx_1 & (l_forward_stq_idx_13 < lcam_stq_idx_1 ^ l_forward_stq_idx_13 < ldq_13_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_13_bits_youngest_stq_idx);
  wire        _GEN_660 = do_ld_search_1 & ldq_13_valid & ldq_13_bits_addr_valid & ~ldq_13_bits_addr_is_virtual & dword_addr_matches_13_1 & (|_mask_overlap_T_54);
  wire        searcher_is_older_27 = lcam_ldq_idx_1 < 5'hD ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'hD;
  wire        _GEN_661 = _GEN_660 & searcher_is_older_27 & _GEN_650;
  wire        _temp_bits_WIRE_1_45 = _GEN_656 ? _GEN_651 : _GEN_658 ? _GEN_659 | _GEN_651 : _GEN_661 | _GEN_651;
  reg         older_nacked_REG_27;
  wire        _GEN_662 = ~_GEN_644 | nacking_loads_13 | older_nacked_REG_27;
  wire        _GEN_663 = searcher_is_older_27 | _GEN_348;
  wire        _GEN_664 = _GEN_656 | _GEN_658;
  reg         io_dmem_s1_kill_1_REG_13;
  wire        _GEN_665 = _GEN_664 | ~_GEN_660 | _GEN_663 | ~_GEN_662;
  reg  [7:0]  casez_tmp_405;
  wire [14:0] _l_mask_mask_T_212 = 15'h1 << ldq_14_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_216 = 15'h3 << {12'h0, ldq_14_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_14_bits_uop_mem_size)
      2'b00:
        casez_tmp_405 = _l_mask_mask_T_212[7:0];
      2'b01:
        casez_tmp_405 = _l_mask_mask_T_216[7:0];
      2'b10:
        casez_tmp_405 = ldq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_405 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_14_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hE;
  wire        l_forwarders_14_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hE;
  wire        l_is_forwarding_14 = l_forwarders_14_0 | l_forwarders_14_1;
  wire [4:0]  l_forward_stq_idx_14 = l_is_forwarding_14 ? (l_forwarders_14_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_14_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_14_bits_forward_stq_idx;
  wire        block_addr_matches_14_0 = lcam_addr_0[39:6] == ldq_14_bits_addr_bits[39:6];
  wire        block_addr_matches_14_1 = lcam_addr_1[39:6] == ldq_14_bits_addr_bits[39:6];
  wire        dword_addr_matches_14_0 = block_addr_matches_14_0 & lcam_addr_0[5:3] == ldq_14_bits_addr_bits[5:3];
  wire        dword_addr_matches_14_1 = block_addr_matches_14_1 & lcam_addr_1[5:3] == ldq_14_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_56 = casez_tmp_405 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_58 = casez_tmp_405 & casez_tmp_388;
  wire        _GEN_666 = fired_release_0 & ldq_14_valid & ldq_14_bits_addr_valid & block_addr_matches_14_0;
  wire        _GEN_667 = ldq_14_bits_executed | ldq_14_bits_succeeded;
  wire        _GEN_668 = _GEN_667 | l_is_forwarding_14;
  wire [31:0] _GEN_669 = ldq_14_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_670 = do_st_search_0 & ldq_14_valid & ldq_14_bits_addr_valid & _GEN_668 & ~ldq_14_bits_addr_is_virtual & _GEN_669[0] & dword_addr_matches_14_0 & (|_mask_overlap_T_56);
  wire        _GEN_671 = ~ldq_14_bits_forward_std_val | l_forward_stq_idx_14 != lcam_stq_idx_0 & (l_forward_stq_idx_14 < lcam_stq_idx_0 ^ l_forward_stq_idx_14 < ldq_14_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_14_bits_youngest_stq_idx);
  wire        _GEN_672 = do_ld_search_0 & ldq_14_valid & ldq_14_bits_addr_valid & ~ldq_14_bits_addr_is_virtual & dword_addr_matches_14_0 & (|_mask_overlap_T_56);
  wire        searcher_is_older_28 = lcam_ldq_idx_0 < 5'hE ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'hE;
  wire        _GEN_673 = _GEN_668 & ~s1_executing_loads_14 & ldq_14_bits_observed;
  wire        _GEN_674 = ~_GEN_666 & (_GEN_670 ? _GEN_671 : _GEN_672 & searcher_is_older_28 & _GEN_673);
  reg         older_nacked_REG_28;
  wire        _GEN_675 = ~_GEN_667 | nacking_loads_14 | older_nacked_REG_28;
  wire        _GEN_676 = searcher_is_older_28 | _GEN_309;
  wire        _GEN_677 = _GEN_666 | _GEN_670;
  reg         io_dmem_s1_kill_0_REG_14;
  wire        _GEN_678 = _GEN_677 | ~_GEN_672 | _GEN_676 | ~_GEN_675;
  wire        _GEN_679 = fired_release_1 & ldq_14_valid & ldq_14_bits_addr_valid & block_addr_matches_14_1;
  wire [31:0] _GEN_680 = ldq_14_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_681 = do_st_search_1 & ldq_14_valid & ldq_14_bits_addr_valid & _GEN_668 & ~ldq_14_bits_addr_is_virtual & _GEN_680[0] & dword_addr_matches_14_1 & (|_mask_overlap_T_58);
  wire        _GEN_682 = ~ldq_14_bits_forward_std_val | l_forward_stq_idx_14 != lcam_stq_idx_1 & (l_forward_stq_idx_14 < lcam_stq_idx_1 ^ l_forward_stq_idx_14 < ldq_14_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_14_bits_youngest_stq_idx);
  wire        _GEN_683 = do_ld_search_1 & ldq_14_valid & ldq_14_bits_addr_valid & ~ldq_14_bits_addr_is_virtual & dword_addr_matches_14_1 & (|_mask_overlap_T_58);
  wire        searcher_is_older_29 = lcam_ldq_idx_1 < 5'hE ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'hE;
  wire        _GEN_684 = _GEN_683 & searcher_is_older_29 & _GEN_673;
  wire        _temp_bits_WIRE_1_46 = _GEN_679 ? _GEN_674 : _GEN_681 ? _GEN_682 | _GEN_674 : _GEN_684 | _GEN_674;
  reg         older_nacked_REG_29;
  wire        _GEN_685 = ~_GEN_667 | nacking_loads_14 | older_nacked_REG_29;
  wire        _GEN_686 = searcher_is_older_29 | _GEN_349;
  wire        _GEN_687 = _GEN_679 | _GEN_681;
  reg         io_dmem_s1_kill_1_REG_14;
  wire        _GEN_688 = _GEN_687 | ~_GEN_683 | _GEN_686 | ~_GEN_685;
  reg  [7:0]  casez_tmp_406;
  wire [14:0] _l_mask_mask_T_227 = 15'h1 << ldq_15_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_231 = 15'h3 << {12'h0, ldq_15_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_15_bits_uop_mem_size)
      2'b00:
        casez_tmp_406 = _l_mask_mask_T_227[7:0];
      2'b01:
        casez_tmp_406 = _l_mask_mask_T_231[7:0];
      2'b10:
        casez_tmp_406 = ldq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_406 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_15_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hF;
  wire        l_forwarders_15_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hF;
  wire        l_is_forwarding_15 = l_forwarders_15_0 | l_forwarders_15_1;
  wire [4:0]  l_forward_stq_idx_15 = l_is_forwarding_15 ? (l_forwarders_15_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_15_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_15_bits_forward_stq_idx;
  wire        block_addr_matches_15_0 = lcam_addr_0[39:6] == ldq_15_bits_addr_bits[39:6];
  wire        block_addr_matches_15_1 = lcam_addr_1[39:6] == ldq_15_bits_addr_bits[39:6];
  wire        dword_addr_matches_15_0 = block_addr_matches_15_0 & lcam_addr_0[5:3] == ldq_15_bits_addr_bits[5:3];
  wire        dword_addr_matches_15_1 = block_addr_matches_15_1 & lcam_addr_1[5:3] == ldq_15_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_60 = casez_tmp_406 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_62 = casez_tmp_406 & casez_tmp_388;
  wire        _GEN_689 = fired_release_0 & ldq_15_valid & ldq_15_bits_addr_valid & block_addr_matches_15_0;
  wire        _GEN_690 = ldq_15_bits_executed | ldq_15_bits_succeeded;
  wire        _GEN_691 = _GEN_690 | l_is_forwarding_15;
  wire [31:0] _GEN_692 = ldq_15_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_693 = do_st_search_0 & ldq_15_valid & ldq_15_bits_addr_valid & _GEN_691 & ~ldq_15_bits_addr_is_virtual & _GEN_692[0] & dword_addr_matches_15_0 & (|_mask_overlap_T_60);
  wire        _GEN_694 = ~ldq_15_bits_forward_std_val | l_forward_stq_idx_15 != lcam_stq_idx_0 & (l_forward_stq_idx_15 < lcam_stq_idx_0 ^ l_forward_stq_idx_15 < ldq_15_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_15_bits_youngest_stq_idx);
  wire        _GEN_695 = do_ld_search_0 & ldq_15_valid & ldq_15_bits_addr_valid & ~ldq_15_bits_addr_is_virtual & dword_addr_matches_15_0 & (|_mask_overlap_T_60);
  wire        searcher_is_older_30 = lcam_ldq_idx_0 < 5'hF ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head[4];
  wire        _GEN_696 = _GEN_691 & ~s1_executing_loads_15 & ldq_15_bits_observed;
  wire        _GEN_697 = ~_GEN_689 & (_GEN_693 ? _GEN_694 : _GEN_695 & searcher_is_older_30 & _GEN_696);
  reg         older_nacked_REG_30;
  wire        _GEN_698 = ~_GEN_690 | nacking_loads_15 | older_nacked_REG_30;
  wire        _GEN_699 = searcher_is_older_30 | _GEN_310;
  wire        _GEN_700 = _GEN_689 | _GEN_693;
  reg         io_dmem_s1_kill_0_REG_15;
  wire        _GEN_701 = _GEN_700 | ~_GEN_695 | _GEN_699 | ~_GEN_698;
  wire        _GEN_702 = fired_release_1 & ldq_15_valid & ldq_15_bits_addr_valid & block_addr_matches_15_1;
  wire [31:0] _GEN_703 = ldq_15_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_704 = do_st_search_1 & ldq_15_valid & ldq_15_bits_addr_valid & _GEN_691 & ~ldq_15_bits_addr_is_virtual & _GEN_703[0] & dword_addr_matches_15_1 & (|_mask_overlap_T_62);
  wire        _GEN_705 = ~ldq_15_bits_forward_std_val | l_forward_stq_idx_15 != lcam_stq_idx_1 & (l_forward_stq_idx_15 < lcam_stq_idx_1 ^ l_forward_stq_idx_15 < ldq_15_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_15_bits_youngest_stq_idx);
  wire        _GEN_706 = do_ld_search_1 & ldq_15_valid & ldq_15_bits_addr_valid & ~ldq_15_bits_addr_is_virtual & dword_addr_matches_15_1 & (|_mask_overlap_T_62);
  wire        searcher_is_older_31 = lcam_ldq_idx_1 < 5'hF ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head[4];
  wire        _GEN_707 = _GEN_706 & searcher_is_older_31 & _GEN_696;
  wire        _temp_bits_WIRE_1_47 = _GEN_702 ? _GEN_697 : _GEN_704 ? _GEN_705 | _GEN_697 : _GEN_707 | _GEN_697;
  reg         older_nacked_REG_31;
  wire        _GEN_708 = ~_GEN_690 | nacking_loads_15 | older_nacked_REG_31;
  wire        _GEN_709 = searcher_is_older_31 | _GEN_350;
  wire        _GEN_710 = _GEN_702 | _GEN_704;
  reg         io_dmem_s1_kill_1_REG_15;
  wire        _GEN_711 = _GEN_710 | ~_GEN_706 | _GEN_709 | ~_GEN_708;
  reg  [7:0]  casez_tmp_407;
  wire [14:0] _l_mask_mask_T_242 = 15'h1 << ldq_16_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_246 = 15'h3 << {12'h0, ldq_16_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_16_bits_uop_mem_size)
      2'b00:
        casez_tmp_407 = _l_mask_mask_T_242[7:0];
      2'b01:
        casez_tmp_407 = _l_mask_mask_T_246[7:0];
      2'b10:
        casez_tmp_407 = ldq_16_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_407 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_16_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h10;
  wire        l_forwarders_16_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h10;
  wire        l_is_forwarding_16 = l_forwarders_16_0 | l_forwarders_16_1;
  wire [4:0]  l_forward_stq_idx_16 = l_is_forwarding_16 ? (l_forwarders_16_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_16_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_16_bits_forward_stq_idx;
  wire        block_addr_matches_16_0 = lcam_addr_0[39:6] == ldq_16_bits_addr_bits[39:6];
  wire        block_addr_matches_16_1 = lcam_addr_1[39:6] == ldq_16_bits_addr_bits[39:6];
  wire        dword_addr_matches_16_0 = block_addr_matches_16_0 & lcam_addr_0[5:3] == ldq_16_bits_addr_bits[5:3];
  wire        dword_addr_matches_16_1 = block_addr_matches_16_1 & lcam_addr_1[5:3] == ldq_16_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_64 = casez_tmp_407 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_66 = casez_tmp_407 & casez_tmp_388;
  wire        _GEN_712 = fired_release_0 & ldq_16_valid & ldq_16_bits_addr_valid & block_addr_matches_16_0;
  wire        _GEN_713 = ldq_16_bits_executed | ldq_16_bits_succeeded;
  wire        _GEN_714 = _GEN_713 | l_is_forwarding_16;
  wire [31:0] _GEN_715 = ldq_16_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_716 = do_st_search_0 & ldq_16_valid & ldq_16_bits_addr_valid & _GEN_714 & ~ldq_16_bits_addr_is_virtual & _GEN_715[0] & dword_addr_matches_16_0 & (|_mask_overlap_T_64);
  wire        _GEN_717 = ~ldq_16_bits_forward_std_val | l_forward_stq_idx_16 != lcam_stq_idx_0 & (l_forward_stq_idx_16 < lcam_stq_idx_0 ^ l_forward_stq_idx_16 < ldq_16_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_16_bits_youngest_stq_idx);
  wire        _GEN_718 = do_ld_search_0 & ldq_16_valid & ldq_16_bits_addr_valid & ~ldq_16_bits_addr_is_virtual & dword_addr_matches_16_0 & (|_mask_overlap_T_64);
  wire        searcher_is_older_32 = lcam_ldq_idx_0[4] ^ lcam_ldq_idx_0 >= ldq_head ^ ldq_head > 5'h10;
  wire        _GEN_719 = _GEN_714 & ~s1_executing_loads_16 & ldq_16_bits_observed;
  wire        _GEN_720 = ~_GEN_712 & (_GEN_716 ? _GEN_717 : _GEN_718 & searcher_is_older_32 & _GEN_719);
  reg         older_nacked_REG_32;
  wire        _GEN_721 = ~_GEN_713 | nacking_loads_16 | older_nacked_REG_32;
  wire        _GEN_722 = searcher_is_older_32 | _GEN_311;
  wire        _GEN_723 = _GEN_712 | _GEN_716;
  reg         io_dmem_s1_kill_0_REG_16;
  wire        _GEN_724 = _GEN_723 | ~_GEN_718 | _GEN_722 | ~_GEN_721;
  wire        _GEN_725 = fired_release_1 & ldq_16_valid & ldq_16_bits_addr_valid & block_addr_matches_16_1;
  wire [31:0] _GEN_726 = ldq_16_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_727 = do_st_search_1 & ldq_16_valid & ldq_16_bits_addr_valid & _GEN_714 & ~ldq_16_bits_addr_is_virtual & _GEN_726[0] & dword_addr_matches_16_1 & (|_mask_overlap_T_66);
  wire        _GEN_728 = ~ldq_16_bits_forward_std_val | l_forward_stq_idx_16 != lcam_stq_idx_1 & (l_forward_stq_idx_16 < lcam_stq_idx_1 ^ l_forward_stq_idx_16 < ldq_16_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_16_bits_youngest_stq_idx);
  wire        _GEN_729 = do_ld_search_1 & ldq_16_valid & ldq_16_bits_addr_valid & ~ldq_16_bits_addr_is_virtual & dword_addr_matches_16_1 & (|_mask_overlap_T_66);
  wire        searcher_is_older_33 = lcam_ldq_idx_1[4] ^ lcam_ldq_idx_1 >= ldq_head ^ ldq_head > 5'h10;
  wire        _GEN_730 = _GEN_729 & searcher_is_older_33 & _GEN_719;
  wire        _temp_bits_WIRE_1_48 = _GEN_725 ? _GEN_720 : _GEN_727 ? _GEN_728 | _GEN_720 : _GEN_730 | _GEN_720;
  reg         older_nacked_REG_33;
  wire        _GEN_731 = ~_GEN_713 | nacking_loads_16 | older_nacked_REG_33;
  wire        _GEN_732 = searcher_is_older_33 | _GEN_351;
  wire        _GEN_733 = _GEN_725 | _GEN_727;
  reg         io_dmem_s1_kill_1_REG_16;
  wire        _GEN_734 = _GEN_733 | ~_GEN_729 | _GEN_732 | ~_GEN_731;
  reg  [7:0]  casez_tmp_408;
  wire [14:0] _l_mask_mask_T_257 = 15'h1 << ldq_17_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_261 = 15'h3 << {12'h0, ldq_17_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_17_bits_uop_mem_size)
      2'b00:
        casez_tmp_408 = _l_mask_mask_T_257[7:0];
      2'b01:
        casez_tmp_408 = _l_mask_mask_T_261[7:0];
      2'b10:
        casez_tmp_408 = ldq_17_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_408 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_17_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h11;
  wire        l_forwarders_17_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h11;
  wire        l_is_forwarding_17 = l_forwarders_17_0 | l_forwarders_17_1;
  wire [4:0]  l_forward_stq_idx_17 = l_is_forwarding_17 ? (l_forwarders_17_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_17_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_17_bits_forward_stq_idx;
  wire        block_addr_matches_17_0 = lcam_addr_0[39:6] == ldq_17_bits_addr_bits[39:6];
  wire        block_addr_matches_17_1 = lcam_addr_1[39:6] == ldq_17_bits_addr_bits[39:6];
  wire        dword_addr_matches_17_0 = block_addr_matches_17_0 & lcam_addr_0[5:3] == ldq_17_bits_addr_bits[5:3];
  wire        dword_addr_matches_17_1 = block_addr_matches_17_1 & lcam_addr_1[5:3] == ldq_17_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_68 = casez_tmp_408 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_70 = casez_tmp_408 & casez_tmp_388;
  wire        _GEN_735 = fired_release_0 & ldq_17_valid & ldq_17_bits_addr_valid & block_addr_matches_17_0;
  wire        _GEN_736 = ldq_17_bits_executed | ldq_17_bits_succeeded;
  wire        _GEN_737 = _GEN_736 | l_is_forwarding_17;
  wire [31:0] _GEN_738 = ldq_17_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_739 = do_st_search_0 & ldq_17_valid & ldq_17_bits_addr_valid & _GEN_737 & ~ldq_17_bits_addr_is_virtual & _GEN_738[0] & dword_addr_matches_17_0 & (|_mask_overlap_T_68);
  wire        _GEN_740 = ~ldq_17_bits_forward_std_val | l_forward_stq_idx_17 != lcam_stq_idx_0 & (l_forward_stq_idx_17 < lcam_stq_idx_0 ^ l_forward_stq_idx_17 < ldq_17_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_17_bits_youngest_stq_idx);
  wire        _GEN_741 = do_ld_search_0 & ldq_17_valid & ldq_17_bits_addr_valid & ~ldq_17_bits_addr_is_virtual & dword_addr_matches_17_0 & (|_mask_overlap_T_68);
  wire        searcher_is_older_34 = lcam_ldq_idx_0 < 5'h11 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h11;
  wire        _GEN_742 = _GEN_737 & ~s1_executing_loads_17 & ldq_17_bits_observed;
  wire        _GEN_743 = ~_GEN_735 & (_GEN_739 ? _GEN_740 : _GEN_741 & searcher_is_older_34 & _GEN_742);
  reg         older_nacked_REG_34;
  wire        _GEN_744 = ~_GEN_736 | nacking_loads_17 | older_nacked_REG_34;
  wire        _GEN_745 = searcher_is_older_34 | _GEN_312;
  wire        _GEN_746 = _GEN_735 | _GEN_739;
  reg         io_dmem_s1_kill_0_REG_17;
  wire        _GEN_747 = _GEN_746 | ~_GEN_741 | _GEN_745 | ~_GEN_744;
  wire        _GEN_748 = fired_release_1 & ldq_17_valid & ldq_17_bits_addr_valid & block_addr_matches_17_1;
  wire [31:0] _GEN_749 = ldq_17_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_750 = do_st_search_1 & ldq_17_valid & ldq_17_bits_addr_valid & _GEN_737 & ~ldq_17_bits_addr_is_virtual & _GEN_749[0] & dword_addr_matches_17_1 & (|_mask_overlap_T_70);
  wire        _GEN_751 = ~ldq_17_bits_forward_std_val | l_forward_stq_idx_17 != lcam_stq_idx_1 & (l_forward_stq_idx_17 < lcam_stq_idx_1 ^ l_forward_stq_idx_17 < ldq_17_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_17_bits_youngest_stq_idx);
  wire        _GEN_752 = do_ld_search_1 & ldq_17_valid & ldq_17_bits_addr_valid & ~ldq_17_bits_addr_is_virtual & dword_addr_matches_17_1 & (|_mask_overlap_T_70);
  wire        searcher_is_older_35 = lcam_ldq_idx_1 < 5'h11 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h11;
  wire        _GEN_753 = _GEN_752 & searcher_is_older_35 & _GEN_742;
  wire        _temp_bits_WIRE_1_49 = _GEN_748 ? _GEN_743 : _GEN_750 ? _GEN_751 | _GEN_743 : _GEN_753 | _GEN_743;
  reg         older_nacked_REG_35;
  wire        _GEN_754 = ~_GEN_736 | nacking_loads_17 | older_nacked_REG_35;
  wire        _GEN_755 = searcher_is_older_35 | _GEN_352;
  wire        _GEN_756 = _GEN_748 | _GEN_750;
  reg         io_dmem_s1_kill_1_REG_17;
  wire        _GEN_757 = _GEN_756 | ~_GEN_752 | _GEN_755 | ~_GEN_754;
  reg  [7:0]  casez_tmp_409;
  wire [14:0] _l_mask_mask_T_272 = 15'h1 << ldq_18_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_276 = 15'h3 << {12'h0, ldq_18_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_18_bits_uop_mem_size)
      2'b00:
        casez_tmp_409 = _l_mask_mask_T_272[7:0];
      2'b01:
        casez_tmp_409 = _l_mask_mask_T_276[7:0];
      2'b10:
        casez_tmp_409 = ldq_18_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_409 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_18_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h12;
  wire        l_forwarders_18_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h12;
  wire        l_is_forwarding_18 = l_forwarders_18_0 | l_forwarders_18_1;
  wire [4:0]  l_forward_stq_idx_18 = l_is_forwarding_18 ? (l_forwarders_18_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_18_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_18_bits_forward_stq_idx;
  wire        block_addr_matches_18_0 = lcam_addr_0[39:6] == ldq_18_bits_addr_bits[39:6];
  wire        block_addr_matches_18_1 = lcam_addr_1[39:6] == ldq_18_bits_addr_bits[39:6];
  wire        dword_addr_matches_18_0 = block_addr_matches_18_0 & lcam_addr_0[5:3] == ldq_18_bits_addr_bits[5:3];
  wire        dword_addr_matches_18_1 = block_addr_matches_18_1 & lcam_addr_1[5:3] == ldq_18_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_72 = casez_tmp_409 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_74 = casez_tmp_409 & casez_tmp_388;
  wire        _GEN_758 = fired_release_0 & ldq_18_valid & ldq_18_bits_addr_valid & block_addr_matches_18_0;
  wire        _GEN_759 = ldq_18_bits_executed | ldq_18_bits_succeeded;
  wire        _GEN_760 = _GEN_759 | l_is_forwarding_18;
  wire [31:0] _GEN_761 = ldq_18_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_762 = do_st_search_0 & ldq_18_valid & ldq_18_bits_addr_valid & _GEN_760 & ~ldq_18_bits_addr_is_virtual & _GEN_761[0] & dword_addr_matches_18_0 & (|_mask_overlap_T_72);
  wire        _GEN_763 = ~ldq_18_bits_forward_std_val | l_forward_stq_idx_18 != lcam_stq_idx_0 & (l_forward_stq_idx_18 < lcam_stq_idx_0 ^ l_forward_stq_idx_18 < ldq_18_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_18_bits_youngest_stq_idx);
  wire        _GEN_764 = do_ld_search_0 & ldq_18_valid & ldq_18_bits_addr_valid & ~ldq_18_bits_addr_is_virtual & dword_addr_matches_18_0 & (|_mask_overlap_T_72);
  wire        searcher_is_older_36 = lcam_ldq_idx_0 < 5'h12 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h12;
  wire        _GEN_765 = _GEN_760 & ~s1_executing_loads_18 & ldq_18_bits_observed;
  wire        _GEN_766 = ~_GEN_758 & (_GEN_762 ? _GEN_763 : _GEN_764 & searcher_is_older_36 & _GEN_765);
  reg         older_nacked_REG_36;
  wire        _GEN_767 = ~_GEN_759 | nacking_loads_18 | older_nacked_REG_36;
  wire        _GEN_768 = searcher_is_older_36 | _GEN_313;
  wire        _GEN_769 = _GEN_758 | _GEN_762;
  reg         io_dmem_s1_kill_0_REG_18;
  wire        _GEN_770 = _GEN_769 | ~_GEN_764 | _GEN_768 | ~_GEN_767;
  wire        _GEN_771 = fired_release_1 & ldq_18_valid & ldq_18_bits_addr_valid & block_addr_matches_18_1;
  wire [31:0] _GEN_772 = ldq_18_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_773 = do_st_search_1 & ldq_18_valid & ldq_18_bits_addr_valid & _GEN_760 & ~ldq_18_bits_addr_is_virtual & _GEN_772[0] & dword_addr_matches_18_1 & (|_mask_overlap_T_74);
  wire        _GEN_774 = ~ldq_18_bits_forward_std_val | l_forward_stq_idx_18 != lcam_stq_idx_1 & (l_forward_stq_idx_18 < lcam_stq_idx_1 ^ l_forward_stq_idx_18 < ldq_18_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_18_bits_youngest_stq_idx);
  wire        _GEN_775 = do_ld_search_1 & ldq_18_valid & ldq_18_bits_addr_valid & ~ldq_18_bits_addr_is_virtual & dword_addr_matches_18_1 & (|_mask_overlap_T_74);
  wire        searcher_is_older_37 = lcam_ldq_idx_1 < 5'h12 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h12;
  wire        _GEN_776 = _GEN_775 & searcher_is_older_37 & _GEN_765;
  wire        _temp_bits_WIRE_1_50 = _GEN_771 ? _GEN_766 : _GEN_773 ? _GEN_774 | _GEN_766 : _GEN_776 | _GEN_766;
  reg         older_nacked_REG_37;
  wire        _GEN_777 = ~_GEN_759 | nacking_loads_18 | older_nacked_REG_37;
  wire        _GEN_778 = searcher_is_older_37 | _GEN_353;
  wire        _GEN_779 = _GEN_771 | _GEN_773;
  reg         io_dmem_s1_kill_1_REG_18;
  wire        _GEN_780 = _GEN_779 | ~_GEN_775 | _GEN_778 | ~_GEN_777;
  reg  [7:0]  casez_tmp_410;
  wire [14:0] _l_mask_mask_T_287 = 15'h1 << ldq_19_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_291 = 15'h3 << {12'h0, ldq_19_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_19_bits_uop_mem_size)
      2'b00:
        casez_tmp_410 = _l_mask_mask_T_287[7:0];
      2'b01:
        casez_tmp_410 = _l_mask_mask_T_291[7:0];
      2'b10:
        casez_tmp_410 = ldq_19_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_410 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_19_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h13;
  wire        l_forwarders_19_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h13;
  wire        l_is_forwarding_19 = l_forwarders_19_0 | l_forwarders_19_1;
  wire [4:0]  l_forward_stq_idx_19 = l_is_forwarding_19 ? (l_forwarders_19_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_19_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_19_bits_forward_stq_idx;
  wire        block_addr_matches_19_0 = lcam_addr_0[39:6] == ldq_19_bits_addr_bits[39:6];
  wire        block_addr_matches_19_1 = lcam_addr_1[39:6] == ldq_19_bits_addr_bits[39:6];
  wire        dword_addr_matches_19_0 = block_addr_matches_19_0 & lcam_addr_0[5:3] == ldq_19_bits_addr_bits[5:3];
  wire        dword_addr_matches_19_1 = block_addr_matches_19_1 & lcam_addr_1[5:3] == ldq_19_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_76 = casez_tmp_410 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_78 = casez_tmp_410 & casez_tmp_388;
  wire        _GEN_781 = fired_release_0 & ldq_19_valid & ldq_19_bits_addr_valid & block_addr_matches_19_0;
  wire        _GEN_782 = ldq_19_bits_executed | ldq_19_bits_succeeded;
  wire        _GEN_783 = _GEN_782 | l_is_forwarding_19;
  wire [31:0] _GEN_784 = ldq_19_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_785 = do_st_search_0 & ldq_19_valid & ldq_19_bits_addr_valid & _GEN_783 & ~ldq_19_bits_addr_is_virtual & _GEN_784[0] & dword_addr_matches_19_0 & (|_mask_overlap_T_76);
  wire        _GEN_786 = ~ldq_19_bits_forward_std_val | l_forward_stq_idx_19 != lcam_stq_idx_0 & (l_forward_stq_idx_19 < lcam_stq_idx_0 ^ l_forward_stq_idx_19 < ldq_19_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_19_bits_youngest_stq_idx);
  wire        _GEN_787 = do_ld_search_0 & ldq_19_valid & ldq_19_bits_addr_valid & ~ldq_19_bits_addr_is_virtual & dword_addr_matches_19_0 & (|_mask_overlap_T_76);
  wire        searcher_is_older_38 = lcam_ldq_idx_0 < 5'h13 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h13;
  wire        _GEN_788 = _GEN_783 & ~s1_executing_loads_19 & ldq_19_bits_observed;
  wire        _GEN_789 = ~_GEN_781 & (_GEN_785 ? _GEN_786 : _GEN_787 & searcher_is_older_38 & _GEN_788);
  reg         older_nacked_REG_38;
  wire        _GEN_790 = ~_GEN_782 | nacking_loads_19 | older_nacked_REG_38;
  wire        _GEN_791 = searcher_is_older_38 | _GEN_314;
  wire        _GEN_792 = _GEN_781 | _GEN_785;
  reg         io_dmem_s1_kill_0_REG_19;
  wire        _GEN_793 = _GEN_792 | ~_GEN_787 | _GEN_791 | ~_GEN_790;
  wire        _GEN_794 = fired_release_1 & ldq_19_valid & ldq_19_bits_addr_valid & block_addr_matches_19_1;
  wire [31:0] _GEN_795 = ldq_19_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_796 = do_st_search_1 & ldq_19_valid & ldq_19_bits_addr_valid & _GEN_783 & ~ldq_19_bits_addr_is_virtual & _GEN_795[0] & dword_addr_matches_19_1 & (|_mask_overlap_T_78);
  wire        _GEN_797 = ~ldq_19_bits_forward_std_val | l_forward_stq_idx_19 != lcam_stq_idx_1 & (l_forward_stq_idx_19 < lcam_stq_idx_1 ^ l_forward_stq_idx_19 < ldq_19_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_19_bits_youngest_stq_idx);
  wire        _GEN_798 = do_ld_search_1 & ldq_19_valid & ldq_19_bits_addr_valid & ~ldq_19_bits_addr_is_virtual & dword_addr_matches_19_1 & (|_mask_overlap_T_78);
  wire        searcher_is_older_39 = lcam_ldq_idx_1 < 5'h13 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h13;
  wire        _GEN_799 = _GEN_798 & searcher_is_older_39 & _GEN_788;
  wire        _temp_bits_WIRE_1_51 = _GEN_794 ? _GEN_789 : _GEN_796 ? _GEN_797 | _GEN_789 : _GEN_799 | _GEN_789;
  reg         older_nacked_REG_39;
  wire        _GEN_800 = ~_GEN_782 | nacking_loads_19 | older_nacked_REG_39;
  wire        _GEN_801 = searcher_is_older_39 | _GEN_354;
  wire        _GEN_802 = _GEN_794 | _GEN_796;
  reg         io_dmem_s1_kill_1_REG_19;
  wire        _GEN_803 = _GEN_802 | ~_GEN_798 | _GEN_801 | ~_GEN_800;
  reg  [7:0]  casez_tmp_411;
  wire [14:0] _l_mask_mask_T_302 = 15'h1 << ldq_20_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_306 = 15'h3 << {12'h0, ldq_20_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_20_bits_uop_mem_size)
      2'b00:
        casez_tmp_411 = _l_mask_mask_T_302[7:0];
      2'b01:
        casez_tmp_411 = _l_mask_mask_T_306[7:0];
      2'b10:
        casez_tmp_411 = ldq_20_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_411 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_20_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h14;
  wire        l_forwarders_20_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h14;
  wire        l_is_forwarding_20 = l_forwarders_20_0 | l_forwarders_20_1;
  wire [4:0]  l_forward_stq_idx_20 = l_is_forwarding_20 ? (l_forwarders_20_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_20_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_20_bits_forward_stq_idx;
  wire        block_addr_matches_20_0 = lcam_addr_0[39:6] == ldq_20_bits_addr_bits[39:6];
  wire        block_addr_matches_20_1 = lcam_addr_1[39:6] == ldq_20_bits_addr_bits[39:6];
  wire        dword_addr_matches_20_0 = block_addr_matches_20_0 & lcam_addr_0[5:3] == ldq_20_bits_addr_bits[5:3];
  wire        dword_addr_matches_20_1 = block_addr_matches_20_1 & lcam_addr_1[5:3] == ldq_20_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_80 = casez_tmp_411 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_82 = casez_tmp_411 & casez_tmp_388;
  wire        _GEN_804 = fired_release_0 & ldq_20_valid & ldq_20_bits_addr_valid & block_addr_matches_20_0;
  wire        _GEN_805 = ldq_20_bits_executed | ldq_20_bits_succeeded;
  wire        _GEN_806 = _GEN_805 | l_is_forwarding_20;
  wire [31:0] _GEN_807 = ldq_20_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_808 = do_st_search_0 & ldq_20_valid & ldq_20_bits_addr_valid & _GEN_806 & ~ldq_20_bits_addr_is_virtual & _GEN_807[0] & dword_addr_matches_20_0 & (|_mask_overlap_T_80);
  wire        _GEN_809 = ~ldq_20_bits_forward_std_val | l_forward_stq_idx_20 != lcam_stq_idx_0 & (l_forward_stq_idx_20 < lcam_stq_idx_0 ^ l_forward_stq_idx_20 < ldq_20_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_20_bits_youngest_stq_idx);
  wire        _GEN_810 = do_ld_search_0 & ldq_20_valid & ldq_20_bits_addr_valid & ~ldq_20_bits_addr_is_virtual & dword_addr_matches_20_0 & (|_mask_overlap_T_80);
  wire        searcher_is_older_40 = lcam_ldq_idx_0 < 5'h14 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h14;
  wire        _GEN_811 = _GEN_806 & ~s1_executing_loads_20 & ldq_20_bits_observed;
  wire        _GEN_812 = ~_GEN_804 & (_GEN_808 ? _GEN_809 : _GEN_810 & searcher_is_older_40 & _GEN_811);
  reg         older_nacked_REG_40;
  wire        _GEN_813 = ~_GEN_805 | nacking_loads_20 | older_nacked_REG_40;
  wire        _GEN_814 = searcher_is_older_40 | _GEN_315;
  wire        _GEN_815 = _GEN_804 | _GEN_808;
  reg         io_dmem_s1_kill_0_REG_20;
  wire        _GEN_816 = _GEN_815 | ~_GEN_810 | _GEN_814 | ~_GEN_813;
  wire        _GEN_817 = fired_release_1 & ldq_20_valid & ldq_20_bits_addr_valid & block_addr_matches_20_1;
  wire [31:0] _GEN_818 = ldq_20_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_819 = do_st_search_1 & ldq_20_valid & ldq_20_bits_addr_valid & _GEN_806 & ~ldq_20_bits_addr_is_virtual & _GEN_818[0] & dword_addr_matches_20_1 & (|_mask_overlap_T_82);
  wire        _GEN_820 = ~ldq_20_bits_forward_std_val | l_forward_stq_idx_20 != lcam_stq_idx_1 & (l_forward_stq_idx_20 < lcam_stq_idx_1 ^ l_forward_stq_idx_20 < ldq_20_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_20_bits_youngest_stq_idx);
  wire        _GEN_821 = do_ld_search_1 & ldq_20_valid & ldq_20_bits_addr_valid & ~ldq_20_bits_addr_is_virtual & dword_addr_matches_20_1 & (|_mask_overlap_T_82);
  wire        searcher_is_older_41 = lcam_ldq_idx_1 < 5'h14 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h14;
  wire        _GEN_822 = _GEN_821 & searcher_is_older_41 & _GEN_811;
  wire        _temp_bits_WIRE_1_52 = _GEN_817 ? _GEN_812 : _GEN_819 ? _GEN_820 | _GEN_812 : _GEN_822 | _GEN_812;
  reg         older_nacked_REG_41;
  wire        _GEN_823 = ~_GEN_805 | nacking_loads_20 | older_nacked_REG_41;
  wire        _GEN_824 = searcher_is_older_41 | _GEN_355;
  wire        _GEN_825 = _GEN_817 | _GEN_819;
  reg         io_dmem_s1_kill_1_REG_20;
  wire        _GEN_826 = _GEN_825 | ~_GEN_821 | _GEN_824 | ~_GEN_823;
  reg  [7:0]  casez_tmp_412;
  wire [14:0] _l_mask_mask_T_317 = 15'h1 << ldq_21_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_321 = 15'h3 << {12'h0, ldq_21_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_21_bits_uop_mem_size)
      2'b00:
        casez_tmp_412 = _l_mask_mask_T_317[7:0];
      2'b01:
        casez_tmp_412 = _l_mask_mask_T_321[7:0];
      2'b10:
        casez_tmp_412 = ldq_21_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_412 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_21_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h15;
  wire        l_forwarders_21_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h15;
  wire        l_is_forwarding_21 = l_forwarders_21_0 | l_forwarders_21_1;
  wire [4:0]  l_forward_stq_idx_21 = l_is_forwarding_21 ? (l_forwarders_21_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_21_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_21_bits_forward_stq_idx;
  wire        block_addr_matches_21_0 = lcam_addr_0[39:6] == ldq_21_bits_addr_bits[39:6];
  wire        block_addr_matches_21_1 = lcam_addr_1[39:6] == ldq_21_bits_addr_bits[39:6];
  wire        dword_addr_matches_21_0 = block_addr_matches_21_0 & lcam_addr_0[5:3] == ldq_21_bits_addr_bits[5:3];
  wire        dword_addr_matches_21_1 = block_addr_matches_21_1 & lcam_addr_1[5:3] == ldq_21_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_84 = casez_tmp_412 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_86 = casez_tmp_412 & casez_tmp_388;
  wire        _GEN_827 = fired_release_0 & ldq_21_valid & ldq_21_bits_addr_valid & block_addr_matches_21_0;
  wire        _GEN_828 = ldq_21_bits_executed | ldq_21_bits_succeeded;
  wire        _GEN_829 = _GEN_828 | l_is_forwarding_21;
  wire [31:0] _GEN_830 = ldq_21_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_831 = do_st_search_0 & ldq_21_valid & ldq_21_bits_addr_valid & _GEN_829 & ~ldq_21_bits_addr_is_virtual & _GEN_830[0] & dword_addr_matches_21_0 & (|_mask_overlap_T_84);
  wire        _GEN_832 = ~ldq_21_bits_forward_std_val | l_forward_stq_idx_21 != lcam_stq_idx_0 & (l_forward_stq_idx_21 < lcam_stq_idx_0 ^ l_forward_stq_idx_21 < ldq_21_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_21_bits_youngest_stq_idx);
  wire        _GEN_833 = do_ld_search_0 & ldq_21_valid & ldq_21_bits_addr_valid & ~ldq_21_bits_addr_is_virtual & dword_addr_matches_21_0 & (|_mask_overlap_T_84);
  wire        searcher_is_older_42 = lcam_ldq_idx_0 < 5'h15 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h15;
  wire        _GEN_834 = _GEN_829 & ~s1_executing_loads_21 & ldq_21_bits_observed;
  wire        _GEN_835 = ~_GEN_827 & (_GEN_831 ? _GEN_832 : _GEN_833 & searcher_is_older_42 & _GEN_834);
  reg         older_nacked_REG_42;
  wire        _GEN_836 = ~_GEN_828 | nacking_loads_21 | older_nacked_REG_42;
  wire        _GEN_837 = searcher_is_older_42 | _GEN_316;
  wire        _GEN_838 = _GEN_827 | _GEN_831;
  reg         io_dmem_s1_kill_0_REG_21;
  wire        _GEN_839 = _GEN_838 | ~_GEN_833 | _GEN_837 | ~_GEN_836;
  wire        _GEN_840 = fired_release_1 & ldq_21_valid & ldq_21_bits_addr_valid & block_addr_matches_21_1;
  wire [31:0] _GEN_841 = ldq_21_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_842 = do_st_search_1 & ldq_21_valid & ldq_21_bits_addr_valid & _GEN_829 & ~ldq_21_bits_addr_is_virtual & _GEN_841[0] & dword_addr_matches_21_1 & (|_mask_overlap_T_86);
  wire        _GEN_843 = ~ldq_21_bits_forward_std_val | l_forward_stq_idx_21 != lcam_stq_idx_1 & (l_forward_stq_idx_21 < lcam_stq_idx_1 ^ l_forward_stq_idx_21 < ldq_21_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_21_bits_youngest_stq_idx);
  wire        _GEN_844 = do_ld_search_1 & ldq_21_valid & ldq_21_bits_addr_valid & ~ldq_21_bits_addr_is_virtual & dword_addr_matches_21_1 & (|_mask_overlap_T_86);
  wire        searcher_is_older_43 = lcam_ldq_idx_1 < 5'h15 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h15;
  wire        _GEN_845 = _GEN_844 & searcher_is_older_43 & _GEN_834;
  wire        _temp_bits_WIRE_1_53 = _GEN_840 ? _GEN_835 : _GEN_842 ? _GEN_843 | _GEN_835 : _GEN_845 | _GEN_835;
  reg         older_nacked_REG_43;
  wire        _GEN_846 = ~_GEN_828 | nacking_loads_21 | older_nacked_REG_43;
  wire        _GEN_847 = searcher_is_older_43 | _GEN_356;
  wire        _GEN_848 = _GEN_840 | _GEN_842;
  reg         io_dmem_s1_kill_1_REG_21;
  wire        _GEN_849 = _GEN_848 | ~_GEN_844 | _GEN_847 | ~_GEN_846;
  reg  [7:0]  casez_tmp_413;
  wire [14:0] _l_mask_mask_T_332 = 15'h1 << ldq_22_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_336 = 15'h3 << {12'h0, ldq_22_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_22_bits_uop_mem_size)
      2'b00:
        casez_tmp_413 = _l_mask_mask_T_332[7:0];
      2'b01:
        casez_tmp_413 = _l_mask_mask_T_336[7:0];
      2'b10:
        casez_tmp_413 = ldq_22_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_413 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_22_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h16;
  wire        l_forwarders_22_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h16;
  wire        l_is_forwarding_22 = l_forwarders_22_0 | l_forwarders_22_1;
  wire [4:0]  l_forward_stq_idx_22 = l_is_forwarding_22 ? (l_forwarders_22_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_22_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_22_bits_forward_stq_idx;
  wire        block_addr_matches_22_0 = lcam_addr_0[39:6] == ldq_22_bits_addr_bits[39:6];
  wire        block_addr_matches_22_1 = lcam_addr_1[39:6] == ldq_22_bits_addr_bits[39:6];
  wire        dword_addr_matches_22_0 = block_addr_matches_22_0 & lcam_addr_0[5:3] == ldq_22_bits_addr_bits[5:3];
  wire        dword_addr_matches_22_1 = block_addr_matches_22_1 & lcam_addr_1[5:3] == ldq_22_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_88 = casez_tmp_413 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_90 = casez_tmp_413 & casez_tmp_388;
  wire        _GEN_850 = fired_release_0 & ldq_22_valid & ldq_22_bits_addr_valid & block_addr_matches_22_0;
  wire        _GEN_851 = ldq_22_bits_executed | ldq_22_bits_succeeded;
  wire        _GEN_852 = _GEN_851 | l_is_forwarding_22;
  wire [31:0] _GEN_853 = ldq_22_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_854 = do_st_search_0 & ldq_22_valid & ldq_22_bits_addr_valid & _GEN_852 & ~ldq_22_bits_addr_is_virtual & _GEN_853[0] & dword_addr_matches_22_0 & (|_mask_overlap_T_88);
  wire        _GEN_855 = ~ldq_22_bits_forward_std_val | l_forward_stq_idx_22 != lcam_stq_idx_0 & (l_forward_stq_idx_22 < lcam_stq_idx_0 ^ l_forward_stq_idx_22 < ldq_22_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_22_bits_youngest_stq_idx);
  wire        _GEN_856 = do_ld_search_0 & ldq_22_valid & ldq_22_bits_addr_valid & ~ldq_22_bits_addr_is_virtual & dword_addr_matches_22_0 & (|_mask_overlap_T_88);
  wire        searcher_is_older_44 = lcam_ldq_idx_0 < 5'h16 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h16;
  wire        _GEN_857 = _GEN_852 & ~s1_executing_loads_22 & ldq_22_bits_observed;
  wire        _GEN_858 = ~_GEN_850 & (_GEN_854 ? _GEN_855 : _GEN_856 & searcher_is_older_44 & _GEN_857);
  reg         older_nacked_REG_44;
  wire        _GEN_859 = ~_GEN_851 | nacking_loads_22 | older_nacked_REG_44;
  wire        _GEN_860 = searcher_is_older_44 | _GEN_317;
  wire        _GEN_861 = _GEN_850 | _GEN_854;
  reg         io_dmem_s1_kill_0_REG_22;
  wire        _GEN_862 = _GEN_861 | ~_GEN_856 | _GEN_860 | ~_GEN_859;
  wire        _GEN_863 = fired_release_1 & ldq_22_valid & ldq_22_bits_addr_valid & block_addr_matches_22_1;
  wire [31:0] _GEN_864 = ldq_22_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_865 = do_st_search_1 & ldq_22_valid & ldq_22_bits_addr_valid & _GEN_852 & ~ldq_22_bits_addr_is_virtual & _GEN_864[0] & dword_addr_matches_22_1 & (|_mask_overlap_T_90);
  wire        _GEN_866 = ~ldq_22_bits_forward_std_val | l_forward_stq_idx_22 != lcam_stq_idx_1 & (l_forward_stq_idx_22 < lcam_stq_idx_1 ^ l_forward_stq_idx_22 < ldq_22_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_22_bits_youngest_stq_idx);
  wire        _GEN_867 = do_ld_search_1 & ldq_22_valid & ldq_22_bits_addr_valid & ~ldq_22_bits_addr_is_virtual & dword_addr_matches_22_1 & (|_mask_overlap_T_90);
  wire        searcher_is_older_45 = lcam_ldq_idx_1 < 5'h16 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h16;
  wire        _GEN_868 = _GEN_867 & searcher_is_older_45 & _GEN_857;
  wire        _temp_bits_WIRE_1_54 = _GEN_863 ? _GEN_858 : _GEN_865 ? _GEN_866 | _GEN_858 : _GEN_868 | _GEN_858;
  reg         older_nacked_REG_45;
  wire        _GEN_869 = ~_GEN_851 | nacking_loads_22 | older_nacked_REG_45;
  wire        _GEN_870 = searcher_is_older_45 | _GEN_357;
  wire        _GEN_871 = _GEN_863 | _GEN_865;
  reg         io_dmem_s1_kill_1_REG_22;
  wire        _GEN_872 = _GEN_871 | ~_GEN_867 | _GEN_870 | ~_GEN_869;
  reg  [7:0]  casez_tmp_414;
  wire [14:0] _l_mask_mask_T_347 = 15'h1 << ldq_23_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_351 = 15'h3 << {12'h0, ldq_23_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_23_bits_uop_mem_size)
      2'b00:
        casez_tmp_414 = _l_mask_mask_T_347[7:0];
      2'b01:
        casez_tmp_414 = _l_mask_mask_T_351[7:0];
      2'b10:
        casez_tmp_414 = ldq_23_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_414 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_23_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h17;
  wire        l_forwarders_23_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h17;
  wire        l_is_forwarding_23 = l_forwarders_23_0 | l_forwarders_23_1;
  wire [4:0]  l_forward_stq_idx_23 = l_is_forwarding_23 ? (l_forwarders_23_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_23_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_23_bits_forward_stq_idx;
  wire        block_addr_matches_23_0 = lcam_addr_0[39:6] == ldq_23_bits_addr_bits[39:6];
  wire        block_addr_matches_23_1 = lcam_addr_1[39:6] == ldq_23_bits_addr_bits[39:6];
  wire        dword_addr_matches_23_0 = block_addr_matches_23_0 & lcam_addr_0[5:3] == ldq_23_bits_addr_bits[5:3];
  wire        dword_addr_matches_23_1 = block_addr_matches_23_1 & lcam_addr_1[5:3] == ldq_23_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_92 = casez_tmp_414 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_94 = casez_tmp_414 & casez_tmp_388;
  wire        _GEN_873 = fired_release_0 & ldq_23_valid & ldq_23_bits_addr_valid & block_addr_matches_23_0;
  wire        _GEN_874 = ldq_23_bits_executed | ldq_23_bits_succeeded;
  wire        _GEN_875 = _GEN_874 | l_is_forwarding_23;
  wire [31:0] _GEN_876 = ldq_23_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_877 = do_st_search_0 & ldq_23_valid & ldq_23_bits_addr_valid & _GEN_875 & ~ldq_23_bits_addr_is_virtual & _GEN_876[0] & dword_addr_matches_23_0 & (|_mask_overlap_T_92);
  wire        _GEN_878 = ~ldq_23_bits_forward_std_val | l_forward_stq_idx_23 != lcam_stq_idx_0 & (l_forward_stq_idx_23 < lcam_stq_idx_0 ^ l_forward_stq_idx_23 < ldq_23_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_23_bits_youngest_stq_idx);
  wire        _GEN_879 = do_ld_search_0 & ldq_23_valid & ldq_23_bits_addr_valid & ~ldq_23_bits_addr_is_virtual & dword_addr_matches_23_0 & (|_mask_overlap_T_92);
  wire        searcher_is_older_46 = lcam_ldq_idx_0 < 5'h17 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h17;
  wire        _GEN_880 = _GEN_875 & ~s1_executing_loads_23 & ldq_23_bits_observed;
  wire        _GEN_881 = ~_GEN_873 & (_GEN_877 ? _GEN_878 : _GEN_879 & searcher_is_older_46 & _GEN_880);
  reg         older_nacked_REG_46;
  wire        _GEN_882 = ~_GEN_874 | nacking_loads_23 | older_nacked_REG_46;
  wire        _GEN_883 = searcher_is_older_46 | _GEN_318;
  wire        _GEN_884 = _GEN_873 | _GEN_877;
  reg         io_dmem_s1_kill_0_REG_23;
  wire        _GEN_885 = _GEN_884 | ~_GEN_879 | _GEN_883 | ~_GEN_882;
  wire        _GEN_886 = fired_release_1 & ldq_23_valid & ldq_23_bits_addr_valid & block_addr_matches_23_1;
  wire [31:0] _GEN_887 = ldq_23_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_888 = do_st_search_1 & ldq_23_valid & ldq_23_bits_addr_valid & _GEN_875 & ~ldq_23_bits_addr_is_virtual & _GEN_887[0] & dword_addr_matches_23_1 & (|_mask_overlap_T_94);
  wire        _GEN_889 = ~ldq_23_bits_forward_std_val | l_forward_stq_idx_23 != lcam_stq_idx_1 & (l_forward_stq_idx_23 < lcam_stq_idx_1 ^ l_forward_stq_idx_23 < ldq_23_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_23_bits_youngest_stq_idx);
  wire        _GEN_890 = do_ld_search_1 & ldq_23_valid & ldq_23_bits_addr_valid & ~ldq_23_bits_addr_is_virtual & dword_addr_matches_23_1 & (|_mask_overlap_T_94);
  wire        searcher_is_older_47 = lcam_ldq_idx_1 < 5'h17 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h17;
  wire        _GEN_891 = _GEN_890 & searcher_is_older_47 & _GEN_880;
  wire        _temp_bits_WIRE_1_55 = _GEN_886 ? _GEN_881 : _GEN_888 ? _GEN_889 | _GEN_881 : _GEN_891 | _GEN_881;
  reg         older_nacked_REG_47;
  wire        _GEN_892 = ~_GEN_874 | nacking_loads_23 | older_nacked_REG_47;
  wire        _GEN_893 = searcher_is_older_47 | _GEN_358;
  wire        _GEN_894 = _GEN_886 | _GEN_888;
  reg         io_dmem_s1_kill_1_REG_23;
  wire        _GEN_895 = _GEN_894 | ~_GEN_890 | _GEN_893 | ~_GEN_892;
  reg  [7:0]  casez_tmp_415;
  wire [14:0] _l_mask_mask_T_362 = 15'h1 << ldq_24_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_366 = 15'h3 << {12'h0, ldq_24_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_24_bits_uop_mem_size)
      2'b00:
        casez_tmp_415 = _l_mask_mask_T_362[7:0];
      2'b01:
        casez_tmp_415 = _l_mask_mask_T_366[7:0];
      2'b10:
        casez_tmp_415 = ldq_24_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_415 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_24_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h18;
  wire        l_forwarders_24_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h18;
  wire        l_is_forwarding_24 = l_forwarders_24_0 | l_forwarders_24_1;
  wire [4:0]  l_forward_stq_idx_24 = l_is_forwarding_24 ? (l_forwarders_24_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_24_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_24_bits_forward_stq_idx;
  wire        block_addr_matches_24_0 = lcam_addr_0[39:6] == ldq_24_bits_addr_bits[39:6];
  wire        block_addr_matches_24_1 = lcam_addr_1[39:6] == ldq_24_bits_addr_bits[39:6];
  wire        dword_addr_matches_24_0 = block_addr_matches_24_0 & lcam_addr_0[5:3] == ldq_24_bits_addr_bits[5:3];
  wire        dword_addr_matches_24_1 = block_addr_matches_24_1 & lcam_addr_1[5:3] == ldq_24_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_96 = casez_tmp_415 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_98 = casez_tmp_415 & casez_tmp_388;
  wire        _GEN_896 = fired_release_0 & ldq_24_valid & ldq_24_bits_addr_valid & block_addr_matches_24_0;
  wire        _GEN_897 = ldq_24_bits_executed | ldq_24_bits_succeeded;
  wire        _GEN_898 = _GEN_897 | l_is_forwarding_24;
  wire [31:0] _GEN_899 = ldq_24_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_900 = do_st_search_0 & ldq_24_valid & ldq_24_bits_addr_valid & _GEN_898 & ~ldq_24_bits_addr_is_virtual & _GEN_899[0] & dword_addr_matches_24_0 & (|_mask_overlap_T_96);
  wire        _GEN_901 = ~ldq_24_bits_forward_std_val | l_forward_stq_idx_24 != lcam_stq_idx_0 & (l_forward_stq_idx_24 < lcam_stq_idx_0 ^ l_forward_stq_idx_24 < ldq_24_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_24_bits_youngest_stq_idx);
  wire        _GEN_902 = do_ld_search_0 & ldq_24_valid & ldq_24_bits_addr_valid & ~ldq_24_bits_addr_is_virtual & dword_addr_matches_24_0 & (|_mask_overlap_T_96);
  wire        searcher_is_older_48 = lcam_ldq_idx_0[4:3] != 2'h3 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h18;
  wire        _GEN_903 = _GEN_898 & ~s1_executing_loads_24 & ldq_24_bits_observed;
  wire        _GEN_904 = ~_GEN_896 & (_GEN_900 ? _GEN_901 : _GEN_902 & searcher_is_older_48 & _GEN_903);
  reg         older_nacked_REG_48;
  wire        _GEN_905 = ~_GEN_897 | nacking_loads_24 | older_nacked_REG_48;
  wire        _GEN_906 = searcher_is_older_48 | _GEN_319;
  wire        _GEN_907 = _GEN_896 | _GEN_900;
  reg         io_dmem_s1_kill_0_REG_24;
  wire        _GEN_908 = _GEN_907 | ~_GEN_902 | _GEN_906 | ~_GEN_905;
  wire        _GEN_909 = fired_release_1 & ldq_24_valid & ldq_24_bits_addr_valid & block_addr_matches_24_1;
  wire [31:0] _GEN_910 = ldq_24_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_911 = do_st_search_1 & ldq_24_valid & ldq_24_bits_addr_valid & _GEN_898 & ~ldq_24_bits_addr_is_virtual & _GEN_910[0] & dword_addr_matches_24_1 & (|_mask_overlap_T_98);
  wire        _GEN_912 = ~ldq_24_bits_forward_std_val | l_forward_stq_idx_24 != lcam_stq_idx_1 & (l_forward_stq_idx_24 < lcam_stq_idx_1 ^ l_forward_stq_idx_24 < ldq_24_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_24_bits_youngest_stq_idx);
  wire        _GEN_913 = do_ld_search_1 & ldq_24_valid & ldq_24_bits_addr_valid & ~ldq_24_bits_addr_is_virtual & dword_addr_matches_24_1 & (|_mask_overlap_T_98);
  wire        searcher_is_older_49 = lcam_ldq_idx_1[4:3] != 2'h3 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h18;
  wire        _GEN_914 = _GEN_913 & searcher_is_older_49 & _GEN_903;
  wire        _temp_bits_WIRE_1_56 = _GEN_909 ? _GEN_904 : _GEN_911 ? _GEN_912 | _GEN_904 : _GEN_914 | _GEN_904;
  reg         older_nacked_REG_49;
  wire        _GEN_915 = ~_GEN_897 | nacking_loads_24 | older_nacked_REG_49;
  wire        _GEN_916 = searcher_is_older_49 | _GEN_359;
  wire        _GEN_917 = _GEN_909 | _GEN_911;
  reg         io_dmem_s1_kill_1_REG_24;
  wire        _GEN_918 = _GEN_917 | ~_GEN_913 | _GEN_916 | ~_GEN_915;
  reg  [7:0]  casez_tmp_416;
  wire [14:0] _l_mask_mask_T_377 = 15'h1 << ldq_25_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_381 = 15'h3 << {12'h0, ldq_25_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_25_bits_uop_mem_size)
      2'b00:
        casez_tmp_416 = _l_mask_mask_T_377[7:0];
      2'b01:
        casez_tmp_416 = _l_mask_mask_T_381[7:0];
      2'b10:
        casez_tmp_416 = ldq_25_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_416 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_25_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h19;
  wire        l_forwarders_25_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h19;
  wire        l_is_forwarding_25 = l_forwarders_25_0 | l_forwarders_25_1;
  wire [4:0]  l_forward_stq_idx_25 = l_is_forwarding_25 ? (l_forwarders_25_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_25_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_25_bits_forward_stq_idx;
  wire        block_addr_matches_25_0 = lcam_addr_0[39:6] == ldq_25_bits_addr_bits[39:6];
  wire        block_addr_matches_25_1 = lcam_addr_1[39:6] == ldq_25_bits_addr_bits[39:6];
  wire        dword_addr_matches_25_0 = block_addr_matches_25_0 & lcam_addr_0[5:3] == ldq_25_bits_addr_bits[5:3];
  wire        dword_addr_matches_25_1 = block_addr_matches_25_1 & lcam_addr_1[5:3] == ldq_25_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_100 = casez_tmp_416 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_102 = casez_tmp_416 & casez_tmp_388;
  wire        _GEN_919 = fired_release_0 & ldq_25_valid & ldq_25_bits_addr_valid & block_addr_matches_25_0;
  wire        _GEN_920 = ldq_25_bits_executed | ldq_25_bits_succeeded;
  wire        _GEN_921 = _GEN_920 | l_is_forwarding_25;
  wire [31:0] _GEN_922 = ldq_25_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_923 = do_st_search_0 & ldq_25_valid & ldq_25_bits_addr_valid & _GEN_921 & ~ldq_25_bits_addr_is_virtual & _GEN_922[0] & dword_addr_matches_25_0 & (|_mask_overlap_T_100);
  wire        _GEN_924 = ~ldq_25_bits_forward_std_val | l_forward_stq_idx_25 != lcam_stq_idx_0 & (l_forward_stq_idx_25 < lcam_stq_idx_0 ^ l_forward_stq_idx_25 < ldq_25_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_25_bits_youngest_stq_idx);
  wire        _GEN_925 = do_ld_search_0 & ldq_25_valid & ldq_25_bits_addr_valid & ~ldq_25_bits_addr_is_virtual & dword_addr_matches_25_0 & (|_mask_overlap_T_100);
  wire        searcher_is_older_50 = lcam_ldq_idx_0 < 5'h19 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h19;
  wire        _GEN_926 = _GEN_921 & ~s1_executing_loads_25 & ldq_25_bits_observed;
  wire        _GEN_927 = ~_GEN_919 & (_GEN_923 ? _GEN_924 : _GEN_925 & searcher_is_older_50 & _GEN_926);
  reg         older_nacked_REG_50;
  wire        _GEN_928 = ~_GEN_920 | nacking_loads_25 | older_nacked_REG_50;
  wire        _GEN_929 = searcher_is_older_50 | _GEN_320;
  wire        _GEN_930 = _GEN_919 | _GEN_923;
  reg         io_dmem_s1_kill_0_REG_25;
  wire        _GEN_931 = _GEN_930 | ~_GEN_925 | _GEN_929 | ~_GEN_928;
  wire        _GEN_932 = fired_release_1 & ldq_25_valid & ldq_25_bits_addr_valid & block_addr_matches_25_1;
  wire [31:0] _GEN_933 = ldq_25_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_934 = do_st_search_1 & ldq_25_valid & ldq_25_bits_addr_valid & _GEN_921 & ~ldq_25_bits_addr_is_virtual & _GEN_933[0] & dword_addr_matches_25_1 & (|_mask_overlap_T_102);
  wire        _GEN_935 = ~ldq_25_bits_forward_std_val | l_forward_stq_idx_25 != lcam_stq_idx_1 & (l_forward_stq_idx_25 < lcam_stq_idx_1 ^ l_forward_stq_idx_25 < ldq_25_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_25_bits_youngest_stq_idx);
  wire        _GEN_936 = do_ld_search_1 & ldq_25_valid & ldq_25_bits_addr_valid & ~ldq_25_bits_addr_is_virtual & dword_addr_matches_25_1 & (|_mask_overlap_T_102);
  wire        searcher_is_older_51 = lcam_ldq_idx_1 < 5'h19 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h19;
  wire        _GEN_937 = _GEN_936 & searcher_is_older_51 & _GEN_926;
  wire        _temp_bits_WIRE_1_57 = _GEN_932 ? _GEN_927 : _GEN_934 ? _GEN_935 | _GEN_927 : _GEN_937 | _GEN_927;
  reg         older_nacked_REG_51;
  wire        _GEN_938 = ~_GEN_920 | nacking_loads_25 | older_nacked_REG_51;
  wire        _GEN_939 = searcher_is_older_51 | _GEN_360;
  wire        _GEN_940 = _GEN_932 | _GEN_934;
  reg         io_dmem_s1_kill_1_REG_25;
  wire        _GEN_941 = _GEN_940 | ~_GEN_936 | _GEN_939 | ~_GEN_938;
  reg  [7:0]  casez_tmp_417;
  wire [14:0] _l_mask_mask_T_392 = 15'h1 << ldq_26_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_396 = 15'h3 << {12'h0, ldq_26_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_26_bits_uop_mem_size)
      2'b00:
        casez_tmp_417 = _l_mask_mask_T_392[7:0];
      2'b01:
        casez_tmp_417 = _l_mask_mask_T_396[7:0];
      2'b10:
        casez_tmp_417 = ldq_26_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_417 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_26_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1A;
  wire        l_forwarders_26_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1A;
  wire        l_is_forwarding_26 = l_forwarders_26_0 | l_forwarders_26_1;
  wire [4:0]  l_forward_stq_idx_26 = l_is_forwarding_26 ? (l_forwarders_26_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_26_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_26_bits_forward_stq_idx;
  wire        block_addr_matches_26_0 = lcam_addr_0[39:6] == ldq_26_bits_addr_bits[39:6];
  wire        block_addr_matches_26_1 = lcam_addr_1[39:6] == ldq_26_bits_addr_bits[39:6];
  wire        dword_addr_matches_26_0 = block_addr_matches_26_0 & lcam_addr_0[5:3] == ldq_26_bits_addr_bits[5:3];
  wire        dword_addr_matches_26_1 = block_addr_matches_26_1 & lcam_addr_1[5:3] == ldq_26_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_104 = casez_tmp_417 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_106 = casez_tmp_417 & casez_tmp_388;
  wire        _GEN_942 = fired_release_0 & ldq_26_valid & ldq_26_bits_addr_valid & block_addr_matches_26_0;
  wire        _GEN_943 = ldq_26_bits_executed | ldq_26_bits_succeeded;
  wire        _GEN_944 = _GEN_943 | l_is_forwarding_26;
  wire [31:0] _GEN_945 = ldq_26_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_946 = do_st_search_0 & ldq_26_valid & ldq_26_bits_addr_valid & _GEN_944 & ~ldq_26_bits_addr_is_virtual & _GEN_945[0] & dword_addr_matches_26_0 & (|_mask_overlap_T_104);
  wire        _GEN_947 = ~ldq_26_bits_forward_std_val | l_forward_stq_idx_26 != lcam_stq_idx_0 & (l_forward_stq_idx_26 < lcam_stq_idx_0 ^ l_forward_stq_idx_26 < ldq_26_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_26_bits_youngest_stq_idx);
  wire        _GEN_948 = do_ld_search_0 & ldq_26_valid & ldq_26_bits_addr_valid & ~ldq_26_bits_addr_is_virtual & dword_addr_matches_26_0 & (|_mask_overlap_T_104);
  wire        searcher_is_older_52 = lcam_ldq_idx_0 < 5'h1A ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h1A;
  wire        _GEN_949 = _GEN_944 & ~s1_executing_loads_26 & ldq_26_bits_observed;
  wire        _GEN_950 = ~_GEN_942 & (_GEN_946 ? _GEN_947 : _GEN_948 & searcher_is_older_52 & _GEN_949);
  reg         older_nacked_REG_52;
  wire        _GEN_951 = ~_GEN_943 | nacking_loads_26 | older_nacked_REG_52;
  wire        _GEN_952 = searcher_is_older_52 | _GEN_321;
  wire        _GEN_953 = _GEN_942 | _GEN_946;
  reg         io_dmem_s1_kill_0_REG_26;
  wire        _GEN_954 = _GEN_953 | ~_GEN_948 | _GEN_952 | ~_GEN_951;
  wire        _GEN_955 = fired_release_1 & ldq_26_valid & ldq_26_bits_addr_valid & block_addr_matches_26_1;
  wire [31:0] _GEN_956 = ldq_26_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_957 = do_st_search_1 & ldq_26_valid & ldq_26_bits_addr_valid & _GEN_944 & ~ldq_26_bits_addr_is_virtual & _GEN_956[0] & dword_addr_matches_26_1 & (|_mask_overlap_T_106);
  wire        _GEN_958 = ~ldq_26_bits_forward_std_val | l_forward_stq_idx_26 != lcam_stq_idx_1 & (l_forward_stq_idx_26 < lcam_stq_idx_1 ^ l_forward_stq_idx_26 < ldq_26_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_26_bits_youngest_stq_idx);
  wire        _GEN_959 = do_ld_search_1 & ldq_26_valid & ldq_26_bits_addr_valid & ~ldq_26_bits_addr_is_virtual & dword_addr_matches_26_1 & (|_mask_overlap_T_106);
  wire        searcher_is_older_53 = lcam_ldq_idx_1 < 5'h1A ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h1A;
  wire        _GEN_960 = _GEN_959 & searcher_is_older_53 & _GEN_949;
  wire        _temp_bits_WIRE_1_58 = _GEN_955 ? _GEN_950 : _GEN_957 ? _GEN_958 | _GEN_950 : _GEN_960 | _GEN_950;
  reg         older_nacked_REG_53;
  wire        _GEN_961 = ~_GEN_943 | nacking_loads_26 | older_nacked_REG_53;
  wire        _GEN_962 = searcher_is_older_53 | _GEN_361;
  wire        _GEN_963 = _GEN_955 | _GEN_957;
  reg         io_dmem_s1_kill_1_REG_26;
  wire        _GEN_964 = _GEN_963 | ~_GEN_959 | _GEN_962 | ~_GEN_961;
  reg  [7:0]  casez_tmp_418;
  wire [14:0] _l_mask_mask_T_407 = 15'h1 << ldq_27_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_411 = 15'h3 << {12'h0, ldq_27_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_27_bits_uop_mem_size)
      2'b00:
        casez_tmp_418 = _l_mask_mask_T_407[7:0];
      2'b01:
        casez_tmp_418 = _l_mask_mask_T_411[7:0];
      2'b10:
        casez_tmp_418 = ldq_27_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_418 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_27_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1B;
  wire        l_forwarders_27_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1B;
  wire        l_is_forwarding_27 = l_forwarders_27_0 | l_forwarders_27_1;
  wire [4:0]  l_forward_stq_idx_27 = l_is_forwarding_27 ? (l_forwarders_27_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_27_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_27_bits_forward_stq_idx;
  wire        block_addr_matches_27_0 = lcam_addr_0[39:6] == ldq_27_bits_addr_bits[39:6];
  wire        block_addr_matches_27_1 = lcam_addr_1[39:6] == ldq_27_bits_addr_bits[39:6];
  wire        dword_addr_matches_27_0 = block_addr_matches_27_0 & lcam_addr_0[5:3] == ldq_27_bits_addr_bits[5:3];
  wire        dword_addr_matches_27_1 = block_addr_matches_27_1 & lcam_addr_1[5:3] == ldq_27_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_108 = casez_tmp_418 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_110 = casez_tmp_418 & casez_tmp_388;
  wire        _GEN_965 = fired_release_0 & ldq_27_valid & ldq_27_bits_addr_valid & block_addr_matches_27_0;
  wire        _GEN_966 = ldq_27_bits_executed | ldq_27_bits_succeeded;
  wire        _GEN_967 = _GEN_966 | l_is_forwarding_27;
  wire [31:0] _GEN_968 = ldq_27_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_969 = do_st_search_0 & ldq_27_valid & ldq_27_bits_addr_valid & _GEN_967 & ~ldq_27_bits_addr_is_virtual & _GEN_968[0] & dword_addr_matches_27_0 & (|_mask_overlap_T_108);
  wire        _GEN_970 = ~ldq_27_bits_forward_std_val | l_forward_stq_idx_27 != lcam_stq_idx_0 & (l_forward_stq_idx_27 < lcam_stq_idx_0 ^ l_forward_stq_idx_27 < ldq_27_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_27_bits_youngest_stq_idx);
  wire        _GEN_971 = do_ld_search_0 & ldq_27_valid & ldq_27_bits_addr_valid & ~ldq_27_bits_addr_is_virtual & dword_addr_matches_27_0 & (|_mask_overlap_T_108);
  wire        searcher_is_older_54 = lcam_ldq_idx_0 < 5'h1B ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h1B;
  wire        _GEN_972 = _GEN_967 & ~s1_executing_loads_27 & ldq_27_bits_observed;
  wire        _GEN_973 = ~_GEN_965 & (_GEN_969 ? _GEN_970 : _GEN_971 & searcher_is_older_54 & _GEN_972);
  reg         older_nacked_REG_54;
  wire        _GEN_974 = ~_GEN_966 | nacking_loads_27 | older_nacked_REG_54;
  wire        _GEN_975 = searcher_is_older_54 | _GEN_322;
  wire        _GEN_976 = _GEN_965 | _GEN_969;
  reg         io_dmem_s1_kill_0_REG_27;
  wire        _GEN_977 = _GEN_976 | ~_GEN_971 | _GEN_975 | ~_GEN_974;
  wire        _GEN_978 = fired_release_1 & ldq_27_valid & ldq_27_bits_addr_valid & block_addr_matches_27_1;
  wire [31:0] _GEN_979 = ldq_27_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_980 = do_st_search_1 & ldq_27_valid & ldq_27_bits_addr_valid & _GEN_967 & ~ldq_27_bits_addr_is_virtual & _GEN_979[0] & dword_addr_matches_27_1 & (|_mask_overlap_T_110);
  wire        _GEN_981 = ~ldq_27_bits_forward_std_val | l_forward_stq_idx_27 != lcam_stq_idx_1 & (l_forward_stq_idx_27 < lcam_stq_idx_1 ^ l_forward_stq_idx_27 < ldq_27_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_27_bits_youngest_stq_idx);
  wire        _GEN_982 = do_ld_search_1 & ldq_27_valid & ldq_27_bits_addr_valid & ~ldq_27_bits_addr_is_virtual & dword_addr_matches_27_1 & (|_mask_overlap_T_110);
  wire        searcher_is_older_55 = lcam_ldq_idx_1 < 5'h1B ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h1B;
  wire        _GEN_983 = _GEN_982 & searcher_is_older_55 & _GEN_972;
  wire        _temp_bits_WIRE_1_59 = _GEN_978 ? _GEN_973 : _GEN_980 ? _GEN_981 | _GEN_973 : _GEN_983 | _GEN_973;
  reg         older_nacked_REG_55;
  wire        _GEN_984 = ~_GEN_966 | nacking_loads_27 | older_nacked_REG_55;
  wire        _GEN_985 = searcher_is_older_55 | _GEN_362;
  wire        _GEN_986 = _GEN_978 | _GEN_980;
  reg         io_dmem_s1_kill_1_REG_27;
  wire        _GEN_987 = _GEN_986 | ~_GEN_982 | _GEN_985 | ~_GEN_984;
  reg  [7:0]  casez_tmp_419;
  wire [14:0] _l_mask_mask_T_422 = 15'h1 << ldq_28_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_426 = 15'h3 << {12'h0, ldq_28_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_28_bits_uop_mem_size)
      2'b00:
        casez_tmp_419 = _l_mask_mask_T_422[7:0];
      2'b01:
        casez_tmp_419 = _l_mask_mask_T_426[7:0];
      2'b10:
        casez_tmp_419 = ldq_28_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_419 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_28_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1C;
  wire        l_forwarders_28_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1C;
  wire        l_is_forwarding_28 = l_forwarders_28_0 | l_forwarders_28_1;
  wire [4:0]  l_forward_stq_idx_28 = l_is_forwarding_28 ? (l_forwarders_28_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_28_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_28_bits_forward_stq_idx;
  wire        block_addr_matches_28_0 = lcam_addr_0[39:6] == ldq_28_bits_addr_bits[39:6];
  wire        block_addr_matches_28_1 = lcam_addr_1[39:6] == ldq_28_bits_addr_bits[39:6];
  wire        dword_addr_matches_28_0 = block_addr_matches_28_0 & lcam_addr_0[5:3] == ldq_28_bits_addr_bits[5:3];
  wire        dword_addr_matches_28_1 = block_addr_matches_28_1 & lcam_addr_1[5:3] == ldq_28_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_112 = casez_tmp_419 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_114 = casez_tmp_419 & casez_tmp_388;
  wire        _GEN_988 = fired_release_0 & ldq_28_valid & ldq_28_bits_addr_valid & block_addr_matches_28_0;
  wire        _GEN_989 = ldq_28_bits_executed | ldq_28_bits_succeeded;
  wire        _GEN_990 = _GEN_989 | l_is_forwarding_28;
  wire [31:0] _GEN_991 = ldq_28_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_992 = do_st_search_0 & ldq_28_valid & ldq_28_bits_addr_valid & _GEN_990 & ~ldq_28_bits_addr_is_virtual & _GEN_991[0] & dword_addr_matches_28_0 & (|_mask_overlap_T_112);
  wire        _GEN_993 = ~ldq_28_bits_forward_std_val | l_forward_stq_idx_28 != lcam_stq_idx_0 & (l_forward_stq_idx_28 < lcam_stq_idx_0 ^ l_forward_stq_idx_28 < ldq_28_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_28_bits_youngest_stq_idx);
  wire        _GEN_994 = do_ld_search_0 & ldq_28_valid & ldq_28_bits_addr_valid & ~ldq_28_bits_addr_is_virtual & dword_addr_matches_28_0 & (|_mask_overlap_T_112);
  wire        searcher_is_older_56 = lcam_ldq_idx_0[4:2] != 3'h7 ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h1C;
  wire        _GEN_995 = _GEN_990 & ~s1_executing_loads_28 & ldq_28_bits_observed;
  wire        _GEN_996 = ~_GEN_988 & (_GEN_992 ? _GEN_993 : _GEN_994 & searcher_is_older_56 & _GEN_995);
  reg         older_nacked_REG_56;
  wire        _GEN_997 = ~_GEN_989 | nacking_loads_28 | older_nacked_REG_56;
  wire        _GEN_998 = searcher_is_older_56 | _GEN_323;
  wire        _GEN_999 = _GEN_988 | _GEN_992;
  reg         io_dmem_s1_kill_0_REG_28;
  wire        _GEN_1000 = _GEN_999 | ~_GEN_994 | _GEN_998 | ~_GEN_997;
  wire        _GEN_1001 = fired_release_1 & ldq_28_valid & ldq_28_bits_addr_valid & block_addr_matches_28_1;
  wire [31:0] _GEN_1002 = ldq_28_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_1003 = do_st_search_1 & ldq_28_valid & ldq_28_bits_addr_valid & _GEN_990 & ~ldq_28_bits_addr_is_virtual & _GEN_1002[0] & dword_addr_matches_28_1 & (|_mask_overlap_T_114);
  wire        _GEN_1004 = ~ldq_28_bits_forward_std_val | l_forward_stq_idx_28 != lcam_stq_idx_1 & (l_forward_stq_idx_28 < lcam_stq_idx_1 ^ l_forward_stq_idx_28 < ldq_28_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_28_bits_youngest_stq_idx);
  wire        _GEN_1005 = do_ld_search_1 & ldq_28_valid & ldq_28_bits_addr_valid & ~ldq_28_bits_addr_is_virtual & dword_addr_matches_28_1 & (|_mask_overlap_T_114);
  wire        searcher_is_older_57 = lcam_ldq_idx_1[4:2] != 3'h7 ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h1C;
  wire        _GEN_1006 = _GEN_1005 & searcher_is_older_57 & _GEN_995;
  wire        _temp_bits_WIRE_1_60 = _GEN_1001 ? _GEN_996 : _GEN_1003 ? _GEN_1004 | _GEN_996 : _GEN_1006 | _GEN_996;
  reg         older_nacked_REG_57;
  wire        _GEN_1007 = ~_GEN_989 | nacking_loads_28 | older_nacked_REG_57;
  wire        _GEN_1008 = searcher_is_older_57 | _GEN_363;
  wire        _GEN_1009 = _GEN_1001 | _GEN_1003;
  reg         io_dmem_s1_kill_1_REG_28;
  wire        _GEN_1010 = _GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~_GEN_1007;
  reg  [7:0]  casez_tmp_420;
  wire [14:0] _l_mask_mask_T_437 = 15'h1 << ldq_29_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_441 = 15'h3 << {12'h0, ldq_29_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_29_bits_uop_mem_size)
      2'b00:
        casez_tmp_420 = _l_mask_mask_T_437[7:0];
      2'b01:
        casez_tmp_420 = _l_mask_mask_T_441[7:0];
      2'b10:
        casez_tmp_420 = ldq_29_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_420 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_29_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1D;
  wire        l_forwarders_29_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1D;
  wire        l_is_forwarding_29 = l_forwarders_29_0 | l_forwarders_29_1;
  wire [4:0]  l_forward_stq_idx_29 = l_is_forwarding_29 ? (l_forwarders_29_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_29_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_29_bits_forward_stq_idx;
  wire        block_addr_matches_29_0 = lcam_addr_0[39:6] == ldq_29_bits_addr_bits[39:6];
  wire        block_addr_matches_29_1 = lcam_addr_1[39:6] == ldq_29_bits_addr_bits[39:6];
  wire        dword_addr_matches_29_0 = block_addr_matches_29_0 & lcam_addr_0[5:3] == ldq_29_bits_addr_bits[5:3];
  wire        dword_addr_matches_29_1 = block_addr_matches_29_1 & lcam_addr_1[5:3] == ldq_29_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_116 = casez_tmp_420 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_118 = casez_tmp_420 & casez_tmp_388;
  wire        _GEN_1011 = fired_release_0 & ldq_29_valid & ldq_29_bits_addr_valid & block_addr_matches_29_0;
  wire        _GEN_1012 = ldq_29_bits_executed | ldq_29_bits_succeeded;
  wire        _GEN_1013 = _GEN_1012 | l_is_forwarding_29;
  wire [31:0] _GEN_1014 = ldq_29_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_1015 = do_st_search_0 & ldq_29_valid & ldq_29_bits_addr_valid & _GEN_1013 & ~ldq_29_bits_addr_is_virtual & _GEN_1014[0] & dword_addr_matches_29_0 & (|_mask_overlap_T_116);
  wire        _GEN_1016 = ~ldq_29_bits_forward_std_val | l_forward_stq_idx_29 != lcam_stq_idx_0 & (l_forward_stq_idx_29 < lcam_stq_idx_0 ^ l_forward_stq_idx_29 < ldq_29_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_29_bits_youngest_stq_idx);
  wire        _GEN_1017 = do_ld_search_0 & ldq_29_valid & ldq_29_bits_addr_valid & ~ldq_29_bits_addr_is_virtual & dword_addr_matches_29_0 & (|_mask_overlap_T_116);
  wire        searcher_is_older_58 = lcam_ldq_idx_0 < 5'h1D ^ lcam_ldq_idx_0 < ldq_head ^ ldq_head > 5'h1D;
  wire        _GEN_1018 = _GEN_1013 & ~s1_executing_loads_29 & ldq_29_bits_observed;
  wire        _GEN_1019 = ~_GEN_1011 & (_GEN_1015 ? _GEN_1016 : _GEN_1017 & searcher_is_older_58 & _GEN_1018);
  reg         older_nacked_REG_58;
  wire        _GEN_1020 = ~_GEN_1012 | nacking_loads_29 | older_nacked_REG_58;
  wire        _GEN_1021 = searcher_is_older_58 | _GEN_324;
  wire        _GEN_1022 = _GEN_1011 | _GEN_1015;
  reg         io_dmem_s1_kill_0_REG_29;
  wire        _GEN_1023 = _GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~_GEN_1020;
  wire        _GEN_1024 = fired_release_1 & ldq_29_valid & ldq_29_bits_addr_valid & block_addr_matches_29_1;
  wire [31:0] _GEN_1025 = ldq_29_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_1026 = do_st_search_1 & ldq_29_valid & ldq_29_bits_addr_valid & _GEN_1013 & ~ldq_29_bits_addr_is_virtual & _GEN_1025[0] & dword_addr_matches_29_1 & (|_mask_overlap_T_118);
  wire        _GEN_1027 = ~ldq_29_bits_forward_std_val | l_forward_stq_idx_29 != lcam_stq_idx_1 & (l_forward_stq_idx_29 < lcam_stq_idx_1 ^ l_forward_stq_idx_29 < ldq_29_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_29_bits_youngest_stq_idx);
  wire        _GEN_1028 = do_ld_search_1 & ldq_29_valid & ldq_29_bits_addr_valid & ~ldq_29_bits_addr_is_virtual & dword_addr_matches_29_1 & (|_mask_overlap_T_118);
  wire        searcher_is_older_59 = lcam_ldq_idx_1 < 5'h1D ^ lcam_ldq_idx_1 < ldq_head ^ ldq_head > 5'h1D;
  wire        _GEN_1029 = _GEN_1028 & searcher_is_older_59 & _GEN_1018;
  wire        _temp_bits_WIRE_1_61 = _GEN_1024 ? _GEN_1019 : _GEN_1026 ? _GEN_1027 | _GEN_1019 : _GEN_1029 | _GEN_1019;
  reg         older_nacked_REG_59;
  wire        _GEN_1030 = ~_GEN_1012 | nacking_loads_29 | older_nacked_REG_59;
  wire        _GEN_1031 = searcher_is_older_59 | _GEN_364;
  wire        _GEN_1032 = _GEN_1024 | _GEN_1026;
  reg         io_dmem_s1_kill_1_REG_29;
  wire        _GEN_1033 = _GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~_GEN_1030;
  reg  [7:0]  casez_tmp_421;
  wire [14:0] _l_mask_mask_T_452 = 15'h1 << ldq_30_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_456 = 15'h3 << {12'h0, ldq_30_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_30_bits_uop_mem_size)
      2'b00:
        casez_tmp_421 = _l_mask_mask_T_452[7:0];
      2'b01:
        casez_tmp_421 = _l_mask_mask_T_456[7:0];
      2'b10:
        casez_tmp_421 = ldq_30_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_421 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_30_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1E;
  wire        l_forwarders_30_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1E;
  wire        l_is_forwarding_30 = l_forwarders_30_0 | l_forwarders_30_1;
  wire [4:0]  l_forward_stq_idx_30 = l_is_forwarding_30 ? (l_forwarders_30_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_30_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_30_bits_forward_stq_idx;
  wire        block_addr_matches_30_0 = lcam_addr_0[39:6] == ldq_30_bits_addr_bits[39:6];
  wire        block_addr_matches_30_1 = lcam_addr_1[39:6] == ldq_30_bits_addr_bits[39:6];
  wire        dword_addr_matches_30_0 = block_addr_matches_30_0 & lcam_addr_0[5:3] == ldq_30_bits_addr_bits[5:3];
  wire        dword_addr_matches_30_1 = block_addr_matches_30_1 & lcam_addr_1[5:3] == ldq_30_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_120 = casez_tmp_421 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_122 = casez_tmp_421 & casez_tmp_388;
  wire        _GEN_1034 = fired_release_0 & ldq_30_valid & ldq_30_bits_addr_valid & block_addr_matches_30_0;
  wire        _GEN_1035 = ldq_30_bits_executed | ldq_30_bits_succeeded;
  wire        _GEN_1036 = _GEN_1035 | l_is_forwarding_30;
  wire [31:0] _GEN_1037 = ldq_30_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_1038 = do_st_search_0 & ldq_30_valid & ldq_30_bits_addr_valid & _GEN_1036 & ~ldq_30_bits_addr_is_virtual & _GEN_1037[0] & dword_addr_matches_30_0 & (|_mask_overlap_T_120);
  wire        _GEN_1039 = ~ldq_30_bits_forward_std_val | l_forward_stq_idx_30 != lcam_stq_idx_0 & (l_forward_stq_idx_30 < lcam_stq_idx_0 ^ l_forward_stq_idx_30 < ldq_30_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_30_bits_youngest_stq_idx);
  wire        _GEN_1040 = do_ld_search_0 & ldq_30_valid & ldq_30_bits_addr_valid & ~ldq_30_bits_addr_is_virtual & dword_addr_matches_30_0 & (|_mask_overlap_T_120);
  wire        searcher_is_older_60 = lcam_ldq_idx_0[4:1] != 4'hF ^ lcam_ldq_idx_0 < ldq_head ^ (&ldq_head);
  wire        _GEN_1041 = _GEN_1036 & ~s1_executing_loads_30 & ldq_30_bits_observed;
  wire        _GEN_1042 = ~_GEN_1034 & (_GEN_1038 ? _GEN_1039 : _GEN_1040 & searcher_is_older_60 & _GEN_1041);
  reg         older_nacked_REG_60;
  wire        _GEN_1043 = ~_GEN_1035 | nacking_loads_30 | older_nacked_REG_60;
  wire        _GEN_1044 = searcher_is_older_60 | _GEN_325;
  wire        _GEN_1045 = _GEN_1034 | _GEN_1038;
  reg         io_dmem_s1_kill_0_REG_30;
  wire        _GEN_1046 = _GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~_GEN_1043;
  wire        _GEN_1047 = fired_release_1 & ldq_30_valid & ldq_30_bits_addr_valid & block_addr_matches_30_1;
  wire [31:0] _GEN_1048 = ldq_30_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_1049 = do_st_search_1 & ldq_30_valid & ldq_30_bits_addr_valid & _GEN_1036 & ~ldq_30_bits_addr_is_virtual & _GEN_1048[0] & dword_addr_matches_30_1 & (|_mask_overlap_T_122);
  wire        _GEN_1050 = ~ldq_30_bits_forward_std_val | l_forward_stq_idx_30 != lcam_stq_idx_1 & (l_forward_stq_idx_30 < lcam_stq_idx_1 ^ l_forward_stq_idx_30 < ldq_30_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_30_bits_youngest_stq_idx);
  wire        _GEN_1051 = do_ld_search_1 & ldq_30_valid & ldq_30_bits_addr_valid & ~ldq_30_bits_addr_is_virtual & dword_addr_matches_30_1 & (|_mask_overlap_T_122);
  wire        searcher_is_older_61 = lcam_ldq_idx_1[4:1] != 4'hF ^ lcam_ldq_idx_1 < ldq_head ^ (&ldq_head);
  wire        _GEN_1052 = _GEN_1051 & searcher_is_older_61 & _GEN_1041;
  wire        _temp_bits_WIRE_1_62 = _GEN_1047 ? _GEN_1042 : _GEN_1049 ? _GEN_1050 | _GEN_1042 : _GEN_1052 | _GEN_1042;
  reg         older_nacked_REG_61;
  wire        _GEN_1053 = ~_GEN_1035 | nacking_loads_30 | older_nacked_REG_61;
  wire        _GEN_1054 = searcher_is_older_61 | _GEN_365;
  wire        _GEN_1055 = _GEN_1047 | _GEN_1049;
  reg         io_dmem_s1_kill_1_REG_30;
  wire        _GEN_1056 = _GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~_GEN_1053;
  reg  [7:0]  casez_tmp_422;
  wire [14:0] _l_mask_mask_T_467 = 15'h1 << ldq_31_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_471 = 15'h3 << {12'h0, ldq_31_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_31_bits_uop_mem_size)
      2'b00:
        casez_tmp_422 = _l_mask_mask_T_467[7:0];
      2'b01:
        casez_tmp_422 = _l_mask_mask_T_471[7:0];
      2'b10:
        casez_tmp_422 = ldq_31_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_422 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_31_0 = wb_forward_valid_0 & (&wb_forward_ldq_idx_0);
  wire        l_forwarders_31_1 = wb_forward_valid_1 & (&wb_forward_ldq_idx_1);
  wire        l_is_forwarding_31 = l_forwarders_31_0 | l_forwarders_31_1;
  wire [4:0]  l_forward_stq_idx_31 = l_is_forwarding_31 ? (l_forwarders_31_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_31_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_31_bits_forward_stq_idx;
  wire        block_addr_matches_31_0 = lcam_addr_0[39:6] == ldq_31_bits_addr_bits[39:6];
  wire        block_addr_matches_31_1 = lcam_addr_1[39:6] == ldq_31_bits_addr_bits[39:6];
  wire        dword_addr_matches_31_0 = block_addr_matches_31_0 & lcam_addr_0[5:3] == ldq_31_bits_addr_bits[5:3];
  wire        dword_addr_matches_31_1 = block_addr_matches_31_1 & lcam_addr_1[5:3] == ldq_31_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_124 = casez_tmp_422 & casez_tmp_387;
  wire [7:0]  _mask_overlap_T_126 = casez_tmp_422 & casez_tmp_388;
  wire        _GEN_1057 = fired_release_0 & ldq_31_valid & ldq_31_bits_addr_valid & block_addr_matches_31_0;
  wire        _GEN_1058 = ldq_31_bits_executed | ldq_31_bits_succeeded;
  wire        _GEN_1059 = _GEN_1058 | l_is_forwarding_31;
  wire [31:0] _GEN_1060 = ldq_31_bits_st_dep_mask >> _GEN_287;
  wire        _GEN_1061 = do_st_search_0 & ldq_31_valid & ldq_31_bits_addr_valid & _GEN_1059 & ~ldq_31_bits_addr_is_virtual & _GEN_1060[0] & dword_addr_matches_31_0 & (|_mask_overlap_T_124);
  wire        _GEN_1062 = ~ldq_31_bits_forward_std_val | l_forward_stq_idx_31 != lcam_stq_idx_0 & (l_forward_stq_idx_31 < lcam_stq_idx_0 ^ l_forward_stq_idx_31 < ldq_31_bits_youngest_stq_idx ^ lcam_stq_idx_0 < ldq_31_bits_youngest_stq_idx);
  wire        _GEN_1063 = do_ld_search_0 & ldq_31_valid & ldq_31_bits_addr_valid & ~ldq_31_bits_addr_is_virtual & dword_addr_matches_31_0 & (|_mask_overlap_T_124);
  wire        searcher_is_older_62 = lcam_ldq_idx_0 != 5'h1F ^ lcam_ldq_idx_0 < ldq_head;
  wire        _GEN_1064 = _GEN_1059 & ~s1_executing_loads_31 & ldq_31_bits_observed;
  wire        _GEN_1065 = ~_GEN_1057 & (_GEN_1061 ? _GEN_1062 : _GEN_1063 & searcher_is_older_62 & _GEN_1064);
  reg         older_nacked_REG_62;
  wire        _GEN_1066 = ~_GEN_1058 | nacking_loads_31 | older_nacked_REG_62;
  wire        _GEN_1067 = _GEN_1057 | _GEN_1061;
  reg         io_dmem_s1_kill_0_REG_31;
  wire        _GEN_1068 = _GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066);
  wire        _GEN_1069 = _GEN_1068 ? (_GEN_1046 ? (_GEN_1023 ? (_GEN_1000 ? (_GEN_977 ? (_GEN_954 ? (_GEN_931 ? (_GEN_908 ? (_GEN_885 ? (_GEN_862 ? (_GEN_839 ? (_GEN_816 ? (_GEN_793 ? (_GEN_770 ? (_GEN_747 ? (_GEN_724 ? (_GEN_701 ? (_GEN_678 ? (_GEN_655 ? (_GEN_632 ? (_GEN_609 ? (_GEN_586 ? (_GEN_563 ? (_GEN_540 ? (_GEN_517 ? (_GEN_494 ? (_GEN_471 ? (_GEN_448 ? (_GEN_425 ? (_GEN_402 ? (_GEN_379 ? ~_GEN_295 & _GEN_291 & ~searcher_is_older & _GEN_326 & io_dmem_s1_kill_0_REG : io_dmem_s1_kill_0_REG_1) : io_dmem_s1_kill_0_REG_2) : io_dmem_s1_kill_0_REG_3) : io_dmem_s1_kill_0_REG_4) : io_dmem_s1_kill_0_REG_5) : io_dmem_s1_kill_0_REG_6) : io_dmem_s1_kill_0_REG_7) : io_dmem_s1_kill_0_REG_8) : io_dmem_s1_kill_0_REG_9) : io_dmem_s1_kill_0_REG_10) : io_dmem_s1_kill_0_REG_11) : io_dmem_s1_kill_0_REG_12) : io_dmem_s1_kill_0_REG_13) : io_dmem_s1_kill_0_REG_14) : io_dmem_s1_kill_0_REG_15) : io_dmem_s1_kill_0_REG_16) : io_dmem_s1_kill_0_REG_17) : io_dmem_s1_kill_0_REG_18) : io_dmem_s1_kill_0_REG_19) : io_dmem_s1_kill_0_REG_20) : io_dmem_s1_kill_0_REG_21) : io_dmem_s1_kill_0_REG_22) : io_dmem_s1_kill_0_REG_23) : io_dmem_s1_kill_0_REG_24) : io_dmem_s1_kill_0_REG_25) : io_dmem_s1_kill_0_REG_26) : io_dmem_s1_kill_0_REG_27) : io_dmem_s1_kill_0_REG_28) : io_dmem_s1_kill_0_REG_29) : io_dmem_s1_kill_0_REG_30) : io_dmem_s1_kill_0_REG_31;
  wire        can_forward_0 = _GEN_1068 & _GEN_1046 & _GEN_1023 & _GEN_1000 & _GEN_977 & _GEN_954 & _GEN_931 & _GEN_908 & _GEN_885 & _GEN_862 & _GEN_839 & _GEN_816 & _GEN_793 & _GEN_770 & _GEN_747 & _GEN_724 & _GEN_701 & _GEN_678 & _GEN_655 & _GEN_632 & _GEN_609 & _GEN_586 & _GEN_563 & _GEN_540 & _GEN_517 & _GEN_494 & _GEN_471 & _GEN_448 & _GEN_425 & _GEN_402 & _GEN_379 & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~_GEN_326) & (_can_forward_T ? ~mem_tlb_uncacheable_0 : ~casez_tmp_389);
  wire        _GEN_1070 = fired_release_1 & ldq_31_valid & ldq_31_bits_addr_valid & block_addr_matches_31_1;
  wire [31:0] _GEN_1071 = ldq_31_bits_st_dep_mask >> _GEN_328;
  wire        _GEN_1072 = do_st_search_1 & ldq_31_valid & ldq_31_bits_addr_valid & _GEN_1059 & ~ldq_31_bits_addr_is_virtual & _GEN_1071[0] & dword_addr_matches_31_1 & (|_mask_overlap_T_126);
  wire        _GEN_1073 = ~ldq_31_bits_forward_std_val | l_forward_stq_idx_31 != lcam_stq_idx_1 & (l_forward_stq_idx_31 < lcam_stq_idx_1 ^ l_forward_stq_idx_31 < ldq_31_bits_youngest_stq_idx ^ lcam_stq_idx_1 < ldq_31_bits_youngest_stq_idx);
  wire        _GEN_1074 = do_ld_search_1 & ldq_31_valid & ldq_31_bits_addr_valid & ~ldq_31_bits_addr_is_virtual & dword_addr_matches_31_1 & (|_mask_overlap_T_126);
  wire        searcher_is_older_63 = lcam_ldq_idx_1 != 5'h1F ^ lcam_ldq_idx_1 < ldq_head;
  wire        _GEN_1075 = _GEN_1074 & searcher_is_older_63 & _GEN_1064;
  wire        _temp_bits_WIRE_1_63 = _GEN_1070 ? _GEN_1065 : _GEN_1072 ? _GEN_1073 | _GEN_1065 : _GEN_1075 | _GEN_1065;
  reg         older_nacked_REG_63;
  wire        _GEN_1076 = ~_GEN_1058 | nacking_loads_31 | older_nacked_REG_63;
  wire        _GEN_1077 = _GEN_1070 | _GEN_1072;
  reg         io_dmem_s1_kill_1_REG_31;
  wire        _GEN_1078 = _GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076);
  wire        _GEN_1079 = _GEN_1078 ? (_GEN_1056 ? (_GEN_1033 ? (_GEN_1010 ? (_GEN_987 ? (_GEN_964 ? (_GEN_941 ? (_GEN_918 ? (_GEN_895 ? (_GEN_872 ? (_GEN_849 ? (_GEN_826 ? (_GEN_803 ? (_GEN_780 ? (_GEN_757 ? (_GEN_734 ? (_GEN_711 ? (_GEN_688 ? (_GEN_665 ? (_GEN_642 ? (_GEN_619 ? (_GEN_596 ? (_GEN_573 ? (_GEN_550 ? (_GEN_527 ? (_GEN_504 ? (_GEN_481 ? (_GEN_458 ? (_GEN_435 ? (_GEN_412 ? (_GEN_389 ? ~_GEN_335 & _GEN_332 & ~searcher_is_older_1 & _GEN_366 & io_dmem_s1_kill_1_REG : io_dmem_s1_kill_1_REG_1) : io_dmem_s1_kill_1_REG_2) : io_dmem_s1_kill_1_REG_3) : io_dmem_s1_kill_1_REG_4) : io_dmem_s1_kill_1_REG_5) : io_dmem_s1_kill_1_REG_6) : io_dmem_s1_kill_1_REG_7) : io_dmem_s1_kill_1_REG_8) : io_dmem_s1_kill_1_REG_9) : io_dmem_s1_kill_1_REG_10) : io_dmem_s1_kill_1_REG_11) : io_dmem_s1_kill_1_REG_12) : io_dmem_s1_kill_1_REG_13) : io_dmem_s1_kill_1_REG_14) : io_dmem_s1_kill_1_REG_15) : io_dmem_s1_kill_1_REG_16) : io_dmem_s1_kill_1_REG_17) : io_dmem_s1_kill_1_REG_18) : io_dmem_s1_kill_1_REG_19) : io_dmem_s1_kill_1_REG_20) : io_dmem_s1_kill_1_REG_21) : io_dmem_s1_kill_1_REG_22) : io_dmem_s1_kill_1_REG_23) : io_dmem_s1_kill_1_REG_24) : io_dmem_s1_kill_1_REG_25) : io_dmem_s1_kill_1_REG_26) : io_dmem_s1_kill_1_REG_27) : io_dmem_s1_kill_1_REG_28) : io_dmem_s1_kill_1_REG_29) : io_dmem_s1_kill_1_REG_30) : io_dmem_s1_kill_1_REG_31;
  wire        can_forward_1 = _GEN_1078 & _GEN_1056 & _GEN_1033 & _GEN_1010 & _GEN_987 & _GEN_964 & _GEN_941 & _GEN_918 & _GEN_895 & _GEN_872 & _GEN_849 & _GEN_826 & _GEN_803 & _GEN_780 & _GEN_757 & _GEN_734 & _GEN_711 & _GEN_688 & _GEN_665 & _GEN_642 & _GEN_619 & _GEN_596 & _GEN_573 & _GEN_550 & _GEN_527 & _GEN_504 & _GEN_481 & _GEN_458 & _GEN_435 & _GEN_412 & _GEN_389 & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~_GEN_366) & (_can_forward_T_6 ? ~mem_tlb_uncacheable_1 : ~casez_tmp_390);
  wire        dword_addr_matches_32_0 = stq_0_bits_addr_valid & ~stq_0_bits_addr_is_virtual & stq_0_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_32_1 = stq_0_bits_addr_valid & ~stq_0_bits_addr_is_virtual & stq_0_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_423;
  wire [14:0] _write_mask_mask_T_2 = 15'h1 << stq_0_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_6 = 15'h3 << {12'h0, stq_0_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_0_bits_uop_mem_size)
      2'b00:
        casez_tmp_423 = _write_mask_mask_T_2[7:0];
      2'b01:
        casez_tmp_423 = _write_mask_mask_T_6[7:0];
      2'b10:
        casez_tmp_423 = stq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_423 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1080 = do_ld_search_0 & stq_0_valid & lcam_st_dep_mask_0[0];
  wire [7:0]  _GEN_1081 = casez_tmp_387 & casez_tmp_423;
  wire        _GEN_1082 = _GEN_1081 == casez_tmp_387 & ~stq_0_bits_uop_is_fence & ~stq_0_bits_uop_is_amo & dword_addr_matches_32_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_32;
  wire        _GEN_1083 = (|_GEN_1081) & dword_addr_matches_32_0;
  reg         io_dmem_s1_kill_0_REG_33;
  wire        _GEN_1084 = stq_0_bits_uop_is_fence | stq_0_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_34;
  wire        _GEN_1085 = _GEN_1080 ? (_GEN_1082 ? io_dmem_s1_kill_0_REG_32 : _GEN_1083 ? io_dmem_s1_kill_0_REG_33 : _GEN_1084 ? io_dmem_s1_kill_0_REG_34 : _GEN_1069) : _GEN_1069;
  wire        _GEN_1086 = do_ld_search_1 & stq_0_valid & lcam_st_dep_mask_1[0];
  wire [7:0]  _GEN_1087 = casez_tmp_388 & casez_tmp_423;
  wire        _GEN_1088 = _GEN_1087 == casez_tmp_388 & ~stq_0_bits_uop_is_fence & ~stq_0_bits_uop_is_amo & dword_addr_matches_32_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_32;
  wire        _GEN_1089 = (|_GEN_1087) & dword_addr_matches_32_1;
  reg         io_dmem_s1_kill_1_REG_33;
  reg         io_dmem_s1_kill_1_REG_34;
  wire        _GEN_1090 = _GEN_1086 ? (_GEN_1088 ? io_dmem_s1_kill_1_REG_32 : _GEN_1089 ? io_dmem_s1_kill_1_REG_33 : _GEN_1084 ? io_dmem_s1_kill_1_REG_34 : _GEN_1079) : _GEN_1079;
  wire        dword_addr_matches_33_0 = stq_1_bits_addr_valid & ~stq_1_bits_addr_is_virtual & stq_1_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_33_1 = stq_1_bits_addr_valid & ~stq_1_bits_addr_is_virtual & stq_1_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_424;
  wire [14:0] _write_mask_mask_T_17 = 15'h1 << stq_1_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_21 = 15'h3 << {12'h0, stq_1_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_1_bits_uop_mem_size)
      2'b00:
        casez_tmp_424 = _write_mask_mask_T_17[7:0];
      2'b01:
        casez_tmp_424 = _write_mask_mask_T_21[7:0];
      2'b10:
        casez_tmp_424 = stq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_424 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1091 = do_ld_search_0 & stq_1_valid & lcam_st_dep_mask_0[1];
  wire [7:0]  _GEN_1092 = casez_tmp_387 & casez_tmp_424;
  wire        _GEN_1093 = _GEN_1092 == casez_tmp_387 & ~stq_1_bits_uop_is_fence & ~stq_1_bits_uop_is_amo & dword_addr_matches_33_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_35;
  wire        _GEN_1094 = (|_GEN_1092) & dword_addr_matches_33_0;
  reg         io_dmem_s1_kill_0_REG_36;
  wire        _GEN_1095 = stq_1_bits_uop_is_fence | stq_1_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_37;
  wire        _GEN_1096 = _GEN_1091 ? (_GEN_1093 ? io_dmem_s1_kill_0_REG_35 : _GEN_1094 ? io_dmem_s1_kill_0_REG_36 : _GEN_1095 ? io_dmem_s1_kill_0_REG_37 : _GEN_1085) : _GEN_1085;
  wire        _GEN_1097 = do_ld_search_1 & stq_1_valid & lcam_st_dep_mask_1[1];
  wire [7:0]  _GEN_1098 = casez_tmp_388 & casez_tmp_424;
  wire        _GEN_1099 = _GEN_1098 == casez_tmp_388 & ~stq_1_bits_uop_is_fence & ~stq_1_bits_uop_is_amo & dword_addr_matches_33_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_35;
  wire        _GEN_1100 = (|_GEN_1098) & dword_addr_matches_33_1;
  reg         io_dmem_s1_kill_1_REG_36;
  reg         io_dmem_s1_kill_1_REG_37;
  wire        _GEN_1101 = _GEN_1097 ? (_GEN_1099 ? io_dmem_s1_kill_1_REG_35 : _GEN_1100 ? io_dmem_s1_kill_1_REG_36 : _GEN_1095 ? io_dmem_s1_kill_1_REG_37 : _GEN_1090) : _GEN_1090;
  wire        dword_addr_matches_34_0 = stq_2_bits_addr_valid & ~stq_2_bits_addr_is_virtual & stq_2_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_34_1 = stq_2_bits_addr_valid & ~stq_2_bits_addr_is_virtual & stq_2_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_425;
  wire [14:0] _write_mask_mask_T_32 = 15'h1 << stq_2_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_36 = 15'h3 << {12'h0, stq_2_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_2_bits_uop_mem_size)
      2'b00:
        casez_tmp_425 = _write_mask_mask_T_32[7:0];
      2'b01:
        casez_tmp_425 = _write_mask_mask_T_36[7:0];
      2'b10:
        casez_tmp_425 = stq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_425 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1102 = do_ld_search_0 & stq_2_valid & lcam_st_dep_mask_0[2];
  wire [7:0]  _GEN_1103 = casez_tmp_387 & casez_tmp_425;
  wire        _GEN_1104 = _GEN_1103 == casez_tmp_387 & ~stq_2_bits_uop_is_fence & ~stq_2_bits_uop_is_amo & dword_addr_matches_34_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_38;
  wire        _GEN_1105 = (|_GEN_1103) & dword_addr_matches_34_0;
  reg         io_dmem_s1_kill_0_REG_39;
  wire        _GEN_1106 = stq_2_bits_uop_is_fence | stq_2_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_40;
  wire        _GEN_1107 = _GEN_1102 ? (_GEN_1104 ? io_dmem_s1_kill_0_REG_38 : _GEN_1105 ? io_dmem_s1_kill_0_REG_39 : _GEN_1106 ? io_dmem_s1_kill_0_REG_40 : _GEN_1096) : _GEN_1096;
  wire        _GEN_1108 = do_ld_search_1 & stq_2_valid & lcam_st_dep_mask_1[2];
  wire [7:0]  _GEN_1109 = casez_tmp_388 & casez_tmp_425;
  wire        _GEN_1110 = _GEN_1109 == casez_tmp_388 & ~stq_2_bits_uop_is_fence & ~stq_2_bits_uop_is_amo & dword_addr_matches_34_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_38;
  wire        _GEN_1111 = (|_GEN_1109) & dword_addr_matches_34_1;
  reg         io_dmem_s1_kill_1_REG_39;
  reg         io_dmem_s1_kill_1_REG_40;
  wire        _GEN_1112 = _GEN_1108 ? (_GEN_1110 ? io_dmem_s1_kill_1_REG_38 : _GEN_1111 ? io_dmem_s1_kill_1_REG_39 : _GEN_1106 ? io_dmem_s1_kill_1_REG_40 : _GEN_1101) : _GEN_1101;
  wire        dword_addr_matches_35_0 = stq_3_bits_addr_valid & ~stq_3_bits_addr_is_virtual & stq_3_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_35_1 = stq_3_bits_addr_valid & ~stq_3_bits_addr_is_virtual & stq_3_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_426;
  wire [14:0] _write_mask_mask_T_47 = 15'h1 << stq_3_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_51 = 15'h3 << {12'h0, stq_3_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_3_bits_uop_mem_size)
      2'b00:
        casez_tmp_426 = _write_mask_mask_T_47[7:0];
      2'b01:
        casez_tmp_426 = _write_mask_mask_T_51[7:0];
      2'b10:
        casez_tmp_426 = stq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_426 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1113 = do_ld_search_0 & stq_3_valid & lcam_st_dep_mask_0[3];
  wire [7:0]  _GEN_1114 = casez_tmp_387 & casez_tmp_426;
  wire        _GEN_1115 = _GEN_1114 == casez_tmp_387 & ~stq_3_bits_uop_is_fence & ~stq_3_bits_uop_is_amo & dword_addr_matches_35_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_41;
  wire        _GEN_1116 = (|_GEN_1114) & dword_addr_matches_35_0;
  reg         io_dmem_s1_kill_0_REG_42;
  wire        _GEN_1117 = stq_3_bits_uop_is_fence | stq_3_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_43;
  wire        _GEN_1118 = _GEN_1113 ? (_GEN_1115 ? io_dmem_s1_kill_0_REG_41 : _GEN_1116 ? io_dmem_s1_kill_0_REG_42 : _GEN_1117 ? io_dmem_s1_kill_0_REG_43 : _GEN_1107) : _GEN_1107;
  wire        _GEN_1119 = do_ld_search_1 & stq_3_valid & lcam_st_dep_mask_1[3];
  wire [7:0]  _GEN_1120 = casez_tmp_388 & casez_tmp_426;
  wire        _GEN_1121 = _GEN_1120 == casez_tmp_388 & ~stq_3_bits_uop_is_fence & ~stq_3_bits_uop_is_amo & dword_addr_matches_35_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_41;
  wire        _GEN_1122 = (|_GEN_1120) & dword_addr_matches_35_1;
  reg         io_dmem_s1_kill_1_REG_42;
  reg         io_dmem_s1_kill_1_REG_43;
  wire        _GEN_1123 = _GEN_1119 ? (_GEN_1121 ? io_dmem_s1_kill_1_REG_41 : _GEN_1122 ? io_dmem_s1_kill_1_REG_42 : _GEN_1117 ? io_dmem_s1_kill_1_REG_43 : _GEN_1112) : _GEN_1112;
  wire        dword_addr_matches_36_0 = stq_4_bits_addr_valid & ~stq_4_bits_addr_is_virtual & stq_4_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_36_1 = stq_4_bits_addr_valid & ~stq_4_bits_addr_is_virtual & stq_4_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_427;
  wire [14:0] _write_mask_mask_T_62 = 15'h1 << stq_4_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_66 = 15'h3 << {12'h0, stq_4_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_4_bits_uop_mem_size)
      2'b00:
        casez_tmp_427 = _write_mask_mask_T_62[7:0];
      2'b01:
        casez_tmp_427 = _write_mask_mask_T_66[7:0];
      2'b10:
        casez_tmp_427 = stq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_427 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1124 = do_ld_search_0 & stq_4_valid & lcam_st_dep_mask_0[4];
  wire [7:0]  _GEN_1125 = casez_tmp_387 & casez_tmp_427;
  wire        _GEN_1126 = _GEN_1125 == casez_tmp_387 & ~stq_4_bits_uop_is_fence & ~stq_4_bits_uop_is_amo & dword_addr_matches_36_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_44;
  wire        _GEN_1127 = (|_GEN_1125) & dword_addr_matches_36_0;
  reg         io_dmem_s1_kill_0_REG_45;
  wire        _GEN_1128 = stq_4_bits_uop_is_fence | stq_4_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_46;
  wire        _GEN_1129 = _GEN_1124 ? (_GEN_1126 ? io_dmem_s1_kill_0_REG_44 : _GEN_1127 ? io_dmem_s1_kill_0_REG_45 : _GEN_1128 ? io_dmem_s1_kill_0_REG_46 : _GEN_1118) : _GEN_1118;
  wire        _GEN_1130 = do_ld_search_1 & stq_4_valid & lcam_st_dep_mask_1[4];
  wire [7:0]  _GEN_1131 = casez_tmp_388 & casez_tmp_427;
  wire        _GEN_1132 = _GEN_1131 == casez_tmp_388 & ~stq_4_bits_uop_is_fence & ~stq_4_bits_uop_is_amo & dword_addr_matches_36_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_44;
  wire        _GEN_1133 = (|_GEN_1131) & dword_addr_matches_36_1;
  reg         io_dmem_s1_kill_1_REG_45;
  reg         io_dmem_s1_kill_1_REG_46;
  wire        _GEN_1134 = _GEN_1130 ? (_GEN_1132 ? io_dmem_s1_kill_1_REG_44 : _GEN_1133 ? io_dmem_s1_kill_1_REG_45 : _GEN_1128 ? io_dmem_s1_kill_1_REG_46 : _GEN_1123) : _GEN_1123;
  wire        dword_addr_matches_37_0 = stq_5_bits_addr_valid & ~stq_5_bits_addr_is_virtual & stq_5_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_37_1 = stq_5_bits_addr_valid & ~stq_5_bits_addr_is_virtual & stq_5_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_428;
  wire [14:0] _write_mask_mask_T_77 = 15'h1 << stq_5_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_81 = 15'h3 << {12'h0, stq_5_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_5_bits_uop_mem_size)
      2'b00:
        casez_tmp_428 = _write_mask_mask_T_77[7:0];
      2'b01:
        casez_tmp_428 = _write_mask_mask_T_81[7:0];
      2'b10:
        casez_tmp_428 = stq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_428 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1135 = do_ld_search_0 & stq_5_valid & lcam_st_dep_mask_0[5];
  wire [7:0]  _GEN_1136 = casez_tmp_387 & casez_tmp_428;
  wire        _GEN_1137 = _GEN_1136 == casez_tmp_387 & ~stq_5_bits_uop_is_fence & ~stq_5_bits_uop_is_amo & dword_addr_matches_37_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_47;
  wire        _GEN_1138 = (|_GEN_1136) & dword_addr_matches_37_0;
  reg         io_dmem_s1_kill_0_REG_48;
  wire        _GEN_1139 = stq_5_bits_uop_is_fence | stq_5_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_49;
  wire        _GEN_1140 = _GEN_1135 ? (_GEN_1137 ? io_dmem_s1_kill_0_REG_47 : _GEN_1138 ? io_dmem_s1_kill_0_REG_48 : _GEN_1139 ? io_dmem_s1_kill_0_REG_49 : _GEN_1129) : _GEN_1129;
  wire        _GEN_1141 = do_ld_search_1 & stq_5_valid & lcam_st_dep_mask_1[5];
  wire [7:0]  _GEN_1142 = casez_tmp_388 & casez_tmp_428;
  wire        _GEN_1143 = _GEN_1142 == casez_tmp_388 & ~stq_5_bits_uop_is_fence & ~stq_5_bits_uop_is_amo & dword_addr_matches_37_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_47;
  wire        _GEN_1144 = (|_GEN_1142) & dword_addr_matches_37_1;
  reg         io_dmem_s1_kill_1_REG_48;
  reg         io_dmem_s1_kill_1_REG_49;
  wire        _GEN_1145 = _GEN_1141 ? (_GEN_1143 ? io_dmem_s1_kill_1_REG_47 : _GEN_1144 ? io_dmem_s1_kill_1_REG_48 : _GEN_1139 ? io_dmem_s1_kill_1_REG_49 : _GEN_1134) : _GEN_1134;
  wire        dword_addr_matches_38_0 = stq_6_bits_addr_valid & ~stq_6_bits_addr_is_virtual & stq_6_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_38_1 = stq_6_bits_addr_valid & ~stq_6_bits_addr_is_virtual & stq_6_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_429;
  wire [14:0] _write_mask_mask_T_92 = 15'h1 << stq_6_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_96 = 15'h3 << {12'h0, stq_6_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_6_bits_uop_mem_size)
      2'b00:
        casez_tmp_429 = _write_mask_mask_T_92[7:0];
      2'b01:
        casez_tmp_429 = _write_mask_mask_T_96[7:0];
      2'b10:
        casez_tmp_429 = stq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_429 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1146 = do_ld_search_0 & stq_6_valid & lcam_st_dep_mask_0[6];
  wire [7:0]  _GEN_1147 = casez_tmp_387 & casez_tmp_429;
  wire        _GEN_1148 = _GEN_1147 == casez_tmp_387 & ~stq_6_bits_uop_is_fence & ~stq_6_bits_uop_is_amo & dword_addr_matches_38_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_50;
  wire        _GEN_1149 = (|_GEN_1147) & dword_addr_matches_38_0;
  reg         io_dmem_s1_kill_0_REG_51;
  wire        _GEN_1150 = stq_6_bits_uop_is_fence | stq_6_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_52;
  wire        _GEN_1151 = _GEN_1146 ? (_GEN_1148 ? io_dmem_s1_kill_0_REG_50 : _GEN_1149 ? io_dmem_s1_kill_0_REG_51 : _GEN_1150 ? io_dmem_s1_kill_0_REG_52 : _GEN_1140) : _GEN_1140;
  wire        _GEN_1152 = do_ld_search_1 & stq_6_valid & lcam_st_dep_mask_1[6];
  wire [7:0]  _GEN_1153 = casez_tmp_388 & casez_tmp_429;
  wire        _GEN_1154 = _GEN_1153 == casez_tmp_388 & ~stq_6_bits_uop_is_fence & ~stq_6_bits_uop_is_amo & dword_addr_matches_38_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_50;
  wire        _GEN_1155 = (|_GEN_1153) & dword_addr_matches_38_1;
  reg         io_dmem_s1_kill_1_REG_51;
  reg         io_dmem_s1_kill_1_REG_52;
  wire        _GEN_1156 = _GEN_1152 ? (_GEN_1154 ? io_dmem_s1_kill_1_REG_50 : _GEN_1155 ? io_dmem_s1_kill_1_REG_51 : _GEN_1150 ? io_dmem_s1_kill_1_REG_52 : _GEN_1145) : _GEN_1145;
  wire        dword_addr_matches_39_0 = stq_7_bits_addr_valid & ~stq_7_bits_addr_is_virtual & stq_7_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_39_1 = stq_7_bits_addr_valid & ~stq_7_bits_addr_is_virtual & stq_7_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_430;
  wire [14:0] _write_mask_mask_T_107 = 15'h1 << stq_7_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_111 = 15'h3 << {12'h0, stq_7_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_7_bits_uop_mem_size)
      2'b00:
        casez_tmp_430 = _write_mask_mask_T_107[7:0];
      2'b01:
        casez_tmp_430 = _write_mask_mask_T_111[7:0];
      2'b10:
        casez_tmp_430 = stq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_430 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1157 = do_ld_search_0 & stq_7_valid & lcam_st_dep_mask_0[7];
  wire [7:0]  _GEN_1158 = casez_tmp_387 & casez_tmp_430;
  wire        _GEN_1159 = _GEN_1158 == casez_tmp_387 & ~stq_7_bits_uop_is_fence & ~stq_7_bits_uop_is_amo & dword_addr_matches_39_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_53;
  wire        _GEN_1160 = (|_GEN_1158) & dword_addr_matches_39_0;
  reg         io_dmem_s1_kill_0_REG_54;
  wire        _GEN_1161 = stq_7_bits_uop_is_fence | stq_7_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_55;
  wire        _GEN_1162 = _GEN_1157 ? (_GEN_1159 ? io_dmem_s1_kill_0_REG_53 : _GEN_1160 ? io_dmem_s1_kill_0_REG_54 : _GEN_1161 ? io_dmem_s1_kill_0_REG_55 : _GEN_1151) : _GEN_1151;
  wire        _GEN_1163 = do_ld_search_1 & stq_7_valid & lcam_st_dep_mask_1[7];
  wire [7:0]  _GEN_1164 = casez_tmp_388 & casez_tmp_430;
  wire        _GEN_1165 = _GEN_1164 == casez_tmp_388 & ~stq_7_bits_uop_is_fence & ~stq_7_bits_uop_is_amo & dword_addr_matches_39_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_53;
  wire        _GEN_1166 = (|_GEN_1164) & dword_addr_matches_39_1;
  reg         io_dmem_s1_kill_1_REG_54;
  reg         io_dmem_s1_kill_1_REG_55;
  wire        _GEN_1167 = _GEN_1163 ? (_GEN_1165 ? io_dmem_s1_kill_1_REG_53 : _GEN_1166 ? io_dmem_s1_kill_1_REG_54 : _GEN_1161 ? io_dmem_s1_kill_1_REG_55 : _GEN_1156) : _GEN_1156;
  wire        dword_addr_matches_40_0 = stq_8_bits_addr_valid & ~stq_8_bits_addr_is_virtual & stq_8_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_40_1 = stq_8_bits_addr_valid & ~stq_8_bits_addr_is_virtual & stq_8_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_431;
  wire [14:0] _write_mask_mask_T_122 = 15'h1 << stq_8_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_126 = 15'h3 << {12'h0, stq_8_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_8_bits_uop_mem_size)
      2'b00:
        casez_tmp_431 = _write_mask_mask_T_122[7:0];
      2'b01:
        casez_tmp_431 = _write_mask_mask_T_126[7:0];
      2'b10:
        casez_tmp_431 = stq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_431 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1168 = do_ld_search_0 & stq_8_valid & lcam_st_dep_mask_0[8];
  wire [7:0]  _GEN_1169 = casez_tmp_387 & casez_tmp_431;
  wire        _GEN_1170 = _GEN_1169 == casez_tmp_387 & ~stq_8_bits_uop_is_fence & ~stq_8_bits_uop_is_amo & dword_addr_matches_40_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_56;
  wire        _GEN_1171 = (|_GEN_1169) & dword_addr_matches_40_0;
  reg         io_dmem_s1_kill_0_REG_57;
  wire        _GEN_1172 = stq_8_bits_uop_is_fence | stq_8_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_58;
  wire        _GEN_1173 = _GEN_1168 ? (_GEN_1170 ? io_dmem_s1_kill_0_REG_56 : _GEN_1171 ? io_dmem_s1_kill_0_REG_57 : _GEN_1172 ? io_dmem_s1_kill_0_REG_58 : _GEN_1162) : _GEN_1162;
  wire        _GEN_1174 = do_ld_search_1 & stq_8_valid & lcam_st_dep_mask_1[8];
  wire [7:0]  _GEN_1175 = casez_tmp_388 & casez_tmp_431;
  wire        _GEN_1176 = _GEN_1175 == casez_tmp_388 & ~stq_8_bits_uop_is_fence & ~stq_8_bits_uop_is_amo & dword_addr_matches_40_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_56;
  wire        _GEN_1177 = (|_GEN_1175) & dword_addr_matches_40_1;
  reg         io_dmem_s1_kill_1_REG_57;
  reg         io_dmem_s1_kill_1_REG_58;
  wire        _GEN_1178 = _GEN_1174 ? (_GEN_1176 ? io_dmem_s1_kill_1_REG_56 : _GEN_1177 ? io_dmem_s1_kill_1_REG_57 : _GEN_1172 ? io_dmem_s1_kill_1_REG_58 : _GEN_1167) : _GEN_1167;
  wire        dword_addr_matches_41_0 = stq_9_bits_addr_valid & ~stq_9_bits_addr_is_virtual & stq_9_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_41_1 = stq_9_bits_addr_valid & ~stq_9_bits_addr_is_virtual & stq_9_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_432;
  wire [14:0] _write_mask_mask_T_137 = 15'h1 << stq_9_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_141 = 15'h3 << {12'h0, stq_9_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_9_bits_uop_mem_size)
      2'b00:
        casez_tmp_432 = _write_mask_mask_T_137[7:0];
      2'b01:
        casez_tmp_432 = _write_mask_mask_T_141[7:0];
      2'b10:
        casez_tmp_432 = stq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_432 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1179 = do_ld_search_0 & stq_9_valid & lcam_st_dep_mask_0[9];
  wire [7:0]  _GEN_1180 = casez_tmp_387 & casez_tmp_432;
  wire        _GEN_1181 = _GEN_1180 == casez_tmp_387 & ~stq_9_bits_uop_is_fence & ~stq_9_bits_uop_is_amo & dword_addr_matches_41_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_59;
  wire        _GEN_1182 = (|_GEN_1180) & dword_addr_matches_41_0;
  reg         io_dmem_s1_kill_0_REG_60;
  wire        _GEN_1183 = stq_9_bits_uop_is_fence | stq_9_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_61;
  wire        _GEN_1184 = _GEN_1179 ? (_GEN_1181 ? io_dmem_s1_kill_0_REG_59 : _GEN_1182 ? io_dmem_s1_kill_0_REG_60 : _GEN_1183 ? io_dmem_s1_kill_0_REG_61 : _GEN_1173) : _GEN_1173;
  wire        _GEN_1185 = do_ld_search_1 & stq_9_valid & lcam_st_dep_mask_1[9];
  wire [7:0]  _GEN_1186 = casez_tmp_388 & casez_tmp_432;
  wire        _GEN_1187 = _GEN_1186 == casez_tmp_388 & ~stq_9_bits_uop_is_fence & ~stq_9_bits_uop_is_amo & dword_addr_matches_41_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_59;
  wire        _GEN_1188 = (|_GEN_1186) & dword_addr_matches_41_1;
  reg         io_dmem_s1_kill_1_REG_60;
  reg         io_dmem_s1_kill_1_REG_61;
  wire        _GEN_1189 = _GEN_1185 ? (_GEN_1187 ? io_dmem_s1_kill_1_REG_59 : _GEN_1188 ? io_dmem_s1_kill_1_REG_60 : _GEN_1183 ? io_dmem_s1_kill_1_REG_61 : _GEN_1178) : _GEN_1178;
  wire        dword_addr_matches_42_0 = stq_10_bits_addr_valid & ~stq_10_bits_addr_is_virtual & stq_10_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_42_1 = stq_10_bits_addr_valid & ~stq_10_bits_addr_is_virtual & stq_10_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_433;
  wire [14:0] _write_mask_mask_T_152 = 15'h1 << stq_10_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_156 = 15'h3 << {12'h0, stq_10_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_10_bits_uop_mem_size)
      2'b00:
        casez_tmp_433 = _write_mask_mask_T_152[7:0];
      2'b01:
        casez_tmp_433 = _write_mask_mask_T_156[7:0];
      2'b10:
        casez_tmp_433 = stq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_433 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1190 = do_ld_search_0 & stq_10_valid & lcam_st_dep_mask_0[10];
  wire [7:0]  _GEN_1191 = casez_tmp_387 & casez_tmp_433;
  wire        _GEN_1192 = _GEN_1191 == casez_tmp_387 & ~stq_10_bits_uop_is_fence & ~stq_10_bits_uop_is_amo & dword_addr_matches_42_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_62;
  wire        _GEN_1193 = (|_GEN_1191) & dword_addr_matches_42_0;
  reg         io_dmem_s1_kill_0_REG_63;
  wire        _GEN_1194 = stq_10_bits_uop_is_fence | stq_10_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_64;
  wire        _GEN_1195 = _GEN_1190 ? (_GEN_1192 ? io_dmem_s1_kill_0_REG_62 : _GEN_1193 ? io_dmem_s1_kill_0_REG_63 : _GEN_1194 ? io_dmem_s1_kill_0_REG_64 : _GEN_1184) : _GEN_1184;
  wire        _GEN_1196 = do_ld_search_1 & stq_10_valid & lcam_st_dep_mask_1[10];
  wire [7:0]  _GEN_1197 = casez_tmp_388 & casez_tmp_433;
  wire        _GEN_1198 = _GEN_1197 == casez_tmp_388 & ~stq_10_bits_uop_is_fence & ~stq_10_bits_uop_is_amo & dword_addr_matches_42_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_62;
  wire        _GEN_1199 = (|_GEN_1197) & dword_addr_matches_42_1;
  reg         io_dmem_s1_kill_1_REG_63;
  reg         io_dmem_s1_kill_1_REG_64;
  wire        _GEN_1200 = _GEN_1196 ? (_GEN_1198 ? io_dmem_s1_kill_1_REG_62 : _GEN_1199 ? io_dmem_s1_kill_1_REG_63 : _GEN_1194 ? io_dmem_s1_kill_1_REG_64 : _GEN_1189) : _GEN_1189;
  wire        dword_addr_matches_43_0 = stq_11_bits_addr_valid & ~stq_11_bits_addr_is_virtual & stq_11_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_43_1 = stq_11_bits_addr_valid & ~stq_11_bits_addr_is_virtual & stq_11_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_434;
  wire [14:0] _write_mask_mask_T_167 = 15'h1 << stq_11_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_171 = 15'h3 << {12'h0, stq_11_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_11_bits_uop_mem_size)
      2'b00:
        casez_tmp_434 = _write_mask_mask_T_167[7:0];
      2'b01:
        casez_tmp_434 = _write_mask_mask_T_171[7:0];
      2'b10:
        casez_tmp_434 = stq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_434 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1201 = do_ld_search_0 & stq_11_valid & lcam_st_dep_mask_0[11];
  wire [7:0]  _GEN_1202 = casez_tmp_387 & casez_tmp_434;
  wire        _GEN_1203 = _GEN_1202 == casez_tmp_387 & ~stq_11_bits_uop_is_fence & ~stq_11_bits_uop_is_amo & dword_addr_matches_43_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_65;
  wire        _GEN_1204 = (|_GEN_1202) & dword_addr_matches_43_0;
  reg         io_dmem_s1_kill_0_REG_66;
  wire        _GEN_1205 = stq_11_bits_uop_is_fence | stq_11_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_67;
  wire        _GEN_1206 = _GEN_1201 ? (_GEN_1203 ? io_dmem_s1_kill_0_REG_65 : _GEN_1204 ? io_dmem_s1_kill_0_REG_66 : _GEN_1205 ? io_dmem_s1_kill_0_REG_67 : _GEN_1195) : _GEN_1195;
  wire        _GEN_1207 = do_ld_search_1 & stq_11_valid & lcam_st_dep_mask_1[11];
  wire [7:0]  _GEN_1208 = casez_tmp_388 & casez_tmp_434;
  wire        _GEN_1209 = _GEN_1208 == casez_tmp_388 & ~stq_11_bits_uop_is_fence & ~stq_11_bits_uop_is_amo & dword_addr_matches_43_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_65;
  wire        _GEN_1210 = (|_GEN_1208) & dword_addr_matches_43_1;
  reg         io_dmem_s1_kill_1_REG_66;
  reg         io_dmem_s1_kill_1_REG_67;
  wire        _GEN_1211 = _GEN_1207 ? (_GEN_1209 ? io_dmem_s1_kill_1_REG_65 : _GEN_1210 ? io_dmem_s1_kill_1_REG_66 : _GEN_1205 ? io_dmem_s1_kill_1_REG_67 : _GEN_1200) : _GEN_1200;
  wire        dword_addr_matches_44_0 = stq_12_bits_addr_valid & ~stq_12_bits_addr_is_virtual & stq_12_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_44_1 = stq_12_bits_addr_valid & ~stq_12_bits_addr_is_virtual & stq_12_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_435;
  wire [14:0] _write_mask_mask_T_182 = 15'h1 << stq_12_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_186 = 15'h3 << {12'h0, stq_12_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_12_bits_uop_mem_size)
      2'b00:
        casez_tmp_435 = _write_mask_mask_T_182[7:0];
      2'b01:
        casez_tmp_435 = _write_mask_mask_T_186[7:0];
      2'b10:
        casez_tmp_435 = stq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_435 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1212 = do_ld_search_0 & stq_12_valid & lcam_st_dep_mask_0[12];
  wire [7:0]  _GEN_1213 = casez_tmp_387 & casez_tmp_435;
  wire        _GEN_1214 = _GEN_1213 == casez_tmp_387 & ~stq_12_bits_uop_is_fence & ~stq_12_bits_uop_is_amo & dword_addr_matches_44_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_68;
  wire        _GEN_1215 = (|_GEN_1213) & dword_addr_matches_44_0;
  reg         io_dmem_s1_kill_0_REG_69;
  wire        _GEN_1216 = stq_12_bits_uop_is_fence | stq_12_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_70;
  wire        _GEN_1217 = _GEN_1212 ? (_GEN_1214 ? io_dmem_s1_kill_0_REG_68 : _GEN_1215 ? io_dmem_s1_kill_0_REG_69 : _GEN_1216 ? io_dmem_s1_kill_0_REG_70 : _GEN_1206) : _GEN_1206;
  wire        _GEN_1218 = do_ld_search_1 & stq_12_valid & lcam_st_dep_mask_1[12];
  wire [7:0]  _GEN_1219 = casez_tmp_388 & casez_tmp_435;
  wire        _GEN_1220 = _GEN_1219 == casez_tmp_388 & ~stq_12_bits_uop_is_fence & ~stq_12_bits_uop_is_amo & dword_addr_matches_44_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_68;
  wire        _GEN_1221 = (|_GEN_1219) & dword_addr_matches_44_1;
  reg         io_dmem_s1_kill_1_REG_69;
  reg         io_dmem_s1_kill_1_REG_70;
  wire        _GEN_1222 = _GEN_1218 ? (_GEN_1220 ? io_dmem_s1_kill_1_REG_68 : _GEN_1221 ? io_dmem_s1_kill_1_REG_69 : _GEN_1216 ? io_dmem_s1_kill_1_REG_70 : _GEN_1211) : _GEN_1211;
  wire        dword_addr_matches_45_0 = stq_13_bits_addr_valid & ~stq_13_bits_addr_is_virtual & stq_13_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_45_1 = stq_13_bits_addr_valid & ~stq_13_bits_addr_is_virtual & stq_13_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_436;
  wire [14:0] _write_mask_mask_T_197 = 15'h1 << stq_13_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_201 = 15'h3 << {12'h0, stq_13_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_13_bits_uop_mem_size)
      2'b00:
        casez_tmp_436 = _write_mask_mask_T_197[7:0];
      2'b01:
        casez_tmp_436 = _write_mask_mask_T_201[7:0];
      2'b10:
        casez_tmp_436 = stq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_436 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1223 = do_ld_search_0 & stq_13_valid & lcam_st_dep_mask_0[13];
  wire [7:0]  _GEN_1224 = casez_tmp_387 & casez_tmp_436;
  wire        _GEN_1225 = _GEN_1224 == casez_tmp_387 & ~stq_13_bits_uop_is_fence & ~stq_13_bits_uop_is_amo & dword_addr_matches_45_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_71;
  wire        _GEN_1226 = (|_GEN_1224) & dword_addr_matches_45_0;
  reg         io_dmem_s1_kill_0_REG_72;
  wire        _GEN_1227 = stq_13_bits_uop_is_fence | stq_13_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_73;
  wire        _GEN_1228 = _GEN_1223 ? (_GEN_1225 ? io_dmem_s1_kill_0_REG_71 : _GEN_1226 ? io_dmem_s1_kill_0_REG_72 : _GEN_1227 ? io_dmem_s1_kill_0_REG_73 : _GEN_1217) : _GEN_1217;
  wire        _GEN_1229 = do_ld_search_1 & stq_13_valid & lcam_st_dep_mask_1[13];
  wire [7:0]  _GEN_1230 = casez_tmp_388 & casez_tmp_436;
  wire        _GEN_1231 = _GEN_1230 == casez_tmp_388 & ~stq_13_bits_uop_is_fence & ~stq_13_bits_uop_is_amo & dword_addr_matches_45_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_71;
  wire        _GEN_1232 = (|_GEN_1230) & dword_addr_matches_45_1;
  reg         io_dmem_s1_kill_1_REG_72;
  reg         io_dmem_s1_kill_1_REG_73;
  wire        _GEN_1233 = _GEN_1229 ? (_GEN_1231 ? io_dmem_s1_kill_1_REG_71 : _GEN_1232 ? io_dmem_s1_kill_1_REG_72 : _GEN_1227 ? io_dmem_s1_kill_1_REG_73 : _GEN_1222) : _GEN_1222;
  wire        dword_addr_matches_46_0 = stq_14_bits_addr_valid & ~stq_14_bits_addr_is_virtual & stq_14_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_46_1 = stq_14_bits_addr_valid & ~stq_14_bits_addr_is_virtual & stq_14_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_437;
  wire [14:0] _write_mask_mask_T_212 = 15'h1 << stq_14_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_216 = 15'h3 << {12'h0, stq_14_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_14_bits_uop_mem_size)
      2'b00:
        casez_tmp_437 = _write_mask_mask_T_212[7:0];
      2'b01:
        casez_tmp_437 = _write_mask_mask_T_216[7:0];
      2'b10:
        casez_tmp_437 = stq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_437 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1234 = do_ld_search_0 & stq_14_valid & lcam_st_dep_mask_0[14];
  wire [7:0]  _GEN_1235 = casez_tmp_387 & casez_tmp_437;
  wire        _GEN_1236 = _GEN_1235 == casez_tmp_387 & ~stq_14_bits_uop_is_fence & ~stq_14_bits_uop_is_amo & dword_addr_matches_46_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_74;
  wire        _GEN_1237 = (|_GEN_1235) & dword_addr_matches_46_0;
  reg         io_dmem_s1_kill_0_REG_75;
  wire        _GEN_1238 = stq_14_bits_uop_is_fence | stq_14_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_76;
  wire        _GEN_1239 = _GEN_1234 ? (_GEN_1236 ? io_dmem_s1_kill_0_REG_74 : _GEN_1237 ? io_dmem_s1_kill_0_REG_75 : _GEN_1238 ? io_dmem_s1_kill_0_REG_76 : _GEN_1228) : _GEN_1228;
  wire        _GEN_1240 = do_ld_search_1 & stq_14_valid & lcam_st_dep_mask_1[14];
  wire [7:0]  _GEN_1241 = casez_tmp_388 & casez_tmp_437;
  wire        _GEN_1242 = _GEN_1241 == casez_tmp_388 & ~stq_14_bits_uop_is_fence & ~stq_14_bits_uop_is_amo & dword_addr_matches_46_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_74;
  wire        _GEN_1243 = (|_GEN_1241) & dword_addr_matches_46_1;
  reg         io_dmem_s1_kill_1_REG_75;
  reg         io_dmem_s1_kill_1_REG_76;
  wire        _GEN_1244 = _GEN_1240 ? (_GEN_1242 ? io_dmem_s1_kill_1_REG_74 : _GEN_1243 ? io_dmem_s1_kill_1_REG_75 : _GEN_1238 ? io_dmem_s1_kill_1_REG_76 : _GEN_1233) : _GEN_1233;
  wire        dword_addr_matches_47_0 = stq_15_bits_addr_valid & ~stq_15_bits_addr_is_virtual & stq_15_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_47_1 = stq_15_bits_addr_valid & ~stq_15_bits_addr_is_virtual & stq_15_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_438;
  wire [14:0] _write_mask_mask_T_227 = 15'h1 << stq_15_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_231 = 15'h3 << {12'h0, stq_15_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_15_bits_uop_mem_size)
      2'b00:
        casez_tmp_438 = _write_mask_mask_T_227[7:0];
      2'b01:
        casez_tmp_438 = _write_mask_mask_T_231[7:0];
      2'b10:
        casez_tmp_438 = stq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_438 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1245 = do_ld_search_0 & stq_15_valid & lcam_st_dep_mask_0[15];
  wire [7:0]  _GEN_1246 = casez_tmp_387 & casez_tmp_438;
  wire        _GEN_1247 = _GEN_1246 == casez_tmp_387 & ~stq_15_bits_uop_is_fence & ~stq_15_bits_uop_is_amo & dword_addr_matches_47_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_77;
  wire        _GEN_1248 = (|_GEN_1246) & dword_addr_matches_47_0;
  reg         io_dmem_s1_kill_0_REG_78;
  wire        _GEN_1249 = stq_15_bits_uop_is_fence | stq_15_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_79;
  wire        _GEN_1250 = _GEN_1245 ? (_GEN_1247 ? io_dmem_s1_kill_0_REG_77 : _GEN_1248 ? io_dmem_s1_kill_0_REG_78 : _GEN_1249 ? io_dmem_s1_kill_0_REG_79 : _GEN_1239) : _GEN_1239;
  wire        _GEN_1251 = do_ld_search_1 & stq_15_valid & lcam_st_dep_mask_1[15];
  wire [7:0]  _GEN_1252 = casez_tmp_388 & casez_tmp_438;
  wire        _GEN_1253 = _GEN_1252 == casez_tmp_388 & ~stq_15_bits_uop_is_fence & ~stq_15_bits_uop_is_amo & dword_addr_matches_47_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_77;
  wire        _GEN_1254 = (|_GEN_1252) & dword_addr_matches_47_1;
  reg         io_dmem_s1_kill_1_REG_78;
  reg         io_dmem_s1_kill_1_REG_79;
  wire        _GEN_1255 = _GEN_1251 ? (_GEN_1253 ? io_dmem_s1_kill_1_REG_77 : _GEN_1254 ? io_dmem_s1_kill_1_REG_78 : _GEN_1249 ? io_dmem_s1_kill_1_REG_79 : _GEN_1244) : _GEN_1244;
  wire        dword_addr_matches_48_0 = stq_16_bits_addr_valid & ~stq_16_bits_addr_is_virtual & stq_16_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_48_1 = stq_16_bits_addr_valid & ~stq_16_bits_addr_is_virtual & stq_16_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_439;
  wire [14:0] _write_mask_mask_T_242 = 15'h1 << stq_16_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_246 = 15'h3 << {12'h0, stq_16_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_16_bits_uop_mem_size)
      2'b00:
        casez_tmp_439 = _write_mask_mask_T_242[7:0];
      2'b01:
        casez_tmp_439 = _write_mask_mask_T_246[7:0];
      2'b10:
        casez_tmp_439 = stq_16_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_439 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1256 = do_ld_search_0 & stq_16_valid & lcam_st_dep_mask_0[16];
  wire [7:0]  _GEN_1257 = casez_tmp_387 & casez_tmp_439;
  wire        _GEN_1258 = _GEN_1257 == casez_tmp_387 & ~stq_16_bits_uop_is_fence & ~stq_16_bits_uop_is_amo & dword_addr_matches_48_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_80;
  wire        _GEN_1259 = (|_GEN_1257) & dword_addr_matches_48_0;
  reg         io_dmem_s1_kill_0_REG_81;
  wire        _GEN_1260 = stq_16_bits_uop_is_fence | stq_16_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_82;
  wire        _GEN_1261 = _GEN_1256 ? (_GEN_1258 ? io_dmem_s1_kill_0_REG_80 : _GEN_1259 ? io_dmem_s1_kill_0_REG_81 : _GEN_1260 ? io_dmem_s1_kill_0_REG_82 : _GEN_1250) : _GEN_1250;
  wire        _GEN_1262 = do_ld_search_1 & stq_16_valid & lcam_st_dep_mask_1[16];
  wire [7:0]  _GEN_1263 = casez_tmp_388 & casez_tmp_439;
  wire        _GEN_1264 = _GEN_1263 == casez_tmp_388 & ~stq_16_bits_uop_is_fence & ~stq_16_bits_uop_is_amo & dword_addr_matches_48_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_80;
  wire        _GEN_1265 = (|_GEN_1263) & dword_addr_matches_48_1;
  reg         io_dmem_s1_kill_1_REG_81;
  reg         io_dmem_s1_kill_1_REG_82;
  wire        _GEN_1266 = _GEN_1262 ? (_GEN_1264 ? io_dmem_s1_kill_1_REG_80 : _GEN_1265 ? io_dmem_s1_kill_1_REG_81 : _GEN_1260 ? io_dmem_s1_kill_1_REG_82 : _GEN_1255) : _GEN_1255;
  wire        dword_addr_matches_49_0 = stq_17_bits_addr_valid & ~stq_17_bits_addr_is_virtual & stq_17_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_49_1 = stq_17_bits_addr_valid & ~stq_17_bits_addr_is_virtual & stq_17_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_440;
  wire [14:0] _write_mask_mask_T_257 = 15'h1 << stq_17_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_261 = 15'h3 << {12'h0, stq_17_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_17_bits_uop_mem_size)
      2'b00:
        casez_tmp_440 = _write_mask_mask_T_257[7:0];
      2'b01:
        casez_tmp_440 = _write_mask_mask_T_261[7:0];
      2'b10:
        casez_tmp_440 = stq_17_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_440 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1267 = do_ld_search_0 & stq_17_valid & lcam_st_dep_mask_0[17];
  wire [7:0]  _GEN_1268 = casez_tmp_387 & casez_tmp_440;
  wire        _GEN_1269 = _GEN_1268 == casez_tmp_387 & ~stq_17_bits_uop_is_fence & ~stq_17_bits_uop_is_amo & dword_addr_matches_49_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_83;
  wire        _GEN_1270 = (|_GEN_1268) & dword_addr_matches_49_0;
  reg         io_dmem_s1_kill_0_REG_84;
  wire        _GEN_1271 = stq_17_bits_uop_is_fence | stq_17_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_85;
  wire        _GEN_1272 = _GEN_1267 ? (_GEN_1269 ? io_dmem_s1_kill_0_REG_83 : _GEN_1270 ? io_dmem_s1_kill_0_REG_84 : _GEN_1271 ? io_dmem_s1_kill_0_REG_85 : _GEN_1261) : _GEN_1261;
  wire        _GEN_1273 = do_ld_search_1 & stq_17_valid & lcam_st_dep_mask_1[17];
  wire [7:0]  _GEN_1274 = casez_tmp_388 & casez_tmp_440;
  wire        _GEN_1275 = _GEN_1274 == casez_tmp_388 & ~stq_17_bits_uop_is_fence & ~stq_17_bits_uop_is_amo & dword_addr_matches_49_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_83;
  wire        _GEN_1276 = (|_GEN_1274) & dword_addr_matches_49_1;
  reg         io_dmem_s1_kill_1_REG_84;
  reg         io_dmem_s1_kill_1_REG_85;
  wire        _GEN_1277 = _GEN_1273 ? (_GEN_1275 ? io_dmem_s1_kill_1_REG_83 : _GEN_1276 ? io_dmem_s1_kill_1_REG_84 : _GEN_1271 ? io_dmem_s1_kill_1_REG_85 : _GEN_1266) : _GEN_1266;
  wire        dword_addr_matches_50_0 = stq_18_bits_addr_valid & ~stq_18_bits_addr_is_virtual & stq_18_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_50_1 = stq_18_bits_addr_valid & ~stq_18_bits_addr_is_virtual & stq_18_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_441;
  wire [14:0] _write_mask_mask_T_272 = 15'h1 << stq_18_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_276 = 15'h3 << {12'h0, stq_18_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_18_bits_uop_mem_size)
      2'b00:
        casez_tmp_441 = _write_mask_mask_T_272[7:0];
      2'b01:
        casez_tmp_441 = _write_mask_mask_T_276[7:0];
      2'b10:
        casez_tmp_441 = stq_18_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_441 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1278 = do_ld_search_0 & stq_18_valid & lcam_st_dep_mask_0[18];
  wire [7:0]  _GEN_1279 = casez_tmp_387 & casez_tmp_441;
  wire        _GEN_1280 = _GEN_1279 == casez_tmp_387 & ~stq_18_bits_uop_is_fence & ~stq_18_bits_uop_is_amo & dword_addr_matches_50_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_86;
  wire        _GEN_1281 = (|_GEN_1279) & dword_addr_matches_50_0;
  reg         io_dmem_s1_kill_0_REG_87;
  wire        _GEN_1282 = stq_18_bits_uop_is_fence | stq_18_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_88;
  wire        _GEN_1283 = _GEN_1278 ? (_GEN_1280 ? io_dmem_s1_kill_0_REG_86 : _GEN_1281 ? io_dmem_s1_kill_0_REG_87 : _GEN_1282 ? io_dmem_s1_kill_0_REG_88 : _GEN_1272) : _GEN_1272;
  wire        _GEN_1284 = do_ld_search_1 & stq_18_valid & lcam_st_dep_mask_1[18];
  wire [7:0]  _GEN_1285 = casez_tmp_388 & casez_tmp_441;
  wire        _GEN_1286 = _GEN_1285 == casez_tmp_388 & ~stq_18_bits_uop_is_fence & ~stq_18_bits_uop_is_amo & dword_addr_matches_50_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_86;
  wire        _GEN_1287 = (|_GEN_1285) & dword_addr_matches_50_1;
  reg         io_dmem_s1_kill_1_REG_87;
  reg         io_dmem_s1_kill_1_REG_88;
  wire        _GEN_1288 = _GEN_1284 ? (_GEN_1286 ? io_dmem_s1_kill_1_REG_86 : _GEN_1287 ? io_dmem_s1_kill_1_REG_87 : _GEN_1282 ? io_dmem_s1_kill_1_REG_88 : _GEN_1277) : _GEN_1277;
  wire        dword_addr_matches_51_0 = stq_19_bits_addr_valid & ~stq_19_bits_addr_is_virtual & stq_19_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_51_1 = stq_19_bits_addr_valid & ~stq_19_bits_addr_is_virtual & stq_19_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_442;
  wire [14:0] _write_mask_mask_T_287 = 15'h1 << stq_19_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_291 = 15'h3 << {12'h0, stq_19_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_19_bits_uop_mem_size)
      2'b00:
        casez_tmp_442 = _write_mask_mask_T_287[7:0];
      2'b01:
        casez_tmp_442 = _write_mask_mask_T_291[7:0];
      2'b10:
        casez_tmp_442 = stq_19_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_442 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1289 = do_ld_search_0 & stq_19_valid & lcam_st_dep_mask_0[19];
  wire [7:0]  _GEN_1290 = casez_tmp_387 & casez_tmp_442;
  wire        _GEN_1291 = _GEN_1290 == casez_tmp_387 & ~stq_19_bits_uop_is_fence & ~stq_19_bits_uop_is_amo & dword_addr_matches_51_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_89;
  wire        _GEN_1292 = (|_GEN_1290) & dword_addr_matches_51_0;
  reg         io_dmem_s1_kill_0_REG_90;
  wire        _GEN_1293 = stq_19_bits_uop_is_fence | stq_19_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_91;
  wire        _GEN_1294 = _GEN_1289 ? (_GEN_1291 ? io_dmem_s1_kill_0_REG_89 : _GEN_1292 ? io_dmem_s1_kill_0_REG_90 : _GEN_1293 ? io_dmem_s1_kill_0_REG_91 : _GEN_1283) : _GEN_1283;
  wire        _GEN_1295 = do_ld_search_1 & stq_19_valid & lcam_st_dep_mask_1[19];
  wire [7:0]  _GEN_1296 = casez_tmp_388 & casez_tmp_442;
  wire        _GEN_1297 = _GEN_1296 == casez_tmp_388 & ~stq_19_bits_uop_is_fence & ~stq_19_bits_uop_is_amo & dword_addr_matches_51_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_89;
  wire        _GEN_1298 = (|_GEN_1296) & dword_addr_matches_51_1;
  reg         io_dmem_s1_kill_1_REG_90;
  reg         io_dmem_s1_kill_1_REG_91;
  wire        _GEN_1299 = _GEN_1295 ? (_GEN_1297 ? io_dmem_s1_kill_1_REG_89 : _GEN_1298 ? io_dmem_s1_kill_1_REG_90 : _GEN_1293 ? io_dmem_s1_kill_1_REG_91 : _GEN_1288) : _GEN_1288;
  wire        dword_addr_matches_52_0 = stq_20_bits_addr_valid & ~stq_20_bits_addr_is_virtual & stq_20_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_52_1 = stq_20_bits_addr_valid & ~stq_20_bits_addr_is_virtual & stq_20_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_443;
  wire [14:0] _write_mask_mask_T_302 = 15'h1 << stq_20_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_306 = 15'h3 << {12'h0, stq_20_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_20_bits_uop_mem_size)
      2'b00:
        casez_tmp_443 = _write_mask_mask_T_302[7:0];
      2'b01:
        casez_tmp_443 = _write_mask_mask_T_306[7:0];
      2'b10:
        casez_tmp_443 = stq_20_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_443 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1300 = do_ld_search_0 & stq_20_valid & lcam_st_dep_mask_0[20];
  wire [7:0]  _GEN_1301 = casez_tmp_387 & casez_tmp_443;
  wire        _GEN_1302 = _GEN_1301 == casez_tmp_387 & ~stq_20_bits_uop_is_fence & ~stq_20_bits_uop_is_amo & dword_addr_matches_52_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_92;
  wire        _GEN_1303 = (|_GEN_1301) & dword_addr_matches_52_0;
  reg         io_dmem_s1_kill_0_REG_93;
  wire        _GEN_1304 = stq_20_bits_uop_is_fence | stq_20_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_94;
  wire        _GEN_1305 = _GEN_1300 ? (_GEN_1302 ? io_dmem_s1_kill_0_REG_92 : _GEN_1303 ? io_dmem_s1_kill_0_REG_93 : _GEN_1304 ? io_dmem_s1_kill_0_REG_94 : _GEN_1294) : _GEN_1294;
  wire        _GEN_1306 = do_ld_search_1 & stq_20_valid & lcam_st_dep_mask_1[20];
  wire [7:0]  _GEN_1307 = casez_tmp_388 & casez_tmp_443;
  wire        _GEN_1308 = _GEN_1307 == casez_tmp_388 & ~stq_20_bits_uop_is_fence & ~stq_20_bits_uop_is_amo & dword_addr_matches_52_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_92;
  wire        _GEN_1309 = (|_GEN_1307) & dword_addr_matches_52_1;
  reg         io_dmem_s1_kill_1_REG_93;
  reg         io_dmem_s1_kill_1_REG_94;
  wire        _GEN_1310 = _GEN_1306 ? (_GEN_1308 ? io_dmem_s1_kill_1_REG_92 : _GEN_1309 ? io_dmem_s1_kill_1_REG_93 : _GEN_1304 ? io_dmem_s1_kill_1_REG_94 : _GEN_1299) : _GEN_1299;
  wire        dword_addr_matches_53_0 = stq_21_bits_addr_valid & ~stq_21_bits_addr_is_virtual & stq_21_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_53_1 = stq_21_bits_addr_valid & ~stq_21_bits_addr_is_virtual & stq_21_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_444;
  wire [14:0] _write_mask_mask_T_317 = 15'h1 << stq_21_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_321 = 15'h3 << {12'h0, stq_21_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_21_bits_uop_mem_size)
      2'b00:
        casez_tmp_444 = _write_mask_mask_T_317[7:0];
      2'b01:
        casez_tmp_444 = _write_mask_mask_T_321[7:0];
      2'b10:
        casez_tmp_444 = stq_21_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_444 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1311 = do_ld_search_0 & stq_21_valid & lcam_st_dep_mask_0[21];
  wire [7:0]  _GEN_1312 = casez_tmp_387 & casez_tmp_444;
  wire        _GEN_1313 = _GEN_1312 == casez_tmp_387 & ~stq_21_bits_uop_is_fence & ~stq_21_bits_uop_is_amo & dword_addr_matches_53_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_95;
  wire        _GEN_1314 = (|_GEN_1312) & dword_addr_matches_53_0;
  reg         io_dmem_s1_kill_0_REG_96;
  wire        _GEN_1315 = stq_21_bits_uop_is_fence | stq_21_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_97;
  wire        _GEN_1316 = _GEN_1311 ? (_GEN_1313 ? io_dmem_s1_kill_0_REG_95 : _GEN_1314 ? io_dmem_s1_kill_0_REG_96 : _GEN_1315 ? io_dmem_s1_kill_0_REG_97 : _GEN_1305) : _GEN_1305;
  wire        _GEN_1317 = do_ld_search_1 & stq_21_valid & lcam_st_dep_mask_1[21];
  wire [7:0]  _GEN_1318 = casez_tmp_388 & casez_tmp_444;
  wire        _GEN_1319 = _GEN_1318 == casez_tmp_388 & ~stq_21_bits_uop_is_fence & ~stq_21_bits_uop_is_amo & dword_addr_matches_53_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_95;
  wire        _GEN_1320 = (|_GEN_1318) & dword_addr_matches_53_1;
  reg         io_dmem_s1_kill_1_REG_96;
  reg         io_dmem_s1_kill_1_REG_97;
  wire        _GEN_1321 = _GEN_1317 ? (_GEN_1319 ? io_dmem_s1_kill_1_REG_95 : _GEN_1320 ? io_dmem_s1_kill_1_REG_96 : _GEN_1315 ? io_dmem_s1_kill_1_REG_97 : _GEN_1310) : _GEN_1310;
  wire        dword_addr_matches_54_0 = stq_22_bits_addr_valid & ~stq_22_bits_addr_is_virtual & stq_22_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_54_1 = stq_22_bits_addr_valid & ~stq_22_bits_addr_is_virtual & stq_22_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_445;
  wire [14:0] _write_mask_mask_T_332 = 15'h1 << stq_22_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_336 = 15'h3 << {12'h0, stq_22_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_22_bits_uop_mem_size)
      2'b00:
        casez_tmp_445 = _write_mask_mask_T_332[7:0];
      2'b01:
        casez_tmp_445 = _write_mask_mask_T_336[7:0];
      2'b10:
        casez_tmp_445 = stq_22_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_445 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1322 = do_ld_search_0 & stq_22_valid & lcam_st_dep_mask_0[22];
  wire [7:0]  _GEN_1323 = casez_tmp_387 & casez_tmp_445;
  wire        _GEN_1324 = _GEN_1323 == casez_tmp_387 & ~stq_22_bits_uop_is_fence & ~stq_22_bits_uop_is_amo & dword_addr_matches_54_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_98;
  wire        _GEN_1325 = (|_GEN_1323) & dword_addr_matches_54_0;
  reg         io_dmem_s1_kill_0_REG_99;
  wire        _GEN_1326 = stq_22_bits_uop_is_fence | stq_22_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_100;
  wire        _GEN_1327 = _GEN_1322 ? (_GEN_1324 ? io_dmem_s1_kill_0_REG_98 : _GEN_1325 ? io_dmem_s1_kill_0_REG_99 : _GEN_1326 ? io_dmem_s1_kill_0_REG_100 : _GEN_1316) : _GEN_1316;
  wire        _GEN_1328 = do_ld_search_1 & stq_22_valid & lcam_st_dep_mask_1[22];
  wire [7:0]  _GEN_1329 = casez_tmp_388 & casez_tmp_445;
  wire        _GEN_1330 = _GEN_1329 == casez_tmp_388 & ~stq_22_bits_uop_is_fence & ~stq_22_bits_uop_is_amo & dword_addr_matches_54_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_98;
  wire        _GEN_1331 = (|_GEN_1329) & dword_addr_matches_54_1;
  reg         io_dmem_s1_kill_1_REG_99;
  reg         io_dmem_s1_kill_1_REG_100;
  wire        _GEN_1332 = _GEN_1328 ? (_GEN_1330 ? io_dmem_s1_kill_1_REG_98 : _GEN_1331 ? io_dmem_s1_kill_1_REG_99 : _GEN_1326 ? io_dmem_s1_kill_1_REG_100 : _GEN_1321) : _GEN_1321;
  wire        dword_addr_matches_55_0 = stq_23_bits_addr_valid & ~stq_23_bits_addr_is_virtual & stq_23_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_55_1 = stq_23_bits_addr_valid & ~stq_23_bits_addr_is_virtual & stq_23_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_446;
  wire [14:0] _write_mask_mask_T_347 = 15'h1 << stq_23_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_351 = 15'h3 << {12'h0, stq_23_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_23_bits_uop_mem_size)
      2'b00:
        casez_tmp_446 = _write_mask_mask_T_347[7:0];
      2'b01:
        casez_tmp_446 = _write_mask_mask_T_351[7:0];
      2'b10:
        casez_tmp_446 = stq_23_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_446 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1333 = do_ld_search_0 & stq_23_valid & lcam_st_dep_mask_0[23];
  wire [7:0]  _GEN_1334 = casez_tmp_387 & casez_tmp_446;
  wire        _GEN_1335 = _GEN_1334 == casez_tmp_387 & ~stq_23_bits_uop_is_fence & ~stq_23_bits_uop_is_amo & dword_addr_matches_55_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_101;
  wire        _GEN_1336 = (|_GEN_1334) & dword_addr_matches_55_0;
  reg         io_dmem_s1_kill_0_REG_102;
  wire        _GEN_1337 = stq_23_bits_uop_is_fence | stq_23_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_103;
  wire        _GEN_1338 = _GEN_1333 ? (_GEN_1335 ? io_dmem_s1_kill_0_REG_101 : _GEN_1336 ? io_dmem_s1_kill_0_REG_102 : _GEN_1337 ? io_dmem_s1_kill_0_REG_103 : _GEN_1327) : _GEN_1327;
  wire        _GEN_1339 = do_ld_search_1 & stq_23_valid & lcam_st_dep_mask_1[23];
  wire [7:0]  _GEN_1340 = casez_tmp_388 & casez_tmp_446;
  wire        _GEN_1341 = _GEN_1340 == casez_tmp_388 & ~stq_23_bits_uop_is_fence & ~stq_23_bits_uop_is_amo & dword_addr_matches_55_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_101;
  wire        _GEN_1342 = (|_GEN_1340) & dword_addr_matches_55_1;
  reg         io_dmem_s1_kill_1_REG_102;
  reg         io_dmem_s1_kill_1_REG_103;
  wire        _GEN_1343 = _GEN_1339 ? (_GEN_1341 ? io_dmem_s1_kill_1_REG_101 : _GEN_1342 ? io_dmem_s1_kill_1_REG_102 : _GEN_1337 ? io_dmem_s1_kill_1_REG_103 : _GEN_1332) : _GEN_1332;
  wire        dword_addr_matches_56_0 = stq_24_bits_addr_valid & ~stq_24_bits_addr_is_virtual & stq_24_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_56_1 = stq_24_bits_addr_valid & ~stq_24_bits_addr_is_virtual & stq_24_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_447;
  wire [14:0] _write_mask_mask_T_362 = 15'h1 << stq_24_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_366 = 15'h3 << {12'h0, stq_24_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_24_bits_uop_mem_size)
      2'b00:
        casez_tmp_447 = _write_mask_mask_T_362[7:0];
      2'b01:
        casez_tmp_447 = _write_mask_mask_T_366[7:0];
      2'b10:
        casez_tmp_447 = stq_24_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_447 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1344 = do_ld_search_0 & stq_24_valid & lcam_st_dep_mask_0[24];
  wire [7:0]  _GEN_1345 = casez_tmp_387 & casez_tmp_447;
  wire        _GEN_1346 = _GEN_1345 == casez_tmp_387 & ~stq_24_bits_uop_is_fence & ~stq_24_bits_uop_is_amo & dword_addr_matches_56_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_104;
  wire        _GEN_1347 = (|_GEN_1345) & dword_addr_matches_56_0;
  reg         io_dmem_s1_kill_0_REG_105;
  wire        _GEN_1348 = stq_24_bits_uop_is_fence | stq_24_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_106;
  wire        _GEN_1349 = _GEN_1344 ? (_GEN_1346 ? io_dmem_s1_kill_0_REG_104 : _GEN_1347 ? io_dmem_s1_kill_0_REG_105 : _GEN_1348 ? io_dmem_s1_kill_0_REG_106 : _GEN_1338) : _GEN_1338;
  wire        _GEN_1350 = do_ld_search_1 & stq_24_valid & lcam_st_dep_mask_1[24];
  wire [7:0]  _GEN_1351 = casez_tmp_388 & casez_tmp_447;
  wire        _GEN_1352 = _GEN_1351 == casez_tmp_388 & ~stq_24_bits_uop_is_fence & ~stq_24_bits_uop_is_amo & dword_addr_matches_56_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_104;
  wire        _GEN_1353 = (|_GEN_1351) & dword_addr_matches_56_1;
  reg         io_dmem_s1_kill_1_REG_105;
  reg         io_dmem_s1_kill_1_REG_106;
  wire        _GEN_1354 = _GEN_1350 ? (_GEN_1352 ? io_dmem_s1_kill_1_REG_104 : _GEN_1353 ? io_dmem_s1_kill_1_REG_105 : _GEN_1348 ? io_dmem_s1_kill_1_REG_106 : _GEN_1343) : _GEN_1343;
  wire        dword_addr_matches_57_0 = stq_25_bits_addr_valid & ~stq_25_bits_addr_is_virtual & stq_25_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_57_1 = stq_25_bits_addr_valid & ~stq_25_bits_addr_is_virtual & stq_25_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_448;
  wire [14:0] _write_mask_mask_T_377 = 15'h1 << stq_25_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_381 = 15'h3 << {12'h0, stq_25_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_25_bits_uop_mem_size)
      2'b00:
        casez_tmp_448 = _write_mask_mask_T_377[7:0];
      2'b01:
        casez_tmp_448 = _write_mask_mask_T_381[7:0];
      2'b10:
        casez_tmp_448 = stq_25_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_448 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1355 = do_ld_search_0 & stq_25_valid & lcam_st_dep_mask_0[25];
  wire [7:0]  _GEN_1356 = casez_tmp_387 & casez_tmp_448;
  wire        _GEN_1357 = _GEN_1356 == casez_tmp_387 & ~stq_25_bits_uop_is_fence & ~stq_25_bits_uop_is_amo & dword_addr_matches_57_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_107;
  wire        _GEN_1358 = (|_GEN_1356) & dword_addr_matches_57_0;
  reg         io_dmem_s1_kill_0_REG_108;
  wire        _GEN_1359 = stq_25_bits_uop_is_fence | stq_25_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_109;
  wire        _GEN_1360 = _GEN_1355 ? (_GEN_1357 ? io_dmem_s1_kill_0_REG_107 : _GEN_1358 ? io_dmem_s1_kill_0_REG_108 : _GEN_1359 ? io_dmem_s1_kill_0_REG_109 : _GEN_1349) : _GEN_1349;
  wire        _GEN_1361 = do_ld_search_1 & stq_25_valid & lcam_st_dep_mask_1[25];
  wire [7:0]  _GEN_1362 = casez_tmp_388 & casez_tmp_448;
  wire        _GEN_1363 = _GEN_1362 == casez_tmp_388 & ~stq_25_bits_uop_is_fence & ~stq_25_bits_uop_is_amo & dword_addr_matches_57_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_107;
  wire        _GEN_1364 = (|_GEN_1362) & dword_addr_matches_57_1;
  reg         io_dmem_s1_kill_1_REG_108;
  reg         io_dmem_s1_kill_1_REG_109;
  wire        _GEN_1365 = _GEN_1361 ? (_GEN_1363 ? io_dmem_s1_kill_1_REG_107 : _GEN_1364 ? io_dmem_s1_kill_1_REG_108 : _GEN_1359 ? io_dmem_s1_kill_1_REG_109 : _GEN_1354) : _GEN_1354;
  wire        dword_addr_matches_58_0 = stq_26_bits_addr_valid & ~stq_26_bits_addr_is_virtual & stq_26_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_58_1 = stq_26_bits_addr_valid & ~stq_26_bits_addr_is_virtual & stq_26_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_449;
  wire [14:0] _write_mask_mask_T_392 = 15'h1 << stq_26_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_396 = 15'h3 << {12'h0, stq_26_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_26_bits_uop_mem_size)
      2'b00:
        casez_tmp_449 = _write_mask_mask_T_392[7:0];
      2'b01:
        casez_tmp_449 = _write_mask_mask_T_396[7:0];
      2'b10:
        casez_tmp_449 = stq_26_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_449 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1366 = do_ld_search_0 & stq_26_valid & lcam_st_dep_mask_0[26];
  wire [7:0]  _GEN_1367 = casez_tmp_387 & casez_tmp_449;
  wire        _GEN_1368 = _GEN_1367 == casez_tmp_387 & ~stq_26_bits_uop_is_fence & ~stq_26_bits_uop_is_amo & dword_addr_matches_58_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_110;
  wire        _GEN_1369 = (|_GEN_1367) & dword_addr_matches_58_0;
  reg         io_dmem_s1_kill_0_REG_111;
  wire        _GEN_1370 = stq_26_bits_uop_is_fence | stq_26_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_112;
  wire        _GEN_1371 = _GEN_1366 ? (_GEN_1368 ? io_dmem_s1_kill_0_REG_110 : _GEN_1369 ? io_dmem_s1_kill_0_REG_111 : _GEN_1370 ? io_dmem_s1_kill_0_REG_112 : _GEN_1360) : _GEN_1360;
  wire        _GEN_1372 = do_ld_search_1 & stq_26_valid & lcam_st_dep_mask_1[26];
  wire [7:0]  _GEN_1373 = casez_tmp_388 & casez_tmp_449;
  wire        _GEN_1374 = _GEN_1373 == casez_tmp_388 & ~stq_26_bits_uop_is_fence & ~stq_26_bits_uop_is_amo & dword_addr_matches_58_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_110;
  wire        _GEN_1375 = (|_GEN_1373) & dword_addr_matches_58_1;
  reg         io_dmem_s1_kill_1_REG_111;
  reg         io_dmem_s1_kill_1_REG_112;
  wire        _GEN_1376 = _GEN_1372 ? (_GEN_1374 ? io_dmem_s1_kill_1_REG_110 : _GEN_1375 ? io_dmem_s1_kill_1_REG_111 : _GEN_1370 ? io_dmem_s1_kill_1_REG_112 : _GEN_1365) : _GEN_1365;
  wire        dword_addr_matches_59_0 = stq_27_bits_addr_valid & ~stq_27_bits_addr_is_virtual & stq_27_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_59_1 = stq_27_bits_addr_valid & ~stq_27_bits_addr_is_virtual & stq_27_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_450;
  wire [14:0] _write_mask_mask_T_407 = 15'h1 << stq_27_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_411 = 15'h3 << {12'h0, stq_27_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_27_bits_uop_mem_size)
      2'b00:
        casez_tmp_450 = _write_mask_mask_T_407[7:0];
      2'b01:
        casez_tmp_450 = _write_mask_mask_T_411[7:0];
      2'b10:
        casez_tmp_450 = stq_27_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_450 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1377 = do_ld_search_0 & stq_27_valid & lcam_st_dep_mask_0[27];
  wire [7:0]  _GEN_1378 = casez_tmp_387 & casez_tmp_450;
  wire        _GEN_1379 = _GEN_1378 == casez_tmp_387 & ~stq_27_bits_uop_is_fence & ~stq_27_bits_uop_is_amo & dword_addr_matches_59_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_113;
  wire        _GEN_1380 = (|_GEN_1378) & dword_addr_matches_59_0;
  reg         io_dmem_s1_kill_0_REG_114;
  wire        _GEN_1381 = stq_27_bits_uop_is_fence | stq_27_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_115;
  wire        _GEN_1382 = _GEN_1377 ? (_GEN_1379 ? io_dmem_s1_kill_0_REG_113 : _GEN_1380 ? io_dmem_s1_kill_0_REG_114 : _GEN_1381 ? io_dmem_s1_kill_0_REG_115 : _GEN_1371) : _GEN_1371;
  wire        _GEN_1383 = do_ld_search_1 & stq_27_valid & lcam_st_dep_mask_1[27];
  wire [7:0]  _GEN_1384 = casez_tmp_388 & casez_tmp_450;
  wire        _GEN_1385 = _GEN_1384 == casez_tmp_388 & ~stq_27_bits_uop_is_fence & ~stq_27_bits_uop_is_amo & dword_addr_matches_59_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_113;
  wire        _GEN_1386 = (|_GEN_1384) & dword_addr_matches_59_1;
  reg         io_dmem_s1_kill_1_REG_114;
  reg         io_dmem_s1_kill_1_REG_115;
  wire        _GEN_1387 = _GEN_1383 ? (_GEN_1385 ? io_dmem_s1_kill_1_REG_113 : _GEN_1386 ? io_dmem_s1_kill_1_REG_114 : _GEN_1381 ? io_dmem_s1_kill_1_REG_115 : _GEN_1376) : _GEN_1376;
  wire        dword_addr_matches_60_0 = stq_28_bits_addr_valid & ~stq_28_bits_addr_is_virtual & stq_28_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_60_1 = stq_28_bits_addr_valid & ~stq_28_bits_addr_is_virtual & stq_28_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_451;
  wire [14:0] _write_mask_mask_T_422 = 15'h1 << stq_28_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_426 = 15'h3 << {12'h0, stq_28_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_28_bits_uop_mem_size)
      2'b00:
        casez_tmp_451 = _write_mask_mask_T_422[7:0];
      2'b01:
        casez_tmp_451 = _write_mask_mask_T_426[7:0];
      2'b10:
        casez_tmp_451 = stq_28_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_451 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1388 = do_ld_search_0 & stq_28_valid & lcam_st_dep_mask_0[28];
  wire [7:0]  _GEN_1389 = casez_tmp_387 & casez_tmp_451;
  wire        _GEN_1390 = _GEN_1389 == casez_tmp_387 & ~stq_28_bits_uop_is_fence & ~stq_28_bits_uop_is_amo & dword_addr_matches_60_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_116;
  wire        _GEN_1391 = (|_GEN_1389) & dword_addr_matches_60_0;
  reg         io_dmem_s1_kill_0_REG_117;
  wire        _GEN_1392 = stq_28_bits_uop_is_fence | stq_28_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_118;
  wire        _GEN_1393 = _GEN_1388 ? (_GEN_1390 ? io_dmem_s1_kill_0_REG_116 : _GEN_1391 ? io_dmem_s1_kill_0_REG_117 : _GEN_1392 ? io_dmem_s1_kill_0_REG_118 : _GEN_1382) : _GEN_1382;
  wire        _GEN_1394 = do_ld_search_1 & stq_28_valid & lcam_st_dep_mask_1[28];
  wire [7:0]  _GEN_1395 = casez_tmp_388 & casez_tmp_451;
  wire        _GEN_1396 = _GEN_1395 == casez_tmp_388 & ~stq_28_bits_uop_is_fence & ~stq_28_bits_uop_is_amo & dword_addr_matches_60_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_116;
  wire        _GEN_1397 = (|_GEN_1395) & dword_addr_matches_60_1;
  reg         io_dmem_s1_kill_1_REG_117;
  reg         io_dmem_s1_kill_1_REG_118;
  wire        _GEN_1398 = _GEN_1394 ? (_GEN_1396 ? io_dmem_s1_kill_1_REG_116 : _GEN_1397 ? io_dmem_s1_kill_1_REG_117 : _GEN_1392 ? io_dmem_s1_kill_1_REG_118 : _GEN_1387) : _GEN_1387;
  wire        dword_addr_matches_61_0 = stq_29_bits_addr_valid & ~stq_29_bits_addr_is_virtual & stq_29_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_61_1 = stq_29_bits_addr_valid & ~stq_29_bits_addr_is_virtual & stq_29_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_452;
  wire [14:0] _write_mask_mask_T_437 = 15'h1 << stq_29_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_441 = 15'h3 << {12'h0, stq_29_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_29_bits_uop_mem_size)
      2'b00:
        casez_tmp_452 = _write_mask_mask_T_437[7:0];
      2'b01:
        casez_tmp_452 = _write_mask_mask_T_441[7:0];
      2'b10:
        casez_tmp_452 = stq_29_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_452 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1399 = do_ld_search_0 & stq_29_valid & lcam_st_dep_mask_0[29];
  wire [7:0]  _GEN_1400 = casez_tmp_387 & casez_tmp_452;
  wire        _GEN_1401 = _GEN_1400 == casez_tmp_387 & ~stq_29_bits_uop_is_fence & ~stq_29_bits_uop_is_amo & dword_addr_matches_61_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_119;
  wire        _GEN_1402 = (|_GEN_1400) & dword_addr_matches_61_0;
  reg         io_dmem_s1_kill_0_REG_120;
  wire        _GEN_1403 = stq_29_bits_uop_is_fence | stq_29_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_121;
  wire        _GEN_1404 = _GEN_1399 ? (_GEN_1401 ? io_dmem_s1_kill_0_REG_119 : _GEN_1402 ? io_dmem_s1_kill_0_REG_120 : _GEN_1403 ? io_dmem_s1_kill_0_REG_121 : _GEN_1393) : _GEN_1393;
  wire        _GEN_1405 = do_ld_search_1 & stq_29_valid & lcam_st_dep_mask_1[29];
  wire [7:0]  _GEN_1406 = casez_tmp_388 & casez_tmp_452;
  wire        _GEN_1407 = _GEN_1406 == casez_tmp_388 & ~stq_29_bits_uop_is_fence & ~stq_29_bits_uop_is_amo & dword_addr_matches_61_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_119;
  wire        _GEN_1408 = (|_GEN_1406) & dword_addr_matches_61_1;
  reg         io_dmem_s1_kill_1_REG_120;
  reg         io_dmem_s1_kill_1_REG_121;
  wire        _GEN_1409 = _GEN_1405 ? (_GEN_1407 ? io_dmem_s1_kill_1_REG_119 : _GEN_1408 ? io_dmem_s1_kill_1_REG_120 : _GEN_1403 ? io_dmem_s1_kill_1_REG_121 : _GEN_1398) : _GEN_1398;
  wire        dword_addr_matches_62_0 = stq_30_bits_addr_valid & ~stq_30_bits_addr_is_virtual & stq_30_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_62_1 = stq_30_bits_addr_valid & ~stq_30_bits_addr_is_virtual & stq_30_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_453;
  wire [14:0] _write_mask_mask_T_452 = 15'h1 << stq_30_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_456 = 15'h3 << {12'h0, stq_30_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_30_bits_uop_mem_size)
      2'b00:
        casez_tmp_453 = _write_mask_mask_T_452[7:0];
      2'b01:
        casez_tmp_453 = _write_mask_mask_T_456[7:0];
      2'b10:
        casez_tmp_453 = stq_30_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_453 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1410 = do_ld_search_0 & stq_30_valid & lcam_st_dep_mask_0[30];
  wire [7:0]  _GEN_1411 = casez_tmp_387 & casez_tmp_453;
  wire        _GEN_1412 = _GEN_1411 == casez_tmp_387 & ~stq_30_bits_uop_is_fence & ~stq_30_bits_uop_is_amo & dword_addr_matches_62_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_122;
  wire        _GEN_1413 = (|_GEN_1411) & dword_addr_matches_62_0;
  reg         io_dmem_s1_kill_0_REG_123;
  wire        _GEN_1414 = stq_30_bits_uop_is_fence | stq_30_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_124;
  wire        _GEN_1415 = _GEN_1410 ? (_GEN_1412 ? io_dmem_s1_kill_0_REG_122 : _GEN_1413 ? io_dmem_s1_kill_0_REG_123 : _GEN_1414 ? io_dmem_s1_kill_0_REG_124 : _GEN_1404) : _GEN_1404;
  wire        _GEN_1416 = do_ld_search_1 & stq_30_valid & lcam_st_dep_mask_1[30];
  wire [7:0]  _GEN_1417 = casez_tmp_388 & casez_tmp_453;
  wire        _GEN_1418 = _GEN_1417 == casez_tmp_388 & ~stq_30_bits_uop_is_fence & ~stq_30_bits_uop_is_amo & dword_addr_matches_62_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_122;
  wire        _GEN_1419 = (|_GEN_1417) & dword_addr_matches_62_1;
  reg         io_dmem_s1_kill_1_REG_123;
  reg         io_dmem_s1_kill_1_REG_124;
  wire        _GEN_1420 = _GEN_1416 ? (_GEN_1418 ? io_dmem_s1_kill_1_REG_122 : _GEN_1419 ? io_dmem_s1_kill_1_REG_123 : _GEN_1414 ? io_dmem_s1_kill_1_REG_124 : _GEN_1409) : _GEN_1409;
  wire        dword_addr_matches_63_0 = stq_31_bits_addr_valid & ~stq_31_bits_addr_is_virtual & stq_31_bits_addr_bits[32:3] == lcam_addr_0[32:3];
  wire        dword_addr_matches_63_1 = stq_31_bits_addr_valid & ~stq_31_bits_addr_is_virtual & stq_31_bits_addr_bits[32:3] == lcam_addr_1[32:3];
  reg  [7:0]  casez_tmp_454;
  wire [14:0] _write_mask_mask_T_467 = 15'h1 << stq_31_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_471 = 15'h3 << {12'h0, stq_31_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_31_bits_uop_mem_size)
      2'b00:
        casez_tmp_454 = _write_mask_mask_T_467[7:0];
      2'b01:
        casez_tmp_454 = _write_mask_mask_T_471[7:0];
      2'b10:
        casez_tmp_454 = stq_31_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_454 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1421 = do_ld_search_0 & stq_31_valid & lcam_st_dep_mask_0[31];
  wire [7:0]  _GEN_1422 = casez_tmp_387 & casez_tmp_454;
  wire        _GEN_1423 = _GEN_1422 == casez_tmp_387 & ~stq_31_bits_uop_is_fence & ~stq_31_bits_uop_is_amo & dword_addr_matches_63_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_125;
  wire        _GEN_1424 = (|_GEN_1422) & dword_addr_matches_63_0;
  reg         io_dmem_s1_kill_0_REG_126;
  wire        _GEN_1425 = stq_31_bits_uop_is_fence | stq_31_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_127;
  wire        _GEN_1426 = do_ld_search_1 & stq_31_valid & lcam_st_dep_mask_1[31];
  wire [7:0]  _GEN_1427 = casez_tmp_388 & casez_tmp_454;
  wire        _GEN_1428 = _GEN_1427 == casez_tmp_388 & ~stq_31_bits_uop_is_fence & ~stq_31_bits_uop_is_amo & dword_addr_matches_63_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_125;
  wire        _GEN_1429 = (|_GEN_1427) & dword_addr_matches_63_1;
  reg         io_dmem_s1_kill_1_REG_126;
  reg         io_dmem_s1_kill_1_REG_127;
  reg         casez_tmp_455;
  always @(*) begin
    casez (_forwarding_age_logic_0_io_forwarding_idx)
      5'b00000:
        casez_tmp_455 = _GEN_1080 & _GEN_1082;
      5'b00001:
        casez_tmp_455 = _GEN_1091 & _GEN_1093;
      5'b00010:
        casez_tmp_455 = _GEN_1102 & _GEN_1104;
      5'b00011:
        casez_tmp_455 = _GEN_1113 & _GEN_1115;
      5'b00100:
        casez_tmp_455 = _GEN_1124 & _GEN_1126;
      5'b00101:
        casez_tmp_455 = _GEN_1135 & _GEN_1137;
      5'b00110:
        casez_tmp_455 = _GEN_1146 & _GEN_1148;
      5'b00111:
        casez_tmp_455 = _GEN_1157 & _GEN_1159;
      5'b01000:
        casez_tmp_455 = _GEN_1168 & _GEN_1170;
      5'b01001:
        casez_tmp_455 = _GEN_1179 & _GEN_1181;
      5'b01010:
        casez_tmp_455 = _GEN_1190 & _GEN_1192;
      5'b01011:
        casez_tmp_455 = _GEN_1201 & _GEN_1203;
      5'b01100:
        casez_tmp_455 = _GEN_1212 & _GEN_1214;
      5'b01101:
        casez_tmp_455 = _GEN_1223 & _GEN_1225;
      5'b01110:
        casez_tmp_455 = _GEN_1234 & _GEN_1236;
      5'b01111:
        casez_tmp_455 = _GEN_1245 & _GEN_1247;
      5'b10000:
        casez_tmp_455 = _GEN_1256 & _GEN_1258;
      5'b10001:
        casez_tmp_455 = _GEN_1267 & _GEN_1269;
      5'b10010:
        casez_tmp_455 = _GEN_1278 & _GEN_1280;
      5'b10011:
        casez_tmp_455 = _GEN_1289 & _GEN_1291;
      5'b10100:
        casez_tmp_455 = _GEN_1300 & _GEN_1302;
      5'b10101:
        casez_tmp_455 = _GEN_1311 & _GEN_1313;
      5'b10110:
        casez_tmp_455 = _GEN_1322 & _GEN_1324;
      5'b10111:
        casez_tmp_455 = _GEN_1333 & _GEN_1335;
      5'b11000:
        casez_tmp_455 = _GEN_1344 & _GEN_1346;
      5'b11001:
        casez_tmp_455 = _GEN_1355 & _GEN_1357;
      5'b11010:
        casez_tmp_455 = _GEN_1366 & _GEN_1368;
      5'b11011:
        casez_tmp_455 = _GEN_1377 & _GEN_1379;
      5'b11100:
        casez_tmp_455 = _GEN_1388 & _GEN_1390;
      5'b11101:
        casez_tmp_455 = _GEN_1399 & _GEN_1401;
      5'b11110:
        casez_tmp_455 = _GEN_1410 & _GEN_1412;
      default:
        casez_tmp_455 = _GEN_1421 & _GEN_1423;
    endcase
  end // always @(*)
  reg         REG_2;
  reg         casez_tmp_456;
  always @(*) begin
    casez (_forwarding_age_logic_1_io_forwarding_idx)
      5'b00000:
        casez_tmp_456 = _GEN_1086 & _GEN_1088;
      5'b00001:
        casez_tmp_456 = _GEN_1097 & _GEN_1099;
      5'b00010:
        casez_tmp_456 = _GEN_1108 & _GEN_1110;
      5'b00011:
        casez_tmp_456 = _GEN_1119 & _GEN_1121;
      5'b00100:
        casez_tmp_456 = _GEN_1130 & _GEN_1132;
      5'b00101:
        casez_tmp_456 = _GEN_1141 & _GEN_1143;
      5'b00110:
        casez_tmp_456 = _GEN_1152 & _GEN_1154;
      5'b00111:
        casez_tmp_456 = _GEN_1163 & _GEN_1165;
      5'b01000:
        casez_tmp_456 = _GEN_1174 & _GEN_1176;
      5'b01001:
        casez_tmp_456 = _GEN_1185 & _GEN_1187;
      5'b01010:
        casez_tmp_456 = _GEN_1196 & _GEN_1198;
      5'b01011:
        casez_tmp_456 = _GEN_1207 & _GEN_1209;
      5'b01100:
        casez_tmp_456 = _GEN_1218 & _GEN_1220;
      5'b01101:
        casez_tmp_456 = _GEN_1229 & _GEN_1231;
      5'b01110:
        casez_tmp_456 = _GEN_1240 & _GEN_1242;
      5'b01111:
        casez_tmp_456 = _GEN_1251 & _GEN_1253;
      5'b10000:
        casez_tmp_456 = _GEN_1262 & _GEN_1264;
      5'b10001:
        casez_tmp_456 = _GEN_1273 & _GEN_1275;
      5'b10010:
        casez_tmp_456 = _GEN_1284 & _GEN_1286;
      5'b10011:
        casez_tmp_456 = _GEN_1295 & _GEN_1297;
      5'b10100:
        casez_tmp_456 = _GEN_1306 & _GEN_1308;
      5'b10101:
        casez_tmp_456 = _GEN_1317 & _GEN_1319;
      5'b10110:
        casez_tmp_456 = _GEN_1328 & _GEN_1330;
      5'b10111:
        casez_tmp_456 = _GEN_1339 & _GEN_1341;
      5'b11000:
        casez_tmp_456 = _GEN_1350 & _GEN_1352;
      5'b11001:
        casez_tmp_456 = _GEN_1361 & _GEN_1363;
      5'b11010:
        casez_tmp_456 = _GEN_1372 & _GEN_1374;
      5'b11011:
        casez_tmp_456 = _GEN_1383 & _GEN_1385;
      5'b11100:
        casez_tmp_456 = _GEN_1394 & _GEN_1396;
      5'b11101:
        casez_tmp_456 = _GEN_1405 & _GEN_1407;
      5'b11110:
        casez_tmp_456 = _GEN_1416 & _GEN_1418;
      default:
        casez_tmp_456 = _GEN_1426 & _GEN_1428;
    endcase
  end // always @(*)
  reg         REG_3;
  wire [5:0]  _l_idx_T_117 =
    _temp_bits_WIRE_1_41 & _temp_bits_T_18
      ? 6'h9
      : _temp_bits_WIRE_1_42 & _temp_bits_T_20 ? 6'hA : _temp_bits_WIRE_1_43 & _temp_bits_T_22 ? 6'hB : _temp_bits_WIRE_1_44 & _temp_bits_T_24 ? 6'hC : _temp_bits_WIRE_1_45 & _temp_bits_T_26 ? 6'hD : _temp_bits_WIRE_1_46 & _temp_bits_T_28 ? 6'hE : _temp_bits_WIRE_1_47 & ~(ldq_head[4]) ? 6'hF : _temp_bits_WIRE_1_48 & _temp_bits_T_32 ? 6'h10 : _temp_bits_WIRE_1_49 & _temp_bits_T_34 ? 6'h11 : _temp_bits_WIRE_1_50 & _temp_bits_T_36 ? 6'h12 : _temp_bits_WIRE_1_51 & _temp_bits_T_38 ? 6'h13 : _temp_bits_WIRE_1_52 & _temp_bits_T_40 ? 6'h14 : _temp_bits_WIRE_1_53 & _temp_bits_T_42 ? 6'h15 : _temp_bits_WIRE_1_54 & _temp_bits_T_44 ? 6'h16 : _temp_bits_WIRE_1_55 & _temp_bits_T_46 ? 6'h17 : _temp_bits_WIRE_1_56 & _temp_bits_T_48 ? 6'h18 : _temp_bits_WIRE_1_57 & _temp_bits_T_50 ? 6'h19 : _temp_bits_WIRE_1_58 & _temp_bits_T_52 ? 6'h1A : _temp_bits_WIRE_1_59 & _temp_bits_T_54 ? 6'h1B : _temp_bits_WIRE_1_60 & _temp_bits_T_56 ? 6'h1C : _temp_bits_WIRE_1_61 & _temp_bits_T_58 ? 6'h1D : _temp_bits_WIRE_1_62 & _temp_bits_T_60 ? 6'h1E : _temp_bits_WIRE_1_63 ? 6'h1F : _temp_bits_WIRE_1_32 ? 6'h20 : _temp_bits_WIRE_1_33 ? 6'h21 : _temp_bits_WIRE_1_34 ? 6'h22 : _temp_bits_WIRE_1_35 ? 6'h23 : _temp_bits_WIRE_1_36 ? 6'h24 : _temp_bits_WIRE_1_37 ? 6'h25 : _temp_bits_WIRE_1_38 ? 6'h26 : _temp_bits_WIRE_1_39 ? 6'h27 : _temp_bits_WIRE_1_40 ? 6'h28 : _temp_bits_WIRE_1_41 ? 6'h29 : _temp_bits_WIRE_1_42 ? 6'h2A : _temp_bits_WIRE_1_43 ? 6'h2B : _temp_bits_WIRE_1_44 ? 6'h2C : _temp_bits_WIRE_1_45 ? 6'h2D : _temp_bits_WIRE_1_46 ? 6'h2E : _temp_bits_WIRE_1_47 ? 6'h2F : _temp_bits_WIRE_1_48 ? 6'h30 : _temp_bits_WIRE_1_49 ? 6'h31 : _temp_bits_WIRE_1_50 ? 6'h32 : _temp_bits_WIRE_1_51 ? 6'h33 : _temp_bits_WIRE_1_52 ? 6'h34 : _temp_bits_WIRE_1_53 ? 6'h35 : _temp_bits_WIRE_1_54 ? 6'h36 : _temp_bits_WIRE_1_55 ? 6'h37 : _temp_bits_WIRE_1_56 ? 6'h38 : _temp_bits_WIRE_1_57 ? 6'h39 : _temp_bits_WIRE_1_58 ? 6'h3A : _temp_bits_WIRE_1_59 ? 6'h3B : _temp_bits_WIRE_1_60 ? 6'h3C : _temp_bits_WIRE_1_61 ? 6'h3D : {5'h1F, ~_temp_bits_WIRE_1_62};
  wire [4:0]  l_idx = _temp_bits_WIRE_1_32 & _temp_bits_T ? 5'h0 : _temp_bits_WIRE_1_33 & _temp_bits_T_2 ? 5'h1 : _temp_bits_WIRE_1_34 & _temp_bits_T_4 ? 5'h2 : _temp_bits_WIRE_1_35 & _temp_bits_T_6 ? 5'h3 : _temp_bits_WIRE_1_36 & _temp_bits_T_8 ? 5'h4 : _temp_bits_WIRE_1_37 & _temp_bits_T_10 ? 5'h5 : _temp_bits_WIRE_1_38 & _temp_bits_T_12 ? 5'h6 : _temp_bits_WIRE_1_39 & _temp_bits_T_14 ? 5'h7 : _temp_bits_WIRE_1_40 & _temp_bits_T_16 ? 5'h8 : _l_idx_T_117[4:0];
  reg         r_xcpt_valid;
  reg  [19:0] r_xcpt_uop_br_mask;
  reg  [6:0]  r_xcpt_uop_rob_idx;
  reg  [4:0]  r_xcpt_cause;
  reg  [39:0] r_xcpt_badvaddr;
  reg  [19:0] casez_tmp_457;
  always @(*) begin
    casez (l_idx)
      5'b00000:
        casez_tmp_457 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_457 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_457 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_457 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_457 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_457 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_457 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_457 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_457 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_457 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_457 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_457 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_457 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_457 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_457 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_457 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_457 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_457 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_457 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_457 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_457 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_457 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_457 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_457 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_457 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_457 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_457 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_457 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_457 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_457 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_457 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_457 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_458;
  always @(*) begin
    casez (l_idx)
      5'b00000:
        casez_tmp_458 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_458 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_458 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_458 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_458 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_458 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_458 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_458 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_458 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_458 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_458 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_458 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_458 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_458 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_458 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_458 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_458 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_458 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_458 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_458 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_458 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_458 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_458 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_458 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_458 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_458 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_458 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_458 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_458 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_458 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_458 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_458 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  wire        _io_core_spec_ld_wakeup_0_valid_output = fired_load_incoming_REG & ~mem_incoming_uop_0_fp_val & (|mem_incoming_uop_0_pdst);
  wire        _io_core_spec_ld_wakeup_1_valid_output = fired_load_incoming_REG_1 & ~mem_incoming_uop_1_fp_val & (|mem_incoming_uop_1_pdst);
  wire        _GEN_1430 = io_dmem_nack_0_valid & io_dmem_nack_0_bits_is_hella;
  wire        _GEN_1431 = hella_state == 3'h4;
  wire        _GEN_1432 = hella_state == 3'h6;
  wire        _GEN_1433 = io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella;
  wire        _GEN_1434 = _GEN_1433 & io_dmem_nack_0_bits_uop_uses_ldq & ~reset;
  reg         casez_tmp_459;
  always @(*) begin
    casez (io_dmem_nack_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_459 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_459 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_459 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_459 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_459 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_459 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_459 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_459 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_459 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_459 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_459 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_459 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_459 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_459 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_459 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_459 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_459 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_459 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_459 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_459 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_459 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_459 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_459 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_459 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_459 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_459 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_459 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_459 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_459 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_459 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_459 = ldq_30_bits_executed;
      default:
        casez_tmp_459 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  wire        _GEN_1435 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h0;
  wire        _GEN_1436 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1;
  wire        _GEN_1437 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h2;
  wire        _GEN_1438 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h3;
  wire        _GEN_1439 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h4;
  wire        _GEN_1440 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h5;
  wire        _GEN_1441 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h6;
  wire        _GEN_1442 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h7;
  wire        _GEN_1443 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h8;
  wire        _GEN_1444 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h9;
  wire        _GEN_1445 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hA;
  wire        _GEN_1446 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hB;
  wire        _GEN_1447 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hC;
  wire        _GEN_1448 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hD;
  wire        _GEN_1449 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hE;
  wire        _GEN_1450 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hF;
  wire        _GEN_1451 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h10;
  wire        _GEN_1452 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h11;
  wire        _GEN_1453 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h12;
  wire        _GEN_1454 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h13;
  wire        _GEN_1455 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h14;
  wire        _GEN_1456 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h15;
  wire        _GEN_1457 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h16;
  wire        _GEN_1458 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h17;
  wire        _GEN_1459 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h18;
  wire        _GEN_1460 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h19;
  wire        _GEN_1461 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1A;
  wire        _GEN_1462 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1B;
  wire        _GEN_1463 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1C;
  wire        _GEN_1464 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1D;
  wire        _GEN_1465 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1E;
  wire        _GEN_1466 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq;
  reg  [6:0]  casez_tmp_460;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_460 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_460 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_460 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_460 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_460 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_460 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_460 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_460 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_460 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_460 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_460 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_460 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_460 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_460 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_460 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_460 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_460 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_460 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_460 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_460 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_460 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_460 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_460 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_460 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_460 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_460 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_460 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_460 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_460 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_460 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_460 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_460 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_461;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_461 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_461 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_461 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_461 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_461 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_461 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_461 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_461 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_461 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_461 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_461 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_461 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_461 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_461 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_461 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_461 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_461 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_461 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_461 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_461 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_461 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_461 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_461 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_461 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_461 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_461 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_461 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_461 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_461 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_461 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_461 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_461 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_462;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_462 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_462 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_462 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_462 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_462 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_462 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_462 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_462 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_462 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_462 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_462 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_462 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_462 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_462 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_462 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_462 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_462 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_462 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_462 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_462 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_462 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_462 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_462 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_462 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_462 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_462 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_462 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_462 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_462 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_462 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_462 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_462 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_463;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_463 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_463 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_463 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_463 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_463 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_463 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_463 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_463 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_463 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_463 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_463 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_463 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_463 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_463 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_463 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_463 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_463 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_463 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_463 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_463 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_463 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_463 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_463 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_463 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_463 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_463 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_463 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_463 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_463 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_463 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_463 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_463 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_464;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_464 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_464 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_464 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_464 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_464 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_464 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_464 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_464 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_464 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_464 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_464 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_464 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_464 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_464 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_464 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_464 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_464 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_464 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_464 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_464 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_464 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_464 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_464 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_464 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_464 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_464 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_464 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_464 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_464 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_464 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_464 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_464 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_465;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_465 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_465 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_465 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_465 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_465 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_465 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_465 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_465 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_465 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_465 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_465 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_465 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_465 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_465 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_465 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_465 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_465 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_465 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_465 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_465 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_465 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_465 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_465 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_465 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_465 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_465 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_465 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_465 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_465 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_465 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_465 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_465 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_466;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_466 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_466 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_466 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_466 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_466 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_466 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_466 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_466 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_466 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_466 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_466 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_466 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_466 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_466 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_466 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_466 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_466 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_466 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_466 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_466 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_466 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_466 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_466 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_466 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_466 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_466 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_466 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_466 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_466 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_466 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_466 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_466 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_467;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_467 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_467 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_467 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_467 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_467 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_467 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_467 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_467 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_467 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_467 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_467 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_467 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_467 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_467 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_467 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_467 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_467 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_467 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_467 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_467 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_467 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_467 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_467 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_467 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_467 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_467 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_467 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_467 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_467 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_467 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_467 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_467 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_468;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_468 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_468 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_468 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_468 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_468 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_468 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_468 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_468 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_468 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_468 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_468 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_468 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_468 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_468 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_468 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_468 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_468 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_468 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_468 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_468 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_468 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_468 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_468 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_468 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_468 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_468 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_468 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_468 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_468 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_468 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_468 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_468 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_469;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_469 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_469 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_469 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_469 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_469 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_469 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_469 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_469 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_469 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_469 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_469 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_469 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_469 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_469 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_469 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_469 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_469 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_469 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_469 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_469 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_469 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_469 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_469 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_469 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_469 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_469 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_469 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_469 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_469 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_469 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_469 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_469 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_470;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_470 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_470 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_470 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_470 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_470 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_470 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_470 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_470 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_470 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_470 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_470 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_470 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_470 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_470 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_470 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_470 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_470 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_470 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_470 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_470 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_470 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_470 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_470 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_470 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_470 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_470 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_470 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_470 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_470 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_470 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_470 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_470 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  wire        send_iresp = casez_tmp_469 == 2'h0;
  wire        send_fresp = casez_tmp_469 == 2'h1;
  reg  [6:0]  casez_tmp_471;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_471 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_471 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_471 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_471 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_471 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_471 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_471 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_471 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_471 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_471 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_471 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_471 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_471 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_471 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_471 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_471 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_471 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_471 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_471 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_471 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_471 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_471 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_471 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_471 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_471 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_471 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_471 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_471 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_471 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_471 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_471 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_471 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_472;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_472 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_472 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_472 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_472 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_472 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_472 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_472 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_472 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_472 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_472 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_472 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_472 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_472 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_472 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_472 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_472 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_472 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_472 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_472 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_472 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_472 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_472 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_472 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_472 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_472 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_472 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_472 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_472 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_472 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_472 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_472 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_472 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_473;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_473 = stq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_473 = stq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_473 = stq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_473 = stq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_473 = stq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_473 = stq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_473 = stq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_473 = stq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_473 = stq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_473 = stq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_473 = stq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_473 = stq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_473 = stq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_473 = stq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_473 = stq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_473 = stq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_473 = stq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_473 = stq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_473 = stq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_473 = stq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_473 = stq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_473 = stq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_473 = stq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_473 = stq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_473 = stq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_473 = stq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_473 = stq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_473 = stq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_473 = stq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_473 = stq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_473 = stq_30_bits_uop_pdst;
      default:
        casez_tmp_473 = stq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_474;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_474 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_474 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_474 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_474 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_474 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_474 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_474 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_474 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_474 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_474 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_474 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_474 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_474 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_474 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_474 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_474 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_474 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_474 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_474 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_474 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_474 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_474 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_474 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_474 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_474 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_474 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_474 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_474 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_474 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_474 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_474 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_474 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_475;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_475 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_475 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_475 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_475 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_475 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_475 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_475 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_475 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_475 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_475 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_475 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_475 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_475 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_475 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_475 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_475 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_475 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_475 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_475 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_475 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_475 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_475 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_475 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_475 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_475 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_475 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_475 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_475 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_475 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_475 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_475 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_475 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_476;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_476 = stq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_476 = stq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_476 = stq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_476 = stq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_476 = stq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_476 = stq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_476 = stq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_476 = stq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_476 = stq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_476 = stq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_476 = stq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_476 = stq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_476 = stq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_476 = stq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_476 = stq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_476 = stq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_476 = stq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_476 = stq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_476 = stq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_476 = stq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_476 = stq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_476 = stq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_476 = stq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_476 = stq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_476 = stq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_476 = stq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_476 = stq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_476 = stq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_476 = stq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_476 = stq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_476 = stq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_476 = stq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  wire        _GEN_1467 = io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_is_amo;
  wire        dmem_resp_fired_0 = io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq | _GEN_1467);
  wire        _GEN_1468 = dmem_resp_fired_0 & wb_forward_valid_0;
  wire        _GEN_1469 = ~dmem_resp_fired_0 & wb_forward_valid_0;
  reg  [6:0]  casez_tmp_477;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_477 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_477 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_477 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_477 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_477 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_477 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_477 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_477 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_477 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_477 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_477 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_477 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_477 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_477 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_477 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_477 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_477 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_477 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_477 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_477 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_477 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_477 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_477 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_477 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_477 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_477 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_477 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_477 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_477 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_477 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_477 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_477 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_478;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_478 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_478 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_478 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_478 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_478 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_478 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_478 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_478 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_478 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_478 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_478 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_478 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_478 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_478 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_478 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_478 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_478 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_478 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_478 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_478 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_478 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_478 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_478 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_478 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_478 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_478 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_478 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_478 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_478 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_478 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_478 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_478 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_479;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_479 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_479 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_479 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_479 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_479 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_479 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_479 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_479 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_479 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_479 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_479 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_479 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_479 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_479 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_479 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_479 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_479 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_479 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_479 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_479 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_479 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_479 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_479 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_479 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_479 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_479 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_479 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_479 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_479 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_479 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_479 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_479 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_480;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_480 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_480 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_480 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_480 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_480 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_480 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_480 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_480 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_480 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_480 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_480 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_480 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_480 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_480 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_480 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_480 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_480 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_480 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_480 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_480 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_480 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_480 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_480 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_480 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_480 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_480 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_480 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_480 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_480 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_480 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_480 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_480 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_481;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_481 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_481 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_481 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_481 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_481 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_481 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_481 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_481 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_481 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_481 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_481 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_481 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_481 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_481 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_481 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_481 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_481 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_481 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_481 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_481 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_481 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_481 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_481 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_481 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_481 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_481 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_481 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_481 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_481 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_481 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_481 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_481 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_482;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_482 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_482 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_482 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_482 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_482 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_482 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_482 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_482 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_482 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_482 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_482 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_482 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_482 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_482 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_482 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_482 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_482 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_482 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_482 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_482 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_482 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_482 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_482 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_482 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_482 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_482 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_482 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_482 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_482 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_482 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_482 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_482 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_483;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_483 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_483 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_483 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_483 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_483 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_483 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_483 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_483 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_483 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_483 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_483 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_483 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_483 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_483 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_483 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_483 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_483 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_483 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_483 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_483 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_483 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_483 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_483 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_483 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_483 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_483 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_483 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_483 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_483 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_483 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_483 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_483 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_484;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_484 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_484 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_484 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_484 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_484 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_484 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_484 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_484 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_484 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_484 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_484 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_484 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_484 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_484 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_484 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_484 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_484 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_484 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_484 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_484 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_484 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_484 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_484 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_484 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_484 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_484 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_484 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_484 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_484 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_484 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_484 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_484 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  reg         casez_tmp_485;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_485 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_485 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_485 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_485 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_485 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_485 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_485 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_485 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_485 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_485 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_485 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_485 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_485 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_485 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_485 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_485 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_485 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_485 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_485 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_485 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_485 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_485 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_485 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_485 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_485 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_485 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_485 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_485 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_485 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_485 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_485 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_485 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_486;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_486 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_486 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_486 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_486 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_486 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_486 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_486 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_486 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_486 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_486 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_486 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_486 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_486 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_486 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_486 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_486 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_486 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_486 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_486 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_486 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_486 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_486 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_486 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_486 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_486 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_486 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_486 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_486 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_486 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_486 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_486 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_486 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_487;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_487 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_487 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_487 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_487 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_487 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_487 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_487 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_487 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_487 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_487 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_487 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_487 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_487 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_487 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_487 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_487 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_487 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_487 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_487 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_487 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_487 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_487 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_487 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_487 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_487 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_487 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_487 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_487 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_487 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_487 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_487 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_487 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_488;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_488 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_488 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_488 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_488 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_488 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_488 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_488 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_488 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_488 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_488 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_488 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_488 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_488 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_488 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_488 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_488 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_488 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_488 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_488 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_488 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_488 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_488 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_488 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_488 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_488 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_488 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_488 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_488 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_488 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_488 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_488 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_488 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  wire        live = (io_core_brupdate_b1_mispredict_mask & casez_tmp_478) == 20'h0;
  reg  [1:0]  casez_tmp_489;
  always @(*) begin
    casez (wb_forward_stq_idx_0)
      5'b00000:
        casez_tmp_489 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_489 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_489 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_489 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_489 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_489 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_489 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_489 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_489 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_489 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_489 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_489 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_489 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_489 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_489 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_489 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_489 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_489 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_489 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_489 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_489 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_489 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_489 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_489 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_489 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_489 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_489 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_489 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_489 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_489 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_489 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_489 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_490;
  always @(*) begin
    casez (wb_forward_stq_idx_0)
      5'b00000:
        casez_tmp_490 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_490 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_490 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_490 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_490 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_490 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_490 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_490 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_490 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_490 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_490 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_490 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_490 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_490 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_490 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_490 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_490 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_490 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_490 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_490 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_490 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_490 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_490 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_490 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_490 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_490 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_490 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_490 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_490 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_490 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_490 = stq_30_bits_data_valid;
      default:
        casez_tmp_490 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_491;
  always @(*) begin
    casez (wb_forward_stq_idx_0)
      5'b00000:
        casez_tmp_491 = stq_0_bits_data_bits;
      5'b00001:
        casez_tmp_491 = stq_1_bits_data_bits;
      5'b00010:
        casez_tmp_491 = stq_2_bits_data_bits;
      5'b00011:
        casez_tmp_491 = stq_3_bits_data_bits;
      5'b00100:
        casez_tmp_491 = stq_4_bits_data_bits;
      5'b00101:
        casez_tmp_491 = stq_5_bits_data_bits;
      5'b00110:
        casez_tmp_491 = stq_6_bits_data_bits;
      5'b00111:
        casez_tmp_491 = stq_7_bits_data_bits;
      5'b01000:
        casez_tmp_491 = stq_8_bits_data_bits;
      5'b01001:
        casez_tmp_491 = stq_9_bits_data_bits;
      5'b01010:
        casez_tmp_491 = stq_10_bits_data_bits;
      5'b01011:
        casez_tmp_491 = stq_11_bits_data_bits;
      5'b01100:
        casez_tmp_491 = stq_12_bits_data_bits;
      5'b01101:
        casez_tmp_491 = stq_13_bits_data_bits;
      5'b01110:
        casez_tmp_491 = stq_14_bits_data_bits;
      5'b01111:
        casez_tmp_491 = stq_15_bits_data_bits;
      5'b10000:
        casez_tmp_491 = stq_16_bits_data_bits;
      5'b10001:
        casez_tmp_491 = stq_17_bits_data_bits;
      5'b10010:
        casez_tmp_491 = stq_18_bits_data_bits;
      5'b10011:
        casez_tmp_491 = stq_19_bits_data_bits;
      5'b10100:
        casez_tmp_491 = stq_20_bits_data_bits;
      5'b10101:
        casez_tmp_491 = stq_21_bits_data_bits;
      5'b10110:
        casez_tmp_491 = stq_22_bits_data_bits;
      5'b10111:
        casez_tmp_491 = stq_23_bits_data_bits;
      5'b11000:
        casez_tmp_491 = stq_24_bits_data_bits;
      5'b11001:
        casez_tmp_491 = stq_25_bits_data_bits;
      5'b11010:
        casez_tmp_491 = stq_26_bits_data_bits;
      5'b11011:
        casez_tmp_491 = stq_27_bits_data_bits;
      5'b11100:
        casez_tmp_491 = stq_28_bits_data_bits;
      5'b11101:
        casez_tmp_491 = stq_29_bits_data_bits;
      5'b11110:
        casez_tmp_491 = stq_30_bits_data_bits;
      default:
        casez_tmp_491 = stq_31_bits_data_bits;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_492;
  always @(*) begin
    casez (casez_tmp_489)
      2'b00:
        casez_tmp_492 = {2{{2{{2{casez_tmp_491[7:0]}}}}}};
      2'b01:
        casez_tmp_492 = {2{{2{casez_tmp_491[15:0]}}}};
      2'b10:
        casez_tmp_492 = {2{casez_tmp_491[31:0]}};
      default:
        casez_tmp_492 = casez_tmp_491;
    endcase
  end // always @(*)
  wire        _GEN_1470 = _GEN_1468 | ~_GEN_1469;
  wire        _io_core_exe_0_iresp_valid_output = _GEN_1470 ? io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq ? send_iresp : _GEN_1467) : casez_tmp_487 == 2'h0 & casez_tmp_490 & live;
  wire        _io_core_exe_0_fresp_valid_output = _GEN_1470 ? _GEN_1466 & send_fresp : casez_tmp_487 == 2'h1 & casez_tmp_490 & live;
  wire [31:0] io_core_exe_0_iresp_bits_data_zeroed = wb_forward_ld_addr_0[2] ? casez_tmp_492[63:32] : casez_tmp_492[31:0];
  wire        _ldq_bits_debug_wb_data_T_1 = casez_tmp_483 == 2'h2;
  wire [15:0] io_core_exe_0_iresp_bits_data_zeroed_1 = wb_forward_ld_addr_0[1] ? io_core_exe_0_iresp_bits_data_zeroed[31:16] : io_core_exe_0_iresp_bits_data_zeroed[15:0];
  wire        _ldq_bits_debug_wb_data_T_10 = casez_tmp_483 == 2'h1;
  wire [7:0]  io_core_exe_0_iresp_bits_data_zeroed_2 = wb_forward_ld_addr_0[0] ? io_core_exe_0_iresp_bits_data_zeroed_1[15:8] : io_core_exe_0_iresp_bits_data_zeroed_1[7:0];
  wire        _ldq_bits_debug_wb_data_T_19 = casez_tmp_483 == 2'h0;
  wire [31:0] io_core_exe_0_fresp_bits_data_zeroed = wb_forward_ld_addr_0[2] ? casez_tmp_492[63:32] : casez_tmp_492[31:0];
  wire [15:0] io_core_exe_0_fresp_bits_data_zeroed_1 = wb_forward_ld_addr_0[1] ? io_core_exe_0_fresp_bits_data_zeroed[31:16] : io_core_exe_0_fresp_bits_data_zeroed[15:0];
  wire [7:0]  io_core_exe_0_fresp_bits_data_zeroed_2 = wb_forward_ld_addr_0[0] ? io_core_exe_0_fresp_bits_data_zeroed_1[15:8] : io_core_exe_0_fresp_bits_data_zeroed_1[7:0];
  wire        _GEN_1471 = io_dmem_nack_1_valid & io_dmem_nack_1_bits_is_hella;
  wire        _GEN_1472 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella;
  wire        _GEN_1473 = _GEN_1472 & io_dmem_nack_1_bits_uop_uses_ldq & ~reset;
  reg         casez_tmp_493;
  always @(*) begin
    casez (io_dmem_nack_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_493 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_493 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_493 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_493 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_493 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_493 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_493 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_493 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_493 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_493 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_493 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_493 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_493 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_493 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_493 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_493 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_493 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_493 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_493 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_493 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_493 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_493 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_493 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_493 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_493 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_493 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_493 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_493 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_493 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_493 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_493 = ldq_30_bits_executed;
      default:
        casez_tmp_493 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  wire        _GEN_1474 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h0;
  wire        _GEN_1475 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1;
  wire        _GEN_1476 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h2;
  wire        _GEN_1477 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h3;
  wire        _GEN_1478 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h4;
  wire        _GEN_1479 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h5;
  wire        _GEN_1480 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h6;
  wire        _GEN_1481 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h7;
  wire        _GEN_1482 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h8;
  wire        _GEN_1483 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h9;
  wire        _GEN_1484 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hA;
  wire        _GEN_1485 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hB;
  wire        _GEN_1486 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hC;
  wire        _GEN_1487 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hD;
  wire        _GEN_1488 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hE;
  wire        _GEN_1489 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hF;
  wire        _GEN_1490 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h10;
  wire        _GEN_1491 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h11;
  wire        _GEN_1492 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h12;
  wire        _GEN_1493 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h13;
  wire        _GEN_1494 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h14;
  wire        _GEN_1495 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h15;
  wire        _GEN_1496 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h16;
  wire        _GEN_1497 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h17;
  wire        _GEN_1498 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h18;
  wire        _GEN_1499 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h19;
  wire        _GEN_1500 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1A;
  wire        _GEN_1501 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1B;
  wire        _GEN_1502 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1C;
  wire        _GEN_1503 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1D;
  wire        _GEN_1504 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1E;
  wire        _GEN_1505 = io_dmem_nack_1_bits_uop_uses_ldq & (&io_dmem_nack_1_bits_uop_ldq_idx);
  assign nacking_loads_0 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1474 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1435;
  assign nacking_loads_1 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1475 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1436;
  assign nacking_loads_2 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1476 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1437;
  assign nacking_loads_3 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1477 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1438;
  assign nacking_loads_4 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1478 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1439;
  assign nacking_loads_5 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1479 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1440;
  assign nacking_loads_6 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1480 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1441;
  assign nacking_loads_7 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1481 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1442;
  assign nacking_loads_8 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1482 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1443;
  assign nacking_loads_9 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1483 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1444;
  assign nacking_loads_10 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1484 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1445;
  assign nacking_loads_11 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1485 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1446;
  assign nacking_loads_12 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1486 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1447;
  assign nacking_loads_13 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1487 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1448;
  assign nacking_loads_14 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1488 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1449;
  assign nacking_loads_15 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1489 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1450;
  assign nacking_loads_16 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1490 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1451;
  assign nacking_loads_17 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1491 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1452;
  assign nacking_loads_18 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1492 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1453;
  assign nacking_loads_19 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1493 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1454;
  assign nacking_loads_20 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1494 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1455;
  assign nacking_loads_21 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1495 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1456;
  assign nacking_loads_22 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1496 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1457;
  assign nacking_loads_23 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1497 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1458;
  assign nacking_loads_24 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1498 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1459;
  assign nacking_loads_25 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1499 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1460;
  assign nacking_loads_26 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1500 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1461;
  assign nacking_loads_27 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1501 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1462;
  assign nacking_loads_28 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1502 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1463;
  assign nacking_loads_29 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1503 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1464;
  assign nacking_loads_30 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1504 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1465;
  assign nacking_loads_31 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_1505 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & (&io_dmem_nack_0_bits_uop_ldq_idx);
  wire        _GEN_1506 = io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq;
  reg  [6:0]  casez_tmp_494;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_494 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_494 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_494 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_494 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_494 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_494 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_494 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_494 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_494 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_494 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_494 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_494 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_494 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_494 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_494 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_494 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_494 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_494 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_494 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_494 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_494 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_494 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_494 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_494 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_494 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_494 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_494 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_494 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_494 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_494 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_494 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_494 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_495;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_495 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_495 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_495 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_495 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_495 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_495 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_495 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_495 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_495 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_495 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_495 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_495 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_495 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_495 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_495 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_495 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_495 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_495 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_495 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_495 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_495 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_495 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_495 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_495 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_495 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_495 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_495 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_495 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_495 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_495 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_495 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_495 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_496;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_496 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_496 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_496 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_496 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_496 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_496 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_496 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_496 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_496 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_496 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_496 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_496 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_496 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_496 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_496 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_496 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_496 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_496 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_496 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_496 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_496 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_496 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_496 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_496 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_496 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_496 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_496 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_496 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_496 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_496 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_496 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_496 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_497;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_497 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_497 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_497 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_497 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_497 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_497 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_497 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_497 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_497 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_497 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_497 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_497 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_497 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_497 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_497 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_497 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_497 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_497 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_497 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_497 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_497 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_497 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_497 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_497 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_497 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_497 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_497 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_497 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_497 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_497 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_497 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_497 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_498;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_498 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_498 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_498 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_498 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_498 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_498 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_498 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_498 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_498 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_498 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_498 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_498 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_498 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_498 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_498 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_498 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_498 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_498 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_498 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_498 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_498 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_498 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_498 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_498 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_498 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_498 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_498 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_498 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_498 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_498 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_498 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_498 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_499;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_499 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_499 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_499 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_499 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_499 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_499 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_499 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_499 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_499 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_499 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_499 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_499 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_499 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_499 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_499 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_499 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_499 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_499 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_499 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_499 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_499 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_499 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_499 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_499 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_499 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_499 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_499 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_499 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_499 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_499 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_499 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_499 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_500;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_500 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_500 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_500 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_500 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_500 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_500 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_500 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_500 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_500 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_500 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_500 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_500 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_500 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_500 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_500 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_500 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_500 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_500 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_500 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_500 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_500 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_500 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_500 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_500 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_500 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_500 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_500 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_500 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_500 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_500 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_500 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_500 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_501;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_501 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_501 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_501 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_501 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_501 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_501 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_501 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_501 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_501 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_501 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_501 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_501 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_501 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_501 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_501 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_501 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_501 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_501 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_501 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_501 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_501 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_501 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_501 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_501 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_501 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_501 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_501 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_501 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_501 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_501 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_501 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_501 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_502;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_502 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_502 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_502 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_502 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_502 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_502 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_502 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_502 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_502 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_502 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_502 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_502 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_502 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_502 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_502 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_502 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_502 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_502 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_502 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_502 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_502 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_502 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_502 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_502 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_502 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_502 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_502 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_502 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_502 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_502 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_502 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_502 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_503;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_503 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_503 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_503 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_503 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_503 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_503 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_503 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_503 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_503 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_503 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_503 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_503 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_503 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_503 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_503 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_503 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_503 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_503 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_503 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_503 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_503 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_503 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_503 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_503 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_503 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_503 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_503 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_503 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_503 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_503 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_503 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_503 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_504;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_504 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_504 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_504 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_504 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_504 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_504 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_504 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_504 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_504 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_504 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_504 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_504 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_504 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_504 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_504 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_504 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_504 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_504 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_504 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_504 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_504 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_504 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_504 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_504 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_504 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_504 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_504 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_504 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_504 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_504 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_504 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_504 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  wire        send_iresp_1 = casez_tmp_503 == 2'h0;
  wire        send_fresp_1 = casez_tmp_503 == 2'h1;
  reg  [6:0]  casez_tmp_505;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_505 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_505 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_505 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_505 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_505 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_505 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_505 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_505 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_505 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_505 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_505 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_505 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_505 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_505 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_505 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_505 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_505 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_505 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_505 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_505 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_505 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_505 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_505 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_505 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_505 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_505 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_505 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_505 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_505 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_505 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_505 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_505 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_506;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_506 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_506 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_506 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_506 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_506 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_506 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_506 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_506 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_506 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_506 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_506 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_506 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_506 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_506 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_506 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_506 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_506 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_506 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_506 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_506 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_506 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_506 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_506 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_506 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_506 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_506 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_506 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_506 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_506 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_506 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_506 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_506 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_507;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_507 = stq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_507 = stq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_507 = stq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_507 = stq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_507 = stq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_507 = stq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_507 = stq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_507 = stq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_507 = stq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_507 = stq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_507 = stq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_507 = stq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_507 = stq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_507 = stq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_507 = stq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_507 = stq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_507 = stq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_507 = stq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_507 = stq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_507 = stq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_507 = stq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_507 = stq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_507 = stq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_507 = stq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_507 = stq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_507 = stq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_507 = stq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_507 = stq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_507 = stq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_507 = stq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_507 = stq_30_bits_uop_pdst;
      default:
        casez_tmp_507 = stq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_508;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_508 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_508 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_508 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_508 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_508 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_508 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_508 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_508 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_508 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_508 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_508 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_508 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_508 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_508 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_508 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_508 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_508 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_508 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_508 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_508 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_508 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_508 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_508 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_508 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_508 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_508 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_508 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_508 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_508 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_508 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_508 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_508 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_509;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_509 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_509 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_509 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_509 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_509 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_509 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_509 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_509 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_509 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_509 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_509 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_509 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_509 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_509 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_509 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_509 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_509 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_509 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_509 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_509 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_509 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_509 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_509 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_509 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_509 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_509 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_509 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_509 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_509 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_509 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_509 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_509 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_510;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_510 = stq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_510 = stq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_510 = stq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_510 = stq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_510 = stq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_510 = stq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_510 = stq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_510 = stq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_510 = stq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_510 = stq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_510 = stq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_510 = stq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_510 = stq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_510 = stq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_510 = stq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_510 = stq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_510 = stq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_510 = stq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_510 = stq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_510 = stq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_510 = stq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_510 = stq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_510 = stq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_510 = stq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_510 = stq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_510 = stq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_510 = stq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_510 = stq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_510 = stq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_510 = stq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_510 = stq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_510 = stq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  wire        _GEN_1507 = io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_is_amo;
  wire        dmem_resp_fired_1 = io_dmem_resp_1_valid & (io_dmem_resp_1_bits_uop_uses_ldq | _GEN_1507);
  wire        _GEN_1508 = dmem_resp_fired_1 & wb_forward_valid_1;
  wire        _GEN_1509 = ~dmem_resp_fired_1 & wb_forward_valid_1;
  reg  [6:0]  casez_tmp_511;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_511 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_511 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_511 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_511 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_511 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_511 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_511 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_511 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_511 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_511 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_511 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_511 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_511 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_511 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_511 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_511 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_511 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_511 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_511 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_511 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_511 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_511 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_511 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_511 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_511 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_511 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_511 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_511 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_511 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_511 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_511 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_511 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  reg  [19:0] casez_tmp_512;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_512 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_512 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_512 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_512 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_512 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_512 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_512 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_512 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_512 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_512 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_512 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_512 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_512 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_512 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_512 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_512 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_512 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_512 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_512 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_512 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_512 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_512 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_512 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_512 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_512 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_512 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_512 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_512 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_512 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_512 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_512 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_512 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_513;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_513 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_513 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_513 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_513 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_513 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_513 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_513 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_513 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_513 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_513 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_513 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_513 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_513 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_513 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_513 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_513 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_513 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_513 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_513 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_513 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_513 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_513 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_513 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_513 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_513 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_513 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_513 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_513 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_513 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_513 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_513 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_513 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_514;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_514 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_514 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_514 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_514 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_514 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_514 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_514 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_514 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_514 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_514 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_514 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_514 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_514 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_514 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_514 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_514 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_514 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_514 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_514 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_514 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_514 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_514 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_514 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_514 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_514 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_514 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_514 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_514 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_514 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_514 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_514 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_514 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  reg  [4:0]  casez_tmp_515;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_515 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_515 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_515 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_515 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_515 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_515 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_515 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_515 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_515 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_515 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_515 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_515 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_515 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_515 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_515 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_515 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_515 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_515 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_515 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_515 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_515 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_515 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_515 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_515 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_515 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_515 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_515 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_515 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_515 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_515 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_515 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_515 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_516;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_516 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_516 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_516 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_516 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_516 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_516 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_516 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_516 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_516 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_516 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_516 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_516 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_516 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_516 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_516 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_516 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_516 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_516 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_516 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_516 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_516 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_516 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_516 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_516 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_516 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_516 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_516 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_516 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_516 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_516 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_516 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_516 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_517;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_517 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_517 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_517 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_517 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_517 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_517 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_517 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_517 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_517 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_517 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_517 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_517 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_517 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_517 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_517 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_517 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_517 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_517 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_517 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_517 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_517 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_517 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_517 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_517 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_517 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_517 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_517 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_517 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_517 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_517 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_517 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_517 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_518;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_518 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_518 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_518 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_518 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_518 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_518 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_518 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_518 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_518 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_518 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_518 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_518 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_518 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_518 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_518 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_518 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_518 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_518 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_518 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_518 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_518 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_518 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_518 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_518 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_518 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_518 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_518 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_518 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_518 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_518 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_518 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_518 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  reg         casez_tmp_519;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_519 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_519 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_519 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_519 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_519 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_519 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_519 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_519 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_519 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_519 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_519 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_519 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_519 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_519 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_519 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_519 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_519 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_519 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_519 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_519 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_519 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_519 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_519 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_519 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_519 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_519 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_519 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_519 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_519 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_519 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_519 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_519 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         casez_tmp_520;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_520 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_520 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_520 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_520 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_520 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_520 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_520 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_520 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_520 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_520 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_520 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_520 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_520 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_520 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_520 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_520 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_520 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_520 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_520 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_520 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_520 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_520 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_520 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_520 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_520 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_520 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_520 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_520 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_520 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_520 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_520 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_520 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_521;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_521 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_521 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_521 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_521 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_521 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_521 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_521 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_521 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_521 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_521 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_521 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_521 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_521 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_521 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_521 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_521 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_521 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_521 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_521 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_521 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_521 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_521 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_521 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_521 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_521 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_521 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_521 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_521 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_521 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_521 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_521 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_521 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_522;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_522 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_522 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_522 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_522 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_522 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_522 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_522 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_522 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_522 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_522 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_522 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_522 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_522 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_522 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_522 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_522 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_522 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_522 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_522 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_522 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_522 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_522 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_522 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_522 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_522 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_522 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_522 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_522 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_522 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_522 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_522 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_522 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  wire        live_1 = (io_core_brupdate_b1_mispredict_mask & casez_tmp_512) == 20'h0;
  reg  [1:0]  casez_tmp_523;
  always @(*) begin
    casez (wb_forward_stq_idx_1)
      5'b00000:
        casez_tmp_523 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_523 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_523 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_523 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_523 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_523 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_523 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_523 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_523 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_523 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_523 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_523 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_523 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_523 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_523 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_523 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_523 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_523 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_523 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_523 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_523 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_523 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_523 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_523 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_523 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_523 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_523 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_523 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_523 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_523 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_523 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_523 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  reg         casez_tmp_524;
  always @(*) begin
    casez (wb_forward_stq_idx_1)
      5'b00000:
        casez_tmp_524 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_524 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_524 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_524 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_524 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_524 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_524 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_524 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_524 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_524 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_524 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_524 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_524 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_524 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_524 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_524 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_524 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_524 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_524 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_524 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_524 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_524 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_524 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_524 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_524 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_524 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_524 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_524 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_524 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_524 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_524 = stq_30_bits_data_valid;
      default:
        casez_tmp_524 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_525;
  always @(*) begin
    casez (wb_forward_stq_idx_1)
      5'b00000:
        casez_tmp_525 = stq_0_bits_data_bits;
      5'b00001:
        casez_tmp_525 = stq_1_bits_data_bits;
      5'b00010:
        casez_tmp_525 = stq_2_bits_data_bits;
      5'b00011:
        casez_tmp_525 = stq_3_bits_data_bits;
      5'b00100:
        casez_tmp_525 = stq_4_bits_data_bits;
      5'b00101:
        casez_tmp_525 = stq_5_bits_data_bits;
      5'b00110:
        casez_tmp_525 = stq_6_bits_data_bits;
      5'b00111:
        casez_tmp_525 = stq_7_bits_data_bits;
      5'b01000:
        casez_tmp_525 = stq_8_bits_data_bits;
      5'b01001:
        casez_tmp_525 = stq_9_bits_data_bits;
      5'b01010:
        casez_tmp_525 = stq_10_bits_data_bits;
      5'b01011:
        casez_tmp_525 = stq_11_bits_data_bits;
      5'b01100:
        casez_tmp_525 = stq_12_bits_data_bits;
      5'b01101:
        casez_tmp_525 = stq_13_bits_data_bits;
      5'b01110:
        casez_tmp_525 = stq_14_bits_data_bits;
      5'b01111:
        casez_tmp_525 = stq_15_bits_data_bits;
      5'b10000:
        casez_tmp_525 = stq_16_bits_data_bits;
      5'b10001:
        casez_tmp_525 = stq_17_bits_data_bits;
      5'b10010:
        casez_tmp_525 = stq_18_bits_data_bits;
      5'b10011:
        casez_tmp_525 = stq_19_bits_data_bits;
      5'b10100:
        casez_tmp_525 = stq_20_bits_data_bits;
      5'b10101:
        casez_tmp_525 = stq_21_bits_data_bits;
      5'b10110:
        casez_tmp_525 = stq_22_bits_data_bits;
      5'b10111:
        casez_tmp_525 = stq_23_bits_data_bits;
      5'b11000:
        casez_tmp_525 = stq_24_bits_data_bits;
      5'b11001:
        casez_tmp_525 = stq_25_bits_data_bits;
      5'b11010:
        casez_tmp_525 = stq_26_bits_data_bits;
      5'b11011:
        casez_tmp_525 = stq_27_bits_data_bits;
      5'b11100:
        casez_tmp_525 = stq_28_bits_data_bits;
      5'b11101:
        casez_tmp_525 = stq_29_bits_data_bits;
      5'b11110:
        casez_tmp_525 = stq_30_bits_data_bits;
      default:
        casez_tmp_525 = stq_31_bits_data_bits;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_526;
  always @(*) begin
    casez (casez_tmp_523)
      2'b00:
        casez_tmp_526 = {2{{2{{2{casez_tmp_525[7:0]}}}}}};
      2'b01:
        casez_tmp_526 = {2{{2{casez_tmp_525[15:0]}}}};
      2'b10:
        casez_tmp_526 = {2{casez_tmp_525[31:0]}};
      default:
        casez_tmp_526 = casez_tmp_525;
    endcase
  end // always @(*)
  wire        _GEN_1510 = _GEN_1508 | ~_GEN_1509;
  wire        _io_core_exe_1_iresp_valid_output = _GEN_1510 ? io_dmem_resp_1_valid & (io_dmem_resp_1_bits_uop_uses_ldq ? send_iresp_1 : _GEN_1507) : casez_tmp_521 == 2'h0 & casez_tmp_524 & live_1;
  wire        _io_core_exe_1_fresp_valid_output = _GEN_1510 ? _GEN_1506 & send_fresp_1 : casez_tmp_521 == 2'h1 & casez_tmp_524 & live_1;
  wire [31:0] io_core_exe_1_iresp_bits_data_zeroed = wb_forward_ld_addr_1[2] ? casez_tmp_526[63:32] : casez_tmp_526[31:0];
  wire        _ldq_bits_debug_wb_data_T_28 = casez_tmp_517 == 2'h2;
  wire [15:0] io_core_exe_1_iresp_bits_data_zeroed_1 = wb_forward_ld_addr_1[1] ? io_core_exe_1_iresp_bits_data_zeroed[31:16] : io_core_exe_1_iresp_bits_data_zeroed[15:0];
  wire        _ldq_bits_debug_wb_data_T_37 = casez_tmp_517 == 2'h1;
  wire [7:0]  io_core_exe_1_iresp_bits_data_zeroed_2 = wb_forward_ld_addr_1[0] ? io_core_exe_1_iresp_bits_data_zeroed_1[15:8] : io_core_exe_1_iresp_bits_data_zeroed_1[7:0];
  wire        _ldq_bits_debug_wb_data_T_46 = casez_tmp_517 == 2'h0;
  wire [31:0] io_core_exe_1_fresp_bits_data_zeroed = wb_forward_ld_addr_1[2] ? casez_tmp_526[63:32] : casez_tmp_526[31:0];
  wire [15:0] io_core_exe_1_fresp_bits_data_zeroed_1 = wb_forward_ld_addr_1[1] ? io_core_exe_1_fresp_bits_data_zeroed[31:16] : io_core_exe_1_fresp_bits_data_zeroed[15:0];
  wire [7:0]  io_core_exe_1_fresp_bits_data_zeroed_2 = wb_forward_ld_addr_1[0] ? io_core_exe_1_fresp_bits_data_zeroed_1[15:8] : io_core_exe_1_fresp_bits_data_zeroed_1[7:0];
  reg         io_core_ld_miss_REG;
  reg         spec_ld_succeed_REG;
  reg  [4:0]  spec_ld_succeed_REG_1;
  reg         spec_ld_succeed_REG_2;
  reg  [4:0]  spec_ld_succeed_REG_3;
  wire [19:0] _GEN_1511 = io_core_brupdate_b1_mispredict_mask & stq_0_bits_uop_br_mask;
  wire [19:0] _GEN_1512 = io_core_brupdate_b1_mispredict_mask & stq_1_bits_uop_br_mask;
  wire [19:0] _GEN_1513 = io_core_brupdate_b1_mispredict_mask & stq_2_bits_uop_br_mask;
  wire [19:0] _GEN_1514 = io_core_brupdate_b1_mispredict_mask & stq_3_bits_uop_br_mask;
  wire [19:0] _GEN_1515 = io_core_brupdate_b1_mispredict_mask & stq_4_bits_uop_br_mask;
  wire [19:0] _GEN_1516 = io_core_brupdate_b1_mispredict_mask & stq_5_bits_uop_br_mask;
  wire [19:0] _GEN_1517 = io_core_brupdate_b1_mispredict_mask & stq_6_bits_uop_br_mask;
  wire [19:0] _GEN_1518 = io_core_brupdate_b1_mispredict_mask & stq_7_bits_uop_br_mask;
  wire [19:0] _GEN_1519 = io_core_brupdate_b1_mispredict_mask & stq_8_bits_uop_br_mask;
  wire [19:0] _GEN_1520 = io_core_brupdate_b1_mispredict_mask & stq_9_bits_uop_br_mask;
  wire [19:0] _GEN_1521 = io_core_brupdate_b1_mispredict_mask & stq_10_bits_uop_br_mask;
  wire [19:0] _GEN_1522 = io_core_brupdate_b1_mispredict_mask & stq_11_bits_uop_br_mask;
  wire [19:0] _GEN_1523 = io_core_brupdate_b1_mispredict_mask & stq_12_bits_uop_br_mask;
  wire [19:0] _GEN_1524 = io_core_brupdate_b1_mispredict_mask & stq_13_bits_uop_br_mask;
  wire [19:0] _GEN_1525 = io_core_brupdate_b1_mispredict_mask & stq_14_bits_uop_br_mask;
  wire [19:0] _GEN_1526 = io_core_brupdate_b1_mispredict_mask & stq_15_bits_uop_br_mask;
  wire [19:0] _GEN_1527 = io_core_brupdate_b1_mispredict_mask & stq_16_bits_uop_br_mask;
  wire [19:0] _GEN_1528 = io_core_brupdate_b1_mispredict_mask & stq_17_bits_uop_br_mask;
  wire [19:0] _GEN_1529 = io_core_brupdate_b1_mispredict_mask & stq_18_bits_uop_br_mask;
  wire [19:0] _GEN_1530 = io_core_brupdate_b1_mispredict_mask & stq_19_bits_uop_br_mask;
  wire [19:0] _GEN_1531 = io_core_brupdate_b1_mispredict_mask & stq_20_bits_uop_br_mask;
  wire [19:0] _GEN_1532 = io_core_brupdate_b1_mispredict_mask & stq_21_bits_uop_br_mask;
  wire [19:0] _GEN_1533 = io_core_brupdate_b1_mispredict_mask & stq_22_bits_uop_br_mask;
  wire [19:0] _GEN_1534 = io_core_brupdate_b1_mispredict_mask & stq_23_bits_uop_br_mask;
  wire [19:0] _GEN_1535 = io_core_brupdate_b1_mispredict_mask & stq_24_bits_uop_br_mask;
  wire [19:0] _GEN_1536 = io_core_brupdate_b1_mispredict_mask & stq_25_bits_uop_br_mask;
  wire [19:0] _GEN_1537 = io_core_brupdate_b1_mispredict_mask & stq_26_bits_uop_br_mask;
  wire [19:0] _GEN_1538 = io_core_brupdate_b1_mispredict_mask & stq_27_bits_uop_br_mask;
  wire [19:0] _GEN_1539 = io_core_brupdate_b1_mispredict_mask & stq_28_bits_uop_br_mask;
  wire [19:0] _GEN_1540 = io_core_brupdate_b1_mispredict_mask & stq_29_bits_uop_br_mask;
  wire [19:0] _GEN_1541 = io_core_brupdate_b1_mispredict_mask & stq_30_bits_uop_br_mask;
  wire [19:0] _GEN_1542 = io_core_brupdate_b1_mispredict_mask & stq_31_bits_uop_br_mask;
  wire        commit_store = io_core_commit_valids_0 & io_core_commit_uops_0_uses_stq;
  wire        commit_load = io_core_commit_valids_0 & io_core_commit_uops_0_uses_ldq;
  wire [4:0]  idx = commit_store ? stq_commit_head : ldq_head;
  wire        _GEN_1543 = ~commit_store & commit_load & ~reset;
  reg         casez_tmp_527;
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_527 = ldq_0_valid;
      5'b00001:
        casez_tmp_527 = ldq_1_valid;
      5'b00010:
        casez_tmp_527 = ldq_2_valid;
      5'b00011:
        casez_tmp_527 = ldq_3_valid;
      5'b00100:
        casez_tmp_527 = ldq_4_valid;
      5'b00101:
        casez_tmp_527 = ldq_5_valid;
      5'b00110:
        casez_tmp_527 = ldq_6_valid;
      5'b00111:
        casez_tmp_527 = ldq_7_valid;
      5'b01000:
        casez_tmp_527 = ldq_8_valid;
      5'b01001:
        casez_tmp_527 = ldq_9_valid;
      5'b01010:
        casez_tmp_527 = ldq_10_valid;
      5'b01011:
        casez_tmp_527 = ldq_11_valid;
      5'b01100:
        casez_tmp_527 = ldq_12_valid;
      5'b01101:
        casez_tmp_527 = ldq_13_valid;
      5'b01110:
        casez_tmp_527 = ldq_14_valid;
      5'b01111:
        casez_tmp_527 = ldq_15_valid;
      5'b10000:
        casez_tmp_527 = ldq_16_valid;
      5'b10001:
        casez_tmp_527 = ldq_17_valid;
      5'b10010:
        casez_tmp_527 = ldq_18_valid;
      5'b10011:
        casez_tmp_527 = ldq_19_valid;
      5'b10100:
        casez_tmp_527 = ldq_20_valid;
      5'b10101:
        casez_tmp_527 = ldq_21_valid;
      5'b10110:
        casez_tmp_527 = ldq_22_valid;
      5'b10111:
        casez_tmp_527 = ldq_23_valid;
      5'b11000:
        casez_tmp_527 = ldq_24_valid;
      5'b11001:
        casez_tmp_527 = ldq_25_valid;
      5'b11010:
        casez_tmp_527 = ldq_26_valid;
      5'b11011:
        casez_tmp_527 = ldq_27_valid;
      5'b11100:
        casez_tmp_527 = ldq_28_valid;
      5'b11101:
        casez_tmp_527 = ldq_29_valid;
      5'b11110:
        casez_tmp_527 = ldq_30_valid;
      default:
        casez_tmp_527 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_528;
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_528 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_528 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_528 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_528 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_528 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_528 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_528 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_528 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_528 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_528 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_528 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_528 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_528 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_528 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_528 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_528 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_528 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_528 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_528 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_528 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_528 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_528 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_528 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_528 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_528 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_528 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_528 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_528 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_528 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_528 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_528 = ldq_30_bits_executed;
      default:
        casez_tmp_528 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg         casez_tmp_529;
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_529 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_529 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_529 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_529 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_529 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_529 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_529 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_529 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_529 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_529 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_529 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_529 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_529 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_529 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_529 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_529 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_529 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_529 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_529 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_529 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_529 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_529 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_529 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_529 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_529 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_529 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_529 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_529 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_529 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_529 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_529 = ldq_30_bits_succeeded;
      default:
        casez_tmp_529 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  reg         casez_tmp_530;
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_530 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_530 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_530 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_530 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_530 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_530 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_530 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_530 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_530 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_530 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_530 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_530 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_530 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_530 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_530 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_530 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_530 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_530 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_530 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_530 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_530 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_530 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_530 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_530 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_530 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_530 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_530 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_530 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_530 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_530 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_530 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_530 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  wire [4:0]  _GEN_1544 = stq_commit_head + 5'h1;
  wire [4:0]  _GEN_1545 = commit_store ? _GEN_1544 : stq_commit_head;
  wire [4:0]  _GEN_1546 = ldq_head + 5'h1;
  wire [4:0]  _GEN_1547 = commit_load ? _GEN_1546 : ldq_head;
  wire        commit_store_1 = io_core_commit_valids_1 & io_core_commit_uops_1_uses_stq;
  wire        commit_load_1 = io_core_commit_valids_1 & io_core_commit_uops_1_uses_ldq;
  wire [4:0]  idx_1 = commit_store_1 ? _GEN_1545 : _GEN_1547;
  wire        _GEN_1548 = ~commit_store_1 & commit_load_1 & ~reset;
  reg         casez_tmp_531;
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_531 = ldq_0_valid;
      5'b00001:
        casez_tmp_531 = ldq_1_valid;
      5'b00010:
        casez_tmp_531 = ldq_2_valid;
      5'b00011:
        casez_tmp_531 = ldq_3_valid;
      5'b00100:
        casez_tmp_531 = ldq_4_valid;
      5'b00101:
        casez_tmp_531 = ldq_5_valid;
      5'b00110:
        casez_tmp_531 = ldq_6_valid;
      5'b00111:
        casez_tmp_531 = ldq_7_valid;
      5'b01000:
        casez_tmp_531 = ldq_8_valid;
      5'b01001:
        casez_tmp_531 = ldq_9_valid;
      5'b01010:
        casez_tmp_531 = ldq_10_valid;
      5'b01011:
        casez_tmp_531 = ldq_11_valid;
      5'b01100:
        casez_tmp_531 = ldq_12_valid;
      5'b01101:
        casez_tmp_531 = ldq_13_valid;
      5'b01110:
        casez_tmp_531 = ldq_14_valid;
      5'b01111:
        casez_tmp_531 = ldq_15_valid;
      5'b10000:
        casez_tmp_531 = ldq_16_valid;
      5'b10001:
        casez_tmp_531 = ldq_17_valid;
      5'b10010:
        casez_tmp_531 = ldq_18_valid;
      5'b10011:
        casez_tmp_531 = ldq_19_valid;
      5'b10100:
        casez_tmp_531 = ldq_20_valid;
      5'b10101:
        casez_tmp_531 = ldq_21_valid;
      5'b10110:
        casez_tmp_531 = ldq_22_valid;
      5'b10111:
        casez_tmp_531 = ldq_23_valid;
      5'b11000:
        casez_tmp_531 = ldq_24_valid;
      5'b11001:
        casez_tmp_531 = ldq_25_valid;
      5'b11010:
        casez_tmp_531 = ldq_26_valid;
      5'b11011:
        casez_tmp_531 = ldq_27_valid;
      5'b11100:
        casez_tmp_531 = ldq_28_valid;
      5'b11101:
        casez_tmp_531 = ldq_29_valid;
      5'b11110:
        casez_tmp_531 = ldq_30_valid;
      default:
        casez_tmp_531 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_532;
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_532 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_532 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_532 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_532 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_532 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_532 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_532 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_532 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_532 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_532 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_532 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_532 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_532 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_532 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_532 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_532 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_532 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_532 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_532 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_532 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_532 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_532 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_532 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_532 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_532 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_532 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_532 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_532 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_532 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_532 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_532 = ldq_30_bits_executed;
      default:
        casez_tmp_532 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg         casez_tmp_533;
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_533 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_533 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_533 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_533 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_533 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_533 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_533 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_533 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_533 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_533 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_533 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_533 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_533 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_533 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_533 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_533 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_533 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_533 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_533 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_533 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_533 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_533 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_533 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_533 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_533 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_533 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_533 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_533 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_533 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_533 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_533 = ldq_30_bits_succeeded;
      default:
        casez_tmp_533 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  reg         casez_tmp_534;
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_534 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_534 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_534 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_534 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_534 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_534 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_534 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_534 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_534 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_534 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_534 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_534 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_534 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_534 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_534 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_534 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_534 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_534 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_534 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_534 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_534 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_534 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_534 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_534 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_534 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_534 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_534 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_534 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_534 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_534 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_534 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_534 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  wire [4:0]  _GEN_1549 = _GEN_1545 + 5'h1;
  wire [4:0]  _GEN_1550 = commit_store_1 ? _GEN_1549 : _GEN_1545;
  wire [4:0]  _GEN_1551 = _GEN_1547 + 5'h1;
  wire [4:0]  _GEN_1552 = commit_load_1 ? _GEN_1551 : _GEN_1547;
  wire        commit_store_2 = io_core_commit_valids_2 & io_core_commit_uops_2_uses_stq;
  wire        commit_load_2 = io_core_commit_valids_2 & io_core_commit_uops_2_uses_ldq;
  wire [4:0]  idx_2 = commit_store_2 ? _GEN_1550 : _GEN_1552;
  wire        _GEN_1553 = ~commit_store_2 & commit_load_2 & ~reset;
  reg         casez_tmp_535;
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_535 = ldq_0_valid;
      5'b00001:
        casez_tmp_535 = ldq_1_valid;
      5'b00010:
        casez_tmp_535 = ldq_2_valid;
      5'b00011:
        casez_tmp_535 = ldq_3_valid;
      5'b00100:
        casez_tmp_535 = ldq_4_valid;
      5'b00101:
        casez_tmp_535 = ldq_5_valid;
      5'b00110:
        casez_tmp_535 = ldq_6_valid;
      5'b00111:
        casez_tmp_535 = ldq_7_valid;
      5'b01000:
        casez_tmp_535 = ldq_8_valid;
      5'b01001:
        casez_tmp_535 = ldq_9_valid;
      5'b01010:
        casez_tmp_535 = ldq_10_valid;
      5'b01011:
        casez_tmp_535 = ldq_11_valid;
      5'b01100:
        casez_tmp_535 = ldq_12_valid;
      5'b01101:
        casez_tmp_535 = ldq_13_valid;
      5'b01110:
        casez_tmp_535 = ldq_14_valid;
      5'b01111:
        casez_tmp_535 = ldq_15_valid;
      5'b10000:
        casez_tmp_535 = ldq_16_valid;
      5'b10001:
        casez_tmp_535 = ldq_17_valid;
      5'b10010:
        casez_tmp_535 = ldq_18_valid;
      5'b10011:
        casez_tmp_535 = ldq_19_valid;
      5'b10100:
        casez_tmp_535 = ldq_20_valid;
      5'b10101:
        casez_tmp_535 = ldq_21_valid;
      5'b10110:
        casez_tmp_535 = ldq_22_valid;
      5'b10111:
        casez_tmp_535 = ldq_23_valid;
      5'b11000:
        casez_tmp_535 = ldq_24_valid;
      5'b11001:
        casez_tmp_535 = ldq_25_valid;
      5'b11010:
        casez_tmp_535 = ldq_26_valid;
      5'b11011:
        casez_tmp_535 = ldq_27_valid;
      5'b11100:
        casez_tmp_535 = ldq_28_valid;
      5'b11101:
        casez_tmp_535 = ldq_29_valid;
      5'b11110:
        casez_tmp_535 = ldq_30_valid;
      default:
        casez_tmp_535 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_536;
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_536 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_536 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_536 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_536 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_536 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_536 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_536 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_536 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_536 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_536 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_536 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_536 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_536 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_536 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_536 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_536 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_536 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_536 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_536 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_536 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_536 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_536 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_536 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_536 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_536 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_536 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_536 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_536 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_536 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_536 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_536 = ldq_30_bits_executed;
      default:
        casez_tmp_536 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg         casez_tmp_537;
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_537 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_537 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_537 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_537 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_537 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_537 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_537 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_537 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_537 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_537 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_537 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_537 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_537 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_537 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_537 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_537 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_537 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_537 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_537 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_537 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_537 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_537 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_537 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_537 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_537 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_537 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_537 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_537 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_537 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_537 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_537 = ldq_30_bits_succeeded;
      default:
        casez_tmp_537 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  reg         casez_tmp_538;
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_538 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_538 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_538 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_538 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_538 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_538 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_538 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_538 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_538 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_538 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_538 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_538 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_538 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_538 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_538 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_538 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_538 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_538 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_538 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_538 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_538 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_538 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_538 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_538 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_538 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_538 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_538 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_538 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_538 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_538 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_538 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_538 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  wire [4:0]  _GEN_1554 = _GEN_1550 + 5'h1;
  wire [4:0]  _GEN_1555 = commit_store_2 ? _GEN_1554 : _GEN_1550;
  wire [4:0]  _GEN_1556 = _GEN_1552 + 5'h1;
  wire [4:0]  _GEN_1557 = commit_load_2 ? _GEN_1556 : _GEN_1552;
  wire        commit_store_3 = io_core_commit_valids_3 & io_core_commit_uops_3_uses_stq;
  wire        commit_load_3 = io_core_commit_valids_3 & io_core_commit_uops_3_uses_ldq;
  wire [4:0]  idx_3 = commit_store_3 ? _GEN_1555 : _GEN_1557;
  wire        _GEN_1558 = ~commit_store_3 & commit_load_3 & ~reset;
  reg         casez_tmp_539;
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_539 = ldq_0_valid;
      5'b00001:
        casez_tmp_539 = ldq_1_valid;
      5'b00010:
        casez_tmp_539 = ldq_2_valid;
      5'b00011:
        casez_tmp_539 = ldq_3_valid;
      5'b00100:
        casez_tmp_539 = ldq_4_valid;
      5'b00101:
        casez_tmp_539 = ldq_5_valid;
      5'b00110:
        casez_tmp_539 = ldq_6_valid;
      5'b00111:
        casez_tmp_539 = ldq_7_valid;
      5'b01000:
        casez_tmp_539 = ldq_8_valid;
      5'b01001:
        casez_tmp_539 = ldq_9_valid;
      5'b01010:
        casez_tmp_539 = ldq_10_valid;
      5'b01011:
        casez_tmp_539 = ldq_11_valid;
      5'b01100:
        casez_tmp_539 = ldq_12_valid;
      5'b01101:
        casez_tmp_539 = ldq_13_valid;
      5'b01110:
        casez_tmp_539 = ldq_14_valid;
      5'b01111:
        casez_tmp_539 = ldq_15_valid;
      5'b10000:
        casez_tmp_539 = ldq_16_valid;
      5'b10001:
        casez_tmp_539 = ldq_17_valid;
      5'b10010:
        casez_tmp_539 = ldq_18_valid;
      5'b10011:
        casez_tmp_539 = ldq_19_valid;
      5'b10100:
        casez_tmp_539 = ldq_20_valid;
      5'b10101:
        casez_tmp_539 = ldq_21_valid;
      5'b10110:
        casez_tmp_539 = ldq_22_valid;
      5'b10111:
        casez_tmp_539 = ldq_23_valid;
      5'b11000:
        casez_tmp_539 = ldq_24_valid;
      5'b11001:
        casez_tmp_539 = ldq_25_valid;
      5'b11010:
        casez_tmp_539 = ldq_26_valid;
      5'b11011:
        casez_tmp_539 = ldq_27_valid;
      5'b11100:
        casez_tmp_539 = ldq_28_valid;
      5'b11101:
        casez_tmp_539 = ldq_29_valid;
      5'b11110:
        casez_tmp_539 = ldq_30_valid;
      default:
        casez_tmp_539 = ldq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_540;
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_540 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_540 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_540 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_540 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_540 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_540 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_540 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_540 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_540 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_540 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_540 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_540 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_540 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_540 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_540 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_540 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_540 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_540 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_540 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_540 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_540 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_540 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_540 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_540 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_540 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_540 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_540 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_540 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_540 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_540 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_540 = ldq_30_bits_executed;
      default:
        casez_tmp_540 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  reg         casez_tmp_541;
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_541 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_541 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_541 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_541 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_541 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_541 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_541 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_541 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_541 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_541 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_541 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_541 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_541 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_541 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_541 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_541 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_541 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_541 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_541 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_541 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_541 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_541 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_541 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_541 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_541 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_541 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_541 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_541 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_541 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_541 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_541 = ldq_30_bits_succeeded;
      default:
        casez_tmp_541 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  reg         casez_tmp_542;
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_542 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_542 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_542 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_542 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_542 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_542 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_542 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_542 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_542 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_542 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_542 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_542 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_542 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_542 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_542 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_542 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_542 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_542 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_542 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_542 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_542 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_542 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_542 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_542 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_542 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_542 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_542 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_542 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_542 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_542 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_542 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_542 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  `ifndef SYNTHESIS
    wire _GEN_1559 = dis_ld_val & ~reset;
    wire _GEN_1560 = ~dis_ld_val & dis_st_val & ~reset;
    wire _GEN_1561 = dis_ld_val_1 & ~reset;
    wire _GEN_1562 = ~dis_ld_val_1 & dis_st_val_1 & ~reset;
    wire _GEN_1563 = dis_ld_val_2 & ~reset;
    wire _GEN_1564 = ~dis_ld_val_2 & dis_st_val_2 & ~reset;
    wire _GEN_1565 = dis_ld_val_3 & ~reset;
    wire _GEN_1566 = ~dis_ld_val_3 & dis_st_val_3 & ~reset;
    wire _GEN_1567 = mem_xcpt_valids_0 & ~reset;
    wire _GEN_1568 = mem_xcpt_valids_1 & ~reset;
    wire _GEN_1569 = ~will_fire_load_incoming_0_will_fire & ~will_fire_load_retry_0_will_fire & ~will_fire_store_commit_0_will_fire;
    wire _GEN_1570 = ~casez_tmp_375 & ~casez_tmp_373;
    wire _GEN_1571 = _GEN_1569 & ~will_fire_load_wakeup_0_will_fire;
    wire _GEN_1572 = ~will_fire_load_incoming_1_will_fire & ~will_fire_load_retry_1_will_fire & ~will_fire_store_commit_1_will_fire;
    wire _GEN_1573 = _GEN_1572 & ~will_fire_load_wakeup_1_will_fire;
    wire _GEN_1574 = _GEN_1431 | _GEN_1432;
    wire _GEN_1575 = _GEN_1466 & ~reset;
    wire _GEN_1576 = _GEN_1506 & ~reset;
    always @(posedge clock) begin
      if (~reset & ~(io_core_brupdate_b2_mispredict | casez_tmp | stq_head == stq_execute_head | stq_tail == stq_execute_head)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: stq_execute_head got off track.\n    at lsu.scala:222 assert (io.core.brupdate.b2.mispredict ||\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1559 & ldq_tail != io_core_dis_uops_0_bits_ldq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1559 & casez_tmp_85) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1560 & stq_tail != io_core_dis_uops_0_bits_stq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1560 & casez_tmp_86) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & dis_ld_val & dis_st_val) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1561 & _GEN_5 != io_core_dis_uops_1_bits_ldq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1561 & casez_tmp_87) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1562 & _GEN_6 != io_core_dis_uops_1_bits_stq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1562 & casez_tmp_88) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & dis_ld_val_1 & dis_st_val_1) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1563 & _GEN_9 != io_core_dis_uops_2_bits_ldq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1563 & casez_tmp_89) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1564 & _GEN_10 != io_core_dis_uops_2_bits_stq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1564 & casez_tmp_90) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & dis_ld_val_2 & dis_st_val_2) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1565 & _GEN_13 != io_core_dis_uops_3_bits_ldq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1565 & casez_tmp_91) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1566 & _GEN_14 != io_core_dis_uops_3_bits_stq_idx) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1566 & casez_tmp_92) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & dis_ld_val_3 & dis_st_val_3) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & exe_req_0_valid & ~(_GEN_18 | will_fire_std_incoming_0_will_fire | will_fire_sfence_0_will_fire)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:566 assert(!(exe_req(w).valid && !(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) || will_fire_std_incoming(w) || will_fire_sfence(w))))\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & exe_req_1_valid & ~(_GEN_144 | will_fire_std_incoming_1_will_fire | will_fire_sfence_1_will_fire)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:566 assert(!(exe_req(w).valid && !(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) || will_fire_std_incoming(w) || will_fire_sfence(w))))\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & ~(~((will_fire_sfence_0_will_fire | will_fire_sfence_1_will_fire) & ~(will_fire_sfence_0_will_fire & will_fire_sfence_1_will_fire)) & ~(will_fire_hella_incoming_0_will_fire & will_fire_hella_incoming_1_will_fire) & ~(will_fire_hella_wakeup_0_will_fire & will_fire_hella_wakeup_1_will_fire) & ~(will_fire_load_retry_0_will_fire & will_fire_load_retry_1_will_fire) & ~(will_fire_sta_retry_0_will_fire & will_fire_sta_retry_1_will_fire) & ~(will_fire_store_commit_0_will_fire & will_fire_store_commit_1_will_fire) & ~(will_fire_load_wakeup_0_will_fire & will_fire_load_wakeup_1_will_fire))) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Some operations is proceeding down multiple pipes\n    at lsu.scala:577 assert((memWidth == 1).B ||\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & ~_will_fire_store_commit_0_T_2 & exe_tlb_uop_0_is_fence) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Fence is pretending to talk to the TLB\n    at lsu.scala:683 assert (!(dtlb.io.req(w).valid && exe_tlb_uop(w).is_fence), \"Fence is pretending to talk to the TLB\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (will_fire_load_incoming_0_will_fire | will_fire_sta_incoming_0_will_fire | will_fire_stad_incoming_0_will_fire) & exe_req_0_bits_mxcpt_valid & ~_will_fire_store_commit_0_T_2 & ~(exe_tlb_uop_0_ctrl_is_load | exe_tlb_uop_0_ctrl_is_sta)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: A uop that's not a load or store-address is throwing a memory exception.\n    at lsu.scala:684 assert (!((will_fire_load_incoming(w) || will_fire_sta_incoming(w) || will_fire_stad_incoming(w)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & ~_will_fire_store_commit_1_T_2 & exe_tlb_uop_1_is_fence) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Fence is pretending to talk to the TLB\n    at lsu.scala:683 assert (!(dtlb.io.req(w).valid && exe_tlb_uop(w).is_fence), \"Fence is pretending to talk to the TLB\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (will_fire_load_incoming_1_will_fire | will_fire_sta_incoming_1_will_fire | will_fire_stad_incoming_1_will_fire) & exe_req_1_bits_mxcpt_valid & ~_will_fire_store_commit_1_T_2 & ~(exe_tlb_uop_1_ctrl_is_load | exe_tlb_uop_1_ctrl_is_sta)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: A uop that's not a load or store-address is throwing a memory exception.\n    at lsu.scala:684 assert (!((will_fire_load_incoming(w) || will_fire_sta_incoming(w) || will_fire_stad_incoming(w)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & ~(exe_tlb_paddr_0 == _dtlb_io_resp_0_paddr | exe_req_0_bits_sfence_valid)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] paddrs should match.\n    at lsu.scala:715 assert (exe_tlb_paddr(w) === dtlb.io.resp(w).paddr || exe_req(w).bits.sfence.valid, \"[lsu] paddrs should match.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1567 & ~REG) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:719 assert(RegNext(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) ||\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1567 & (mem_xcpt_uops_0_uses_ldq ^ ~mem_xcpt_uops_0_uses_stq)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:722 assert(mem_xcpt_uops(w).uses_ldq ^ mem_xcpt_uops(w).uses_stq)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & ~(exe_tlb_paddr_1 == _dtlb_io_resp_1_paddr | exe_req_1_bits_sfence_valid)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] paddrs should match.\n    at lsu.scala:715 assert (exe_tlb_paddr(w) === dtlb.io.resp(w).paddr || exe_req(w).bits.sfence.valid, \"[lsu] paddrs should match.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1568 & ~REG_1) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:719 assert(RegNext(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) ||\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1568 & (mem_xcpt_uops_1_uses_ldq ^ ~mem_xcpt_uops_1_uses_stq)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:722 assert(mem_xcpt_uops(w).uses_ldq ^ mem_xcpt_uops(w).uses_stq)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (will_fire_load_incoming_0_will_fire & ~reset & casez_tmp_97) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:773 assert(!ldq_incoming_e(w).bits.executed)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~will_fire_load_incoming_0_will_fire & will_fire_load_retry_0_will_fire & ~reset & casez_tmp_204) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:780 assert(!ldq_retry_e.bits.executed)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1569 & will_fire_load_wakeup_0_will_fire & ~reset & ~_GEN_1570) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:802 assert(!ldq_wakeup_e.bits.executed && !ldq_wakeup_e.bits.addr_is_virtual)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1571 & will_fire_hella_incoming_0_will_fire & ~reset & ~_GEN_2) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:804 assert(hella_state === h_s1)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1571 & ~will_fire_hella_incoming_0_will_fire & will_fire_hella_wakeup_0_will_fire & ~reset & ~_GEN_1) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:821 assert(hella_state === h_replay)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_275 & ~reset & will_fire_load_incoming_0_will_fire & casez_tmp_96) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Incoming load is overwriting a valid address\n    at lsu.scala:845 assert(!(will_fire_load_incoming(w) && ldq_incoming_e(w).bits.addr.valid),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_278 & ~reset & will_fire_sta_incoming_0_will_fire & casez_tmp_111) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid address\n    at lsu.scala:859 assert(!(will_fire_sta_incoming(w) && stq_incoming_e(w).bits.addr.valid),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_279 & ~reset & casez_tmp_381) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid data entry\n    at lsu.scala:878 assert(!(stq(sidx).bits.data.valid),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (will_fire_load_incoming_1_will_fire & ~reset & casez_tmp_103) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:773 assert(!ldq_incoming_e(w).bits.executed)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~will_fire_load_incoming_1_will_fire & will_fire_load_retry_1_will_fire & ~reset & casez_tmp_204) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:780 assert(!ldq_retry_e.bits.executed)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1572 & will_fire_load_wakeup_1_will_fire & ~reset & ~_GEN_1570) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:802 assert(!ldq_wakeup_e.bits.executed && !ldq_wakeup_e.bits.addr_is_virtual)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1573 & will_fire_hella_incoming_1_will_fire & ~reset & ~_GEN_2) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:804 assert(hella_state === h_s1)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1573 & ~will_fire_hella_incoming_1_will_fire & will_fire_hella_wakeup_1_will_fire & ~reset & ~_GEN_1) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:821 assert(hella_state === h_replay)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_281 & ~reset & will_fire_load_incoming_1_will_fire & casez_tmp_102) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Incoming load is overwriting a valid address\n    at lsu.scala:845 assert(!(will_fire_load_incoming(w) && ldq_incoming_e(w).bits.addr.valid),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_283 & ~reset & will_fire_sta_incoming_1_will_fire & casez_tmp_120) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid address\n    at lsu.scala:859 assert(!(will_fire_sta_incoming(w) && stq_incoming_e(w).bits.addr.valid),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_stq_bits_data_bits_T_2 & ~reset & casez_tmp_382) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] Incoming store is overwriting a valid data entry\n    at lsu.scala:878 assert(!(stq(sidx).bits.data.valid),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1430 & ~reset & ~_GEN_1574) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1291 assert(hella_state === h_wait || hella_state === h_dead)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1434 & ~casez_tmp_459) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1295 assert(ldq(io.dmem.nack(w).bits.uop.ldq_idx).bits.executed)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1433 & ~io_dmem_nack_0_bits_uop_uses_ldq & ~reset & ~io_dmem_nack_0_bits_uop_uses_stq) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1301 assert(io.dmem.nack(w).bits.uop.uses_stq)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1575 & io_dmem_resp_0_bits_is_hella) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1312 assert(!io.dmem.resp(w).bits.is_hella)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1575 & (send_iresp ^ ~send_fresp)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1324 assert(send_iresp ^ send_fresp)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & ~reset & io_dmem_resp_0_bits_is_hella) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1332 assert(!io.dmem.resp(w).bits.is_hella)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1471 & ~reset & ~_GEN_1574) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1291 assert(hella_state === h_wait || hella_state === h_dead)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1473 & ~casez_tmp_493) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1295 assert(ldq(io.dmem.nack(w).bits.uop.ldq_idx).bits.executed)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1472 & ~io_dmem_nack_1_bits_uop_uses_ldq & ~reset & ~io_dmem_nack_1_bits_uop_uses_stq) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1301 assert(io.dmem.nack(w).bits.uop.uses_stq)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1576 & io_dmem_resp_1_bits_is_hella) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1312 assert(!io.dmem.resp(w).bits.is_hella)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1576 & (send_iresp_1 ^ ~send_fresp_1)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1324 assert(send_iresp ^ send_fresp)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & ~reset & io_dmem_resp_1_bits_is_hella) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at lsu.scala:1332 assert(!io.dmem.resp(w).bits.is_hella)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1511) & stq_0_valid & stq_0_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1512) & stq_1_valid & stq_1_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1513) & stq_2_valid & stq_2_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1514) & stq_3_valid & stq_3_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1515) & stq_4_valid & stq_4_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1516) & stq_5_valid & stq_5_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1517) & stq_6_valid & stq_6_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1518) & stq_7_valid & stq_7_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1519) & stq_8_valid & stq_8_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1520) & stq_9_valid & stq_9_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1521) & stq_10_valid & stq_10_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1522) & stq_11_valid & stq_11_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1523) & stq_12_valid & stq_12_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1524) & stq_13_valid & stq_13_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1525) & stq_14_valid & stq_14_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1526) & stq_15_valid & stq_15_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1527) & stq_16_valid & stq_16_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1528) & stq_17_valid & stq_17_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1529) & stq_18_valid & stq_18_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1530) & stq_19_valid & stq_19_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1531) & stq_20_valid & stq_20_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1532) & stq_21_valid & stq_21_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1533) & stq_22_valid & stq_22_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1534) & stq_23_valid & stq_23_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1535) & stq_24_valid & stq_24_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1536) & stq_25_valid & stq_25_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1537) & stq_26_valid & stq_26_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1538) & stq_27_valid & stq_27_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1539) & stq_28_valid & stq_28_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1540) & stq_29_valid & stq_29_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1541) & stq_30_valid & stq_30_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|_GEN_1542) & stq_31_valid & stq_31_bits_committed) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1543 & ~casez_tmp_527) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1543 & ~((casez_tmp_528 | casez_tmp_530) & casez_tmp_529)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1548 & ~casez_tmp_531) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1548 & ~((casez_tmp_532 | casez_tmp_534) & casez_tmp_533)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1553 & ~casez_tmp_535) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1553 & ~((casez_tmp_536 | casez_tmp_538) & casez_tmp_537)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1558 & ~casez_tmp_539) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_1558 & ~((casez_tmp_540 | casez_tmp_542) & casez_tmp_541)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
        if (`STOP_COND_)
          $fatal;
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  reg         casez_tmp_543;
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_543 = stq_0_valid;
      5'b00001:
        casez_tmp_543 = stq_1_valid;
      5'b00010:
        casez_tmp_543 = stq_2_valid;
      5'b00011:
        casez_tmp_543 = stq_3_valid;
      5'b00100:
        casez_tmp_543 = stq_4_valid;
      5'b00101:
        casez_tmp_543 = stq_5_valid;
      5'b00110:
        casez_tmp_543 = stq_6_valid;
      5'b00111:
        casez_tmp_543 = stq_7_valid;
      5'b01000:
        casez_tmp_543 = stq_8_valid;
      5'b01001:
        casez_tmp_543 = stq_9_valid;
      5'b01010:
        casez_tmp_543 = stq_10_valid;
      5'b01011:
        casez_tmp_543 = stq_11_valid;
      5'b01100:
        casez_tmp_543 = stq_12_valid;
      5'b01101:
        casez_tmp_543 = stq_13_valid;
      5'b01110:
        casez_tmp_543 = stq_14_valid;
      5'b01111:
        casez_tmp_543 = stq_15_valid;
      5'b10000:
        casez_tmp_543 = stq_16_valid;
      5'b10001:
        casez_tmp_543 = stq_17_valid;
      5'b10010:
        casez_tmp_543 = stq_18_valid;
      5'b10011:
        casez_tmp_543 = stq_19_valid;
      5'b10100:
        casez_tmp_543 = stq_20_valid;
      5'b10101:
        casez_tmp_543 = stq_21_valid;
      5'b10110:
        casez_tmp_543 = stq_22_valid;
      5'b10111:
        casez_tmp_543 = stq_23_valid;
      5'b11000:
        casez_tmp_543 = stq_24_valid;
      5'b11001:
        casez_tmp_543 = stq_25_valid;
      5'b11010:
        casez_tmp_543 = stq_26_valid;
      5'b11011:
        casez_tmp_543 = stq_27_valid;
      5'b11100:
        casez_tmp_543 = stq_28_valid;
      5'b11101:
        casez_tmp_543 = stq_29_valid;
      5'b11110:
        casez_tmp_543 = stq_30_valid;
      default:
        casez_tmp_543 = stq_31_valid;
    endcase
  end // always @(*)
  reg         casez_tmp_544;
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_544 = stq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_544 = stq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_544 = stq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_544 = stq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_544 = stq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_544 = stq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_544 = stq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_544 = stq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_544 = stq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_544 = stq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_544 = stq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_544 = stq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_544 = stq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_544 = stq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_544 = stq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_544 = stq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_544 = stq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_544 = stq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_544 = stq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_544 = stq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_544 = stq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_544 = stq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_544 = stq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_544 = stq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_544 = stq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_544 = stq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_544 = stq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_544 = stq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_544 = stq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_544 = stq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_544 = stq_30_bits_uop_is_fence;
      default:
        casez_tmp_544 = stq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  reg         casez_tmp_545;
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_545 = stq_0_bits_committed;
      5'b00001:
        casez_tmp_545 = stq_1_bits_committed;
      5'b00010:
        casez_tmp_545 = stq_2_bits_committed;
      5'b00011:
        casez_tmp_545 = stq_3_bits_committed;
      5'b00100:
        casez_tmp_545 = stq_4_bits_committed;
      5'b00101:
        casez_tmp_545 = stq_5_bits_committed;
      5'b00110:
        casez_tmp_545 = stq_6_bits_committed;
      5'b00111:
        casez_tmp_545 = stq_7_bits_committed;
      5'b01000:
        casez_tmp_545 = stq_8_bits_committed;
      5'b01001:
        casez_tmp_545 = stq_9_bits_committed;
      5'b01010:
        casez_tmp_545 = stq_10_bits_committed;
      5'b01011:
        casez_tmp_545 = stq_11_bits_committed;
      5'b01100:
        casez_tmp_545 = stq_12_bits_committed;
      5'b01101:
        casez_tmp_545 = stq_13_bits_committed;
      5'b01110:
        casez_tmp_545 = stq_14_bits_committed;
      5'b01111:
        casez_tmp_545 = stq_15_bits_committed;
      5'b10000:
        casez_tmp_545 = stq_16_bits_committed;
      5'b10001:
        casez_tmp_545 = stq_17_bits_committed;
      5'b10010:
        casez_tmp_545 = stq_18_bits_committed;
      5'b10011:
        casez_tmp_545 = stq_19_bits_committed;
      5'b10100:
        casez_tmp_545 = stq_20_bits_committed;
      5'b10101:
        casez_tmp_545 = stq_21_bits_committed;
      5'b10110:
        casez_tmp_545 = stq_22_bits_committed;
      5'b10111:
        casez_tmp_545 = stq_23_bits_committed;
      5'b11000:
        casez_tmp_545 = stq_24_bits_committed;
      5'b11001:
        casez_tmp_545 = stq_25_bits_committed;
      5'b11010:
        casez_tmp_545 = stq_26_bits_committed;
      5'b11011:
        casez_tmp_545 = stq_27_bits_committed;
      5'b11100:
        casez_tmp_545 = stq_28_bits_committed;
      5'b11101:
        casez_tmp_545 = stq_29_bits_committed;
      5'b11110:
        casez_tmp_545 = stq_30_bits_committed;
      default:
        casez_tmp_545 = stq_31_bits_committed;
    endcase
  end // always @(*)
  reg         casez_tmp_546;
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_546 = stq_0_bits_succeeded;
      5'b00001:
        casez_tmp_546 = stq_1_bits_succeeded;
      5'b00010:
        casez_tmp_546 = stq_2_bits_succeeded;
      5'b00011:
        casez_tmp_546 = stq_3_bits_succeeded;
      5'b00100:
        casez_tmp_546 = stq_4_bits_succeeded;
      5'b00101:
        casez_tmp_546 = stq_5_bits_succeeded;
      5'b00110:
        casez_tmp_546 = stq_6_bits_succeeded;
      5'b00111:
        casez_tmp_546 = stq_7_bits_succeeded;
      5'b01000:
        casez_tmp_546 = stq_8_bits_succeeded;
      5'b01001:
        casez_tmp_546 = stq_9_bits_succeeded;
      5'b01010:
        casez_tmp_546 = stq_10_bits_succeeded;
      5'b01011:
        casez_tmp_546 = stq_11_bits_succeeded;
      5'b01100:
        casez_tmp_546 = stq_12_bits_succeeded;
      5'b01101:
        casez_tmp_546 = stq_13_bits_succeeded;
      5'b01110:
        casez_tmp_546 = stq_14_bits_succeeded;
      5'b01111:
        casez_tmp_546 = stq_15_bits_succeeded;
      5'b10000:
        casez_tmp_546 = stq_16_bits_succeeded;
      5'b10001:
        casez_tmp_546 = stq_17_bits_succeeded;
      5'b10010:
        casez_tmp_546 = stq_18_bits_succeeded;
      5'b10011:
        casez_tmp_546 = stq_19_bits_succeeded;
      5'b10100:
        casez_tmp_546 = stq_20_bits_succeeded;
      5'b10101:
        casez_tmp_546 = stq_21_bits_succeeded;
      5'b10110:
        casez_tmp_546 = stq_22_bits_succeeded;
      5'b10111:
        casez_tmp_546 = stq_23_bits_succeeded;
      5'b11000:
        casez_tmp_546 = stq_24_bits_succeeded;
      5'b11001:
        casez_tmp_546 = stq_25_bits_succeeded;
      5'b11010:
        casez_tmp_546 = stq_26_bits_succeeded;
      5'b11011:
        casez_tmp_546 = stq_27_bits_succeeded;
      5'b11100:
        casez_tmp_546 = stq_28_bits_succeeded;
      5'b11101:
        casez_tmp_546 = stq_29_bits_succeeded;
      5'b11110:
        casez_tmp_546 = stq_30_bits_succeeded;
      default:
        casez_tmp_546 = stq_31_bits_succeeded;
    endcase
  end // always @(*)
  wire        _GEN_1577 = casez_tmp_543 & casez_tmp_545;
  wire        _GEN_1578 = casez_tmp_544 & ~io_dmem_ordered;
  assign store_needs_order = _GEN_1577 & _GEN_1578;
  wire        clear_store = _GEN_1577 & (casez_tmp_544 ? io_dmem_ordered : casez_tmp_546);
  wire        _io_hellacache_req_ready_output = hella_state == 3'h0;
  wire        _GEN_1579 = _io_hellacache_req_ready_output & io_hellacache_req_valid;
  assign _GEN_0 = ~_io_hellacache_req_ready_output;
  wire        _GEN_1580 = hella_state == 3'h3;
  wire        _GEN_1581 = _io_hellacache_req_ready_output | _GEN_2;
  wire        _GEN_1582 = hella_state == 3'h2;
  wire        _GEN_1583 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_is_hella;
  wire        _GEN_1584 = io_dmem_resp_1_valid & io_dmem_resp_1_bits_is_hella;
  assign _GEN = ~(_io_hellacache_req_ready_output | _GEN_2 | _GEN_1580 | _GEN_1582 | _GEN_1431);
  reg  [2:0]  casez_tmp_547;
  wire        _GEN_1585 = will_fire_hella_incoming_1_will_fire & dmem_req_fire_1;
  wire [2:0]  _GEN_1586 = _GEN_1432 & (_GEN_1584 | _GEN_1583) ? 3'h0 : hella_state;
  always @(*) begin
    casez (hella_state)
      3'b000:
        casez_tmp_547 = _GEN_1579 ? 3'h1 : hella_state;
      3'b001:
        casez_tmp_547 = io_hellacache_s1_kill ? (_GEN_1585 ? 3'h6 : 3'h0) : {2'h1, ~_GEN_1585};
      3'b010:
        casez_tmp_547 = {1'h1, |{hella_xcpt_ma_ld, hella_xcpt_ma_st, hella_xcpt_pf_ld, hella_xcpt_pf_st, hella_xcpt_gf_ld, hella_xcpt_gf_st, hella_xcpt_ae_ld, hella_xcpt_ae_st}, 1'h0};
      3'b011:
        casez_tmp_547 = 3'h0;
      3'b100:
        casez_tmp_547 = _GEN_1584 ? 3'h0 : _GEN_1471 ? 3'h5 : _GEN_1583 ? 3'h0 : _GEN_1430 ? 3'h5 : hella_state;
      3'b101:
        casez_tmp_547 = will_fire_hella_wakeup_1_will_fire & dmem_req_fire_1 ? 3'h4 : hella_state;
      3'b110:
        casez_tmp_547 = _GEN_1586;
      default:
        casez_tmp_547 = _GEN_1586;
    endcase
  end // always @(*)
  wire        _GEN_1587 = stq_execute_head < stq_head;
  wire [31:0] _ldq_31_bits_st_dep_mask_T = 32'h1 << stq_head;
  wire [31:0] _GEN_1588 = {32{~clear_store}};
  wire [31:0] next_live_store_mask = (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & live_store_mask;
  wire        _GEN_1589 = dis_ld_val & ldq_tail == 5'h0;
  wire        _GEN_1590 = dis_ld_val & ldq_tail == 5'h1;
  wire        _GEN_1591 = dis_ld_val & ldq_tail == 5'h2;
  wire        _GEN_1592 = dis_ld_val & ldq_tail == 5'h3;
  wire        _GEN_1593 = dis_ld_val & ldq_tail == 5'h4;
  wire        _GEN_1594 = dis_ld_val & ldq_tail == 5'h5;
  wire        _GEN_1595 = dis_ld_val & ldq_tail == 5'h6;
  wire        _GEN_1596 = dis_ld_val & ldq_tail == 5'h7;
  wire        _GEN_1597 = dis_ld_val & ldq_tail == 5'h8;
  wire        _GEN_1598 = dis_ld_val & ldq_tail == 5'h9;
  wire        _GEN_1599 = dis_ld_val & ldq_tail == 5'hA;
  wire        _GEN_1600 = dis_ld_val & ldq_tail == 5'hB;
  wire        _GEN_1601 = dis_ld_val & ldq_tail == 5'hC;
  wire        _GEN_1602 = dis_ld_val & ldq_tail == 5'hD;
  wire        _GEN_1603 = dis_ld_val & ldq_tail == 5'hE;
  wire        _GEN_1604 = dis_ld_val & ldq_tail == 5'hF;
  wire        _GEN_1605 = dis_ld_val & ldq_tail == 5'h10;
  wire        _GEN_1606 = dis_ld_val & ldq_tail == 5'h11;
  wire        _GEN_1607 = dis_ld_val & ldq_tail == 5'h12;
  wire        _GEN_1608 = dis_ld_val & ldq_tail == 5'h13;
  wire        _GEN_1609 = dis_ld_val & ldq_tail == 5'h14;
  wire        _GEN_1610 = dis_ld_val & ldq_tail == 5'h15;
  wire        _GEN_1611 = dis_ld_val & ldq_tail == 5'h16;
  wire        _GEN_1612 = dis_ld_val & ldq_tail == 5'h17;
  wire        _GEN_1613 = dis_ld_val & ldq_tail == 5'h18;
  wire        _GEN_1614 = dis_ld_val & ldq_tail == 5'h19;
  wire        _GEN_1615 = dis_ld_val & ldq_tail == 5'h1A;
  wire        _GEN_1616 = dis_ld_val & ldq_tail == 5'h1B;
  wire        _GEN_1617 = dis_ld_val & ldq_tail == 5'h1C;
  wire        _GEN_1618 = dis_ld_val & ldq_tail == 5'h1D;
  wire        _GEN_1619 = dis_ld_val & ldq_tail == 5'h1E;
  wire        _GEN_1620 = dis_ld_val & (&ldq_tail);
  wire        _GEN_1621 = dis_st_val & stq_tail == 5'h0;
  wire        _GEN_1622 = dis_st_val & stq_tail == 5'h1;
  wire        _GEN_1623 = dis_st_val & stq_tail == 5'h2;
  wire        _GEN_1624 = dis_st_val & stq_tail == 5'h3;
  wire        _GEN_1625 = dis_st_val & stq_tail == 5'h4;
  wire        _GEN_1626 = dis_st_val & stq_tail == 5'h5;
  wire        _GEN_1627 = dis_st_val & stq_tail == 5'h6;
  wire        _GEN_1628 = dis_st_val & stq_tail == 5'h7;
  wire        _GEN_1629 = dis_st_val & stq_tail == 5'h8;
  wire        _GEN_1630 = dis_st_val & stq_tail == 5'h9;
  wire        _GEN_1631 = dis_st_val & stq_tail == 5'hA;
  wire        _GEN_1632 = dis_st_val & stq_tail == 5'hB;
  wire        _GEN_1633 = dis_st_val & stq_tail == 5'hC;
  wire        _GEN_1634 = dis_st_val & stq_tail == 5'hD;
  wire        _GEN_1635 = dis_st_val & stq_tail == 5'hE;
  wire        _GEN_1636 = dis_st_val & stq_tail == 5'hF;
  wire        _GEN_1637 = dis_st_val & stq_tail == 5'h10;
  wire        _GEN_1638 = dis_st_val & stq_tail == 5'h11;
  wire        _GEN_1639 = dis_st_val & stq_tail == 5'h12;
  wire        _GEN_1640 = dis_st_val & stq_tail == 5'h13;
  wire        _GEN_1641 = dis_st_val & stq_tail == 5'h14;
  wire        _GEN_1642 = dis_st_val & stq_tail == 5'h15;
  wire        _GEN_1643 = dis_st_val & stq_tail == 5'h16;
  wire        _GEN_1644 = dis_st_val & stq_tail == 5'h17;
  wire        _GEN_1645 = dis_st_val & stq_tail == 5'h18;
  wire        _GEN_1646 = dis_st_val & stq_tail == 5'h19;
  wire        _GEN_1647 = dis_st_val & stq_tail == 5'h1A;
  wire        _GEN_1648 = dis_st_val & stq_tail == 5'h1B;
  wire        _GEN_1649 = dis_st_val & stq_tail == 5'h1C;
  wire        _GEN_1650 = dis_st_val & stq_tail == 5'h1D;
  wire        _GEN_1651 = dis_st_val & stq_tail == 5'h1E;
  wire        _GEN_1652 = dis_st_val & (&stq_tail);
  wire        _GEN_1653 = dis_ld_val | ~_GEN_1621;
  wire        _GEN_1654 = dis_ld_val | ~_GEN_1622;
  wire        _GEN_1655 = dis_ld_val | ~_GEN_1623;
  wire        _GEN_1656 = dis_ld_val | ~_GEN_1624;
  wire        _GEN_1657 = dis_ld_val | ~_GEN_1625;
  wire        _GEN_1658 = dis_ld_val | ~_GEN_1626;
  wire        _GEN_1659 = dis_ld_val | ~_GEN_1627;
  wire        _GEN_1660 = dis_ld_val | ~_GEN_1628;
  wire        _GEN_1661 = dis_ld_val | ~_GEN_1629;
  wire        _GEN_1662 = dis_ld_val | ~_GEN_1630;
  wire        _GEN_1663 = dis_ld_val | ~_GEN_1631;
  wire        _GEN_1664 = dis_ld_val | ~_GEN_1632;
  wire        _GEN_1665 = dis_ld_val | ~_GEN_1633;
  wire        _GEN_1666 = dis_ld_val | ~_GEN_1634;
  wire        _GEN_1667 = dis_ld_val | ~_GEN_1635;
  wire        _GEN_1668 = dis_ld_val | ~_GEN_1636;
  wire        _GEN_1669 = dis_ld_val | ~_GEN_1637;
  wire        _GEN_1670 = dis_ld_val | ~_GEN_1638;
  wire        _GEN_1671 = dis_ld_val | ~_GEN_1639;
  wire        _GEN_1672 = dis_ld_val | ~_GEN_1640;
  wire        _GEN_1673 = dis_ld_val | ~_GEN_1641;
  wire        _GEN_1674 = dis_ld_val | ~_GEN_1642;
  wire        _GEN_1675 = dis_ld_val | ~_GEN_1643;
  wire        _GEN_1676 = dis_ld_val | ~_GEN_1644;
  wire        _GEN_1677 = dis_ld_val | ~_GEN_1645;
  wire        _GEN_1678 = dis_ld_val | ~_GEN_1646;
  wire        _GEN_1679 = dis_ld_val | ~_GEN_1647;
  wire        _GEN_1680 = dis_ld_val | ~_GEN_1648;
  wire        _GEN_1681 = dis_ld_val | ~_GEN_1649;
  wire        _GEN_1682 = dis_ld_val | ~_GEN_1650;
  wire        _GEN_1683 = dis_ld_val | ~_GEN_1651;
  wire        _GEN_1684 = dis_ld_val | ~_GEN_1652;
  wire [31:0] _GEN_1685 = {32{dis_st_val}} & 32'h1 << stq_tail | next_live_store_mask;
  wire        _GEN_1686 = _GEN_5 == 5'h0;
  wire        _GEN_1687 = _GEN_1686 | _GEN_1589;
  wire        _GEN_1688 = dis_ld_val_1 ? _GEN_1687 | ldq_0_valid : _GEN_1589 | ldq_0_valid;
  wire        _GEN_1689 = _GEN_5 == 5'h1;
  wire        _GEN_1690 = _GEN_1689 | _GEN_1590;
  wire        _GEN_1691 = dis_ld_val_1 ? _GEN_1690 | ldq_1_valid : _GEN_1590 | ldq_1_valid;
  wire        _GEN_1692 = _GEN_5 == 5'h2;
  wire        _GEN_1693 = _GEN_1692 | _GEN_1591;
  wire        _GEN_1694 = dis_ld_val_1 ? _GEN_1693 | ldq_2_valid : _GEN_1591 | ldq_2_valid;
  wire        _GEN_1695 = _GEN_5 == 5'h3;
  wire        _GEN_1696 = _GEN_1695 | _GEN_1592;
  wire        _GEN_1697 = dis_ld_val_1 ? _GEN_1696 | ldq_3_valid : _GEN_1592 | ldq_3_valid;
  wire        _GEN_1698 = _GEN_5 == 5'h4;
  wire        _GEN_1699 = _GEN_1698 | _GEN_1593;
  wire        _GEN_1700 = dis_ld_val_1 ? _GEN_1699 | ldq_4_valid : _GEN_1593 | ldq_4_valid;
  wire        _GEN_1701 = _GEN_5 == 5'h5;
  wire        _GEN_1702 = _GEN_1701 | _GEN_1594;
  wire        _GEN_1703 = dis_ld_val_1 ? _GEN_1702 | ldq_5_valid : _GEN_1594 | ldq_5_valid;
  wire        _GEN_1704 = _GEN_5 == 5'h6;
  wire        _GEN_1705 = _GEN_1704 | _GEN_1595;
  wire        _GEN_1706 = dis_ld_val_1 ? _GEN_1705 | ldq_6_valid : _GEN_1595 | ldq_6_valid;
  wire        _GEN_1707 = _GEN_5 == 5'h7;
  wire        _GEN_1708 = _GEN_1707 | _GEN_1596;
  wire        _GEN_1709 = dis_ld_val_1 ? _GEN_1708 | ldq_7_valid : _GEN_1596 | ldq_7_valid;
  wire        _GEN_1710 = _GEN_5 == 5'h8;
  wire        _GEN_1711 = _GEN_1710 | _GEN_1597;
  wire        _GEN_1712 = dis_ld_val_1 ? _GEN_1711 | ldq_8_valid : _GEN_1597 | ldq_8_valid;
  wire        _GEN_1713 = _GEN_5 == 5'h9;
  wire        _GEN_1714 = _GEN_1713 | _GEN_1598;
  wire        _GEN_1715 = dis_ld_val_1 ? _GEN_1714 | ldq_9_valid : _GEN_1598 | ldq_9_valid;
  wire        _GEN_1716 = _GEN_5 == 5'hA;
  wire        _GEN_1717 = _GEN_1716 | _GEN_1599;
  wire        _GEN_1718 = dis_ld_val_1 ? _GEN_1717 | ldq_10_valid : _GEN_1599 | ldq_10_valid;
  wire        _GEN_1719 = _GEN_5 == 5'hB;
  wire        _GEN_1720 = _GEN_1719 | _GEN_1600;
  wire        _GEN_1721 = dis_ld_val_1 ? _GEN_1720 | ldq_11_valid : _GEN_1600 | ldq_11_valid;
  wire        _GEN_1722 = _GEN_5 == 5'hC;
  wire        _GEN_1723 = _GEN_1722 | _GEN_1601;
  wire        _GEN_1724 = dis_ld_val_1 ? _GEN_1723 | ldq_12_valid : _GEN_1601 | ldq_12_valid;
  wire        _GEN_1725 = _GEN_5 == 5'hD;
  wire        _GEN_1726 = _GEN_1725 | _GEN_1602;
  wire        _GEN_1727 = dis_ld_val_1 ? _GEN_1726 | ldq_13_valid : _GEN_1602 | ldq_13_valid;
  wire        _GEN_1728 = _GEN_5 == 5'hE;
  wire        _GEN_1729 = _GEN_1728 | _GEN_1603;
  wire        _GEN_1730 = dis_ld_val_1 ? _GEN_1729 | ldq_14_valid : _GEN_1603 | ldq_14_valid;
  wire        _GEN_1731 = _GEN_5 == 5'hF;
  wire        _GEN_1732 = _GEN_1731 | _GEN_1604;
  wire        _GEN_1733 = dis_ld_val_1 ? _GEN_1732 | ldq_15_valid : _GEN_1604 | ldq_15_valid;
  wire        _GEN_1734 = _GEN_5 == 5'h10;
  wire        _GEN_1735 = _GEN_1734 | _GEN_1605;
  wire        _GEN_1736 = dis_ld_val_1 ? _GEN_1735 | ldq_16_valid : _GEN_1605 | ldq_16_valid;
  wire        _GEN_1737 = _GEN_5 == 5'h11;
  wire        _GEN_1738 = _GEN_1737 | _GEN_1606;
  wire        _GEN_1739 = dis_ld_val_1 ? _GEN_1738 | ldq_17_valid : _GEN_1606 | ldq_17_valid;
  wire        _GEN_1740 = _GEN_5 == 5'h12;
  wire        _GEN_1741 = _GEN_1740 | _GEN_1607;
  wire        _GEN_1742 = dis_ld_val_1 ? _GEN_1741 | ldq_18_valid : _GEN_1607 | ldq_18_valid;
  wire        _GEN_1743 = _GEN_5 == 5'h13;
  wire        _GEN_1744 = _GEN_1743 | _GEN_1608;
  wire        _GEN_1745 = dis_ld_val_1 ? _GEN_1744 | ldq_19_valid : _GEN_1608 | ldq_19_valid;
  wire        _GEN_1746 = _GEN_5 == 5'h14;
  wire        _GEN_1747 = _GEN_1746 | _GEN_1609;
  wire        _GEN_1748 = dis_ld_val_1 ? _GEN_1747 | ldq_20_valid : _GEN_1609 | ldq_20_valid;
  wire        _GEN_1749 = _GEN_5 == 5'h15;
  wire        _GEN_1750 = _GEN_1749 | _GEN_1610;
  wire        _GEN_1751 = dis_ld_val_1 ? _GEN_1750 | ldq_21_valid : _GEN_1610 | ldq_21_valid;
  wire        _GEN_1752 = _GEN_5 == 5'h16;
  wire        _GEN_1753 = _GEN_1752 | _GEN_1611;
  wire        _GEN_1754 = dis_ld_val_1 ? _GEN_1753 | ldq_22_valid : _GEN_1611 | ldq_22_valid;
  wire        _GEN_1755 = _GEN_5 == 5'h17;
  wire        _GEN_1756 = _GEN_1755 | _GEN_1612;
  wire        _GEN_1757 = dis_ld_val_1 ? _GEN_1756 | ldq_23_valid : _GEN_1612 | ldq_23_valid;
  wire        _GEN_1758 = _GEN_5 == 5'h18;
  wire        _GEN_1759 = _GEN_1758 | _GEN_1613;
  wire        _GEN_1760 = dis_ld_val_1 ? _GEN_1759 | ldq_24_valid : _GEN_1613 | ldq_24_valid;
  wire        _GEN_1761 = _GEN_5 == 5'h19;
  wire        _GEN_1762 = _GEN_1761 | _GEN_1614;
  wire        _GEN_1763 = dis_ld_val_1 ? _GEN_1762 | ldq_25_valid : _GEN_1614 | ldq_25_valid;
  wire        _GEN_1764 = _GEN_5 == 5'h1A;
  wire        _GEN_1765 = _GEN_1764 | _GEN_1615;
  wire        _GEN_1766 = dis_ld_val_1 ? _GEN_1765 | ldq_26_valid : _GEN_1615 | ldq_26_valid;
  wire        _GEN_1767 = _GEN_5 == 5'h1B;
  wire        _GEN_1768 = _GEN_1767 | _GEN_1616;
  wire        _GEN_1769 = dis_ld_val_1 ? _GEN_1768 | ldq_27_valid : _GEN_1616 | ldq_27_valid;
  wire        _GEN_1770 = _GEN_5 == 5'h1C;
  wire        _GEN_1771 = _GEN_1770 | _GEN_1617;
  wire        _GEN_1772 = dis_ld_val_1 ? _GEN_1771 | ldq_28_valid : _GEN_1617 | ldq_28_valid;
  wire        _GEN_1773 = _GEN_5 == 5'h1D;
  wire        _GEN_1774 = _GEN_1773 | _GEN_1618;
  wire        _GEN_1775 = dis_ld_val_1 ? _GEN_1774 | ldq_29_valid : _GEN_1618 | ldq_29_valid;
  wire        _GEN_1776 = _GEN_5 == 5'h1E;
  wire        _GEN_1777 = _GEN_1776 | _GEN_1619;
  wire        _GEN_1778 = dis_ld_val_1 ? _GEN_1777 | ldq_30_valid : _GEN_1619 | ldq_30_valid;
  wire        _GEN_1779 = (&_GEN_5) | _GEN_1620;
  wire        _GEN_1780 = dis_ld_val_1 ? _GEN_1779 | ldq_31_valid : _GEN_1620 | ldq_31_valid;
  wire        _GEN_1781 = dis_ld_val_1 & _GEN_1686;
  wire        _GEN_1782 = dis_ld_val_1 & _GEN_1689;
  wire        _GEN_1783 = dis_ld_val_1 & _GEN_1692;
  wire        _GEN_1784 = dis_ld_val_1 & _GEN_1695;
  wire        _GEN_1785 = dis_ld_val_1 & _GEN_1698;
  wire        _GEN_1786 = dis_ld_val_1 & _GEN_1701;
  wire        _GEN_1787 = dis_ld_val_1 & _GEN_1704;
  wire        _GEN_1788 = dis_ld_val_1 & _GEN_1707;
  wire        _GEN_1789 = dis_ld_val_1 & _GEN_1710;
  wire        _GEN_1790 = dis_ld_val_1 & _GEN_1713;
  wire        _GEN_1791 = dis_ld_val_1 & _GEN_1716;
  wire        _GEN_1792 = dis_ld_val_1 & _GEN_1719;
  wire        _GEN_1793 = dis_ld_val_1 & _GEN_1722;
  wire        _GEN_1794 = dis_ld_val_1 & _GEN_1725;
  wire        _GEN_1795 = dis_ld_val_1 & _GEN_1728;
  wire        _GEN_1796 = dis_ld_val_1 & _GEN_1731;
  wire        _GEN_1797 = dis_ld_val_1 & _GEN_1734;
  wire        _GEN_1798 = dis_ld_val_1 & _GEN_1737;
  wire        _GEN_1799 = dis_ld_val_1 & _GEN_1740;
  wire        _GEN_1800 = dis_ld_val_1 & _GEN_1743;
  wire        _GEN_1801 = dis_ld_val_1 & _GEN_1746;
  wire        _GEN_1802 = dis_ld_val_1 & _GEN_1749;
  wire        _GEN_1803 = dis_ld_val_1 & _GEN_1752;
  wire        _GEN_1804 = dis_ld_val_1 & _GEN_1755;
  wire        _GEN_1805 = dis_ld_val_1 & _GEN_1758;
  wire        _GEN_1806 = dis_ld_val_1 & _GEN_1761;
  wire        _GEN_1807 = dis_ld_val_1 & _GEN_1764;
  wire        _GEN_1808 = dis_ld_val_1 & _GEN_1767;
  wire        _GEN_1809 = dis_ld_val_1 & _GEN_1770;
  wire        _GEN_1810 = dis_ld_val_1 & _GEN_1773;
  wire        _GEN_1811 = dis_ld_val_1 & _GEN_1776;
  wire        _GEN_1812 = dis_ld_val_1 & (&_GEN_5);
  wire        _GEN_1813 = dis_ld_val_1 ? ~_GEN_1687 & ldq_0_bits_addr_valid : ~_GEN_1589 & ldq_0_bits_addr_valid;
  wire        _GEN_1814 = dis_ld_val_1 ? ~_GEN_1690 & ldq_1_bits_addr_valid : ~_GEN_1590 & ldq_1_bits_addr_valid;
  wire        _GEN_1815 = dis_ld_val_1 ? ~_GEN_1693 & ldq_2_bits_addr_valid : ~_GEN_1591 & ldq_2_bits_addr_valid;
  wire        _GEN_1816 = dis_ld_val_1 ? ~_GEN_1696 & ldq_3_bits_addr_valid : ~_GEN_1592 & ldq_3_bits_addr_valid;
  wire        _GEN_1817 = dis_ld_val_1 ? ~_GEN_1699 & ldq_4_bits_addr_valid : ~_GEN_1593 & ldq_4_bits_addr_valid;
  wire        _GEN_1818 = dis_ld_val_1 ? ~_GEN_1702 & ldq_5_bits_addr_valid : ~_GEN_1594 & ldq_5_bits_addr_valid;
  wire        _GEN_1819 = dis_ld_val_1 ? ~_GEN_1705 & ldq_6_bits_addr_valid : ~_GEN_1595 & ldq_6_bits_addr_valid;
  wire        _GEN_1820 = dis_ld_val_1 ? ~_GEN_1708 & ldq_7_bits_addr_valid : ~_GEN_1596 & ldq_7_bits_addr_valid;
  wire        _GEN_1821 = dis_ld_val_1 ? ~_GEN_1711 & ldq_8_bits_addr_valid : ~_GEN_1597 & ldq_8_bits_addr_valid;
  wire        _GEN_1822 = dis_ld_val_1 ? ~_GEN_1714 & ldq_9_bits_addr_valid : ~_GEN_1598 & ldq_9_bits_addr_valid;
  wire        _GEN_1823 = dis_ld_val_1 ? ~_GEN_1717 & ldq_10_bits_addr_valid : ~_GEN_1599 & ldq_10_bits_addr_valid;
  wire        _GEN_1824 = dis_ld_val_1 ? ~_GEN_1720 & ldq_11_bits_addr_valid : ~_GEN_1600 & ldq_11_bits_addr_valid;
  wire        _GEN_1825 = dis_ld_val_1 ? ~_GEN_1723 & ldq_12_bits_addr_valid : ~_GEN_1601 & ldq_12_bits_addr_valid;
  wire        _GEN_1826 = dis_ld_val_1 ? ~_GEN_1726 & ldq_13_bits_addr_valid : ~_GEN_1602 & ldq_13_bits_addr_valid;
  wire        _GEN_1827 = dis_ld_val_1 ? ~_GEN_1729 & ldq_14_bits_addr_valid : ~_GEN_1603 & ldq_14_bits_addr_valid;
  wire        _GEN_1828 = dis_ld_val_1 ? ~_GEN_1732 & ldq_15_bits_addr_valid : ~_GEN_1604 & ldq_15_bits_addr_valid;
  wire        _GEN_1829 = dis_ld_val_1 ? ~_GEN_1735 & ldq_16_bits_addr_valid : ~_GEN_1605 & ldq_16_bits_addr_valid;
  wire        _GEN_1830 = dis_ld_val_1 ? ~_GEN_1738 & ldq_17_bits_addr_valid : ~_GEN_1606 & ldq_17_bits_addr_valid;
  wire        _GEN_1831 = dis_ld_val_1 ? ~_GEN_1741 & ldq_18_bits_addr_valid : ~_GEN_1607 & ldq_18_bits_addr_valid;
  wire        _GEN_1832 = dis_ld_val_1 ? ~_GEN_1744 & ldq_19_bits_addr_valid : ~_GEN_1608 & ldq_19_bits_addr_valid;
  wire        _GEN_1833 = dis_ld_val_1 ? ~_GEN_1747 & ldq_20_bits_addr_valid : ~_GEN_1609 & ldq_20_bits_addr_valid;
  wire        _GEN_1834 = dis_ld_val_1 ? ~_GEN_1750 & ldq_21_bits_addr_valid : ~_GEN_1610 & ldq_21_bits_addr_valid;
  wire        _GEN_1835 = dis_ld_val_1 ? ~_GEN_1753 & ldq_22_bits_addr_valid : ~_GEN_1611 & ldq_22_bits_addr_valid;
  wire        _GEN_1836 = dis_ld_val_1 ? ~_GEN_1756 & ldq_23_bits_addr_valid : ~_GEN_1612 & ldq_23_bits_addr_valid;
  wire        _GEN_1837 = dis_ld_val_1 ? ~_GEN_1759 & ldq_24_bits_addr_valid : ~_GEN_1613 & ldq_24_bits_addr_valid;
  wire        _GEN_1838 = dis_ld_val_1 ? ~_GEN_1762 & ldq_25_bits_addr_valid : ~_GEN_1614 & ldq_25_bits_addr_valid;
  wire        _GEN_1839 = dis_ld_val_1 ? ~_GEN_1765 & ldq_26_bits_addr_valid : ~_GEN_1615 & ldq_26_bits_addr_valid;
  wire        _GEN_1840 = dis_ld_val_1 ? ~_GEN_1768 & ldq_27_bits_addr_valid : ~_GEN_1616 & ldq_27_bits_addr_valid;
  wire        _GEN_1841 = dis_ld_val_1 ? ~_GEN_1771 & ldq_28_bits_addr_valid : ~_GEN_1617 & ldq_28_bits_addr_valid;
  wire        _GEN_1842 = dis_ld_val_1 ? ~_GEN_1774 & ldq_29_bits_addr_valid : ~_GEN_1618 & ldq_29_bits_addr_valid;
  wire        _GEN_1843 = dis_ld_val_1 ? ~_GEN_1777 & ldq_30_bits_addr_valid : ~_GEN_1619 & ldq_30_bits_addr_valid;
  wire        _GEN_1844 = dis_ld_val_1 ? ~_GEN_1779 & ldq_31_bits_addr_valid : ~_GEN_1620 & ldq_31_bits_addr_valid;
  wire        _GEN_1845 = dis_ld_val_1 ? ~_GEN_1687 & ldq_0_bits_executed : ~_GEN_1589 & ldq_0_bits_executed;
  wire        _GEN_1846 = dis_ld_val_1 ? ~_GEN_1690 & ldq_1_bits_executed : ~_GEN_1590 & ldq_1_bits_executed;
  wire        _GEN_1847 = dis_ld_val_1 ? ~_GEN_1693 & ldq_2_bits_executed : ~_GEN_1591 & ldq_2_bits_executed;
  wire        _GEN_1848 = dis_ld_val_1 ? ~_GEN_1696 & ldq_3_bits_executed : ~_GEN_1592 & ldq_3_bits_executed;
  wire        _GEN_1849 = dis_ld_val_1 ? ~_GEN_1699 & ldq_4_bits_executed : ~_GEN_1593 & ldq_4_bits_executed;
  wire        _GEN_1850 = dis_ld_val_1 ? ~_GEN_1702 & ldq_5_bits_executed : ~_GEN_1594 & ldq_5_bits_executed;
  wire        _GEN_1851 = dis_ld_val_1 ? ~_GEN_1705 & ldq_6_bits_executed : ~_GEN_1595 & ldq_6_bits_executed;
  wire        _GEN_1852 = dis_ld_val_1 ? ~_GEN_1708 & ldq_7_bits_executed : ~_GEN_1596 & ldq_7_bits_executed;
  wire        _GEN_1853 = dis_ld_val_1 ? ~_GEN_1711 & ldq_8_bits_executed : ~_GEN_1597 & ldq_8_bits_executed;
  wire        _GEN_1854 = dis_ld_val_1 ? ~_GEN_1714 & ldq_9_bits_executed : ~_GEN_1598 & ldq_9_bits_executed;
  wire        _GEN_1855 = dis_ld_val_1 ? ~_GEN_1717 & ldq_10_bits_executed : ~_GEN_1599 & ldq_10_bits_executed;
  wire        _GEN_1856 = dis_ld_val_1 ? ~_GEN_1720 & ldq_11_bits_executed : ~_GEN_1600 & ldq_11_bits_executed;
  wire        _GEN_1857 = dis_ld_val_1 ? ~_GEN_1723 & ldq_12_bits_executed : ~_GEN_1601 & ldq_12_bits_executed;
  wire        _GEN_1858 = dis_ld_val_1 ? ~_GEN_1726 & ldq_13_bits_executed : ~_GEN_1602 & ldq_13_bits_executed;
  wire        _GEN_1859 = dis_ld_val_1 ? ~_GEN_1729 & ldq_14_bits_executed : ~_GEN_1603 & ldq_14_bits_executed;
  wire        _GEN_1860 = dis_ld_val_1 ? ~_GEN_1732 & ldq_15_bits_executed : ~_GEN_1604 & ldq_15_bits_executed;
  wire        _GEN_1861 = dis_ld_val_1 ? ~_GEN_1735 & ldq_16_bits_executed : ~_GEN_1605 & ldq_16_bits_executed;
  wire        _GEN_1862 = dis_ld_val_1 ? ~_GEN_1738 & ldq_17_bits_executed : ~_GEN_1606 & ldq_17_bits_executed;
  wire        _GEN_1863 = dis_ld_val_1 ? ~_GEN_1741 & ldq_18_bits_executed : ~_GEN_1607 & ldq_18_bits_executed;
  wire        _GEN_1864 = dis_ld_val_1 ? ~_GEN_1744 & ldq_19_bits_executed : ~_GEN_1608 & ldq_19_bits_executed;
  wire        _GEN_1865 = dis_ld_val_1 ? ~_GEN_1747 & ldq_20_bits_executed : ~_GEN_1609 & ldq_20_bits_executed;
  wire        _GEN_1866 = dis_ld_val_1 ? ~_GEN_1750 & ldq_21_bits_executed : ~_GEN_1610 & ldq_21_bits_executed;
  wire        _GEN_1867 = dis_ld_val_1 ? ~_GEN_1753 & ldq_22_bits_executed : ~_GEN_1611 & ldq_22_bits_executed;
  wire        _GEN_1868 = dis_ld_val_1 ? ~_GEN_1756 & ldq_23_bits_executed : ~_GEN_1612 & ldq_23_bits_executed;
  wire        _GEN_1869 = dis_ld_val_1 ? ~_GEN_1759 & ldq_24_bits_executed : ~_GEN_1613 & ldq_24_bits_executed;
  wire        _GEN_1870 = dis_ld_val_1 ? ~_GEN_1762 & ldq_25_bits_executed : ~_GEN_1614 & ldq_25_bits_executed;
  wire        _GEN_1871 = dis_ld_val_1 ? ~_GEN_1765 & ldq_26_bits_executed : ~_GEN_1615 & ldq_26_bits_executed;
  wire        _GEN_1872 = dis_ld_val_1 ? ~_GEN_1768 & ldq_27_bits_executed : ~_GEN_1616 & ldq_27_bits_executed;
  wire        _GEN_1873 = dis_ld_val_1 ? ~_GEN_1771 & ldq_28_bits_executed : ~_GEN_1617 & ldq_28_bits_executed;
  wire        _GEN_1874 = dis_ld_val_1 ? ~_GEN_1774 & ldq_29_bits_executed : ~_GEN_1618 & ldq_29_bits_executed;
  wire        _GEN_1875 = dis_ld_val_1 ? ~_GEN_1777 & ldq_30_bits_executed : ~_GEN_1619 & ldq_30_bits_executed;
  wire        _GEN_1876 = dis_ld_val_1 ? ~_GEN_1779 & ldq_31_bits_executed : ~_GEN_1620 & ldq_31_bits_executed;
  wire        _GEN_1877 = dis_ld_val_1 ? ~_GEN_1687 & ldq_0_bits_succeeded : ~_GEN_1589 & ldq_0_bits_succeeded;
  wire        _GEN_1878 = dis_ld_val_1 ? ~_GEN_1690 & ldq_1_bits_succeeded : ~_GEN_1590 & ldq_1_bits_succeeded;
  wire        _GEN_1879 = dis_ld_val_1 ? ~_GEN_1693 & ldq_2_bits_succeeded : ~_GEN_1591 & ldq_2_bits_succeeded;
  wire        _GEN_1880 = dis_ld_val_1 ? ~_GEN_1696 & ldq_3_bits_succeeded : ~_GEN_1592 & ldq_3_bits_succeeded;
  wire        _GEN_1881 = dis_ld_val_1 ? ~_GEN_1699 & ldq_4_bits_succeeded : ~_GEN_1593 & ldq_4_bits_succeeded;
  wire        _GEN_1882 = dis_ld_val_1 ? ~_GEN_1702 & ldq_5_bits_succeeded : ~_GEN_1594 & ldq_5_bits_succeeded;
  wire        _GEN_1883 = dis_ld_val_1 ? ~_GEN_1705 & ldq_6_bits_succeeded : ~_GEN_1595 & ldq_6_bits_succeeded;
  wire        _GEN_1884 = dis_ld_val_1 ? ~_GEN_1708 & ldq_7_bits_succeeded : ~_GEN_1596 & ldq_7_bits_succeeded;
  wire        _GEN_1885 = dis_ld_val_1 ? ~_GEN_1711 & ldq_8_bits_succeeded : ~_GEN_1597 & ldq_8_bits_succeeded;
  wire        _GEN_1886 = dis_ld_val_1 ? ~_GEN_1714 & ldq_9_bits_succeeded : ~_GEN_1598 & ldq_9_bits_succeeded;
  wire        _GEN_1887 = dis_ld_val_1 ? ~_GEN_1717 & ldq_10_bits_succeeded : ~_GEN_1599 & ldq_10_bits_succeeded;
  wire        _GEN_1888 = dis_ld_val_1 ? ~_GEN_1720 & ldq_11_bits_succeeded : ~_GEN_1600 & ldq_11_bits_succeeded;
  wire        _GEN_1889 = dis_ld_val_1 ? ~_GEN_1723 & ldq_12_bits_succeeded : ~_GEN_1601 & ldq_12_bits_succeeded;
  wire        _GEN_1890 = dis_ld_val_1 ? ~_GEN_1726 & ldq_13_bits_succeeded : ~_GEN_1602 & ldq_13_bits_succeeded;
  wire        _GEN_1891 = dis_ld_val_1 ? ~_GEN_1729 & ldq_14_bits_succeeded : ~_GEN_1603 & ldq_14_bits_succeeded;
  wire        _GEN_1892 = dis_ld_val_1 ? ~_GEN_1732 & ldq_15_bits_succeeded : ~_GEN_1604 & ldq_15_bits_succeeded;
  wire        _GEN_1893 = dis_ld_val_1 ? ~_GEN_1735 & ldq_16_bits_succeeded : ~_GEN_1605 & ldq_16_bits_succeeded;
  wire        _GEN_1894 = dis_ld_val_1 ? ~_GEN_1738 & ldq_17_bits_succeeded : ~_GEN_1606 & ldq_17_bits_succeeded;
  wire        _GEN_1895 = dis_ld_val_1 ? ~_GEN_1741 & ldq_18_bits_succeeded : ~_GEN_1607 & ldq_18_bits_succeeded;
  wire        _GEN_1896 = dis_ld_val_1 ? ~_GEN_1744 & ldq_19_bits_succeeded : ~_GEN_1608 & ldq_19_bits_succeeded;
  wire        _GEN_1897 = dis_ld_val_1 ? ~_GEN_1747 & ldq_20_bits_succeeded : ~_GEN_1609 & ldq_20_bits_succeeded;
  wire        _GEN_1898 = dis_ld_val_1 ? ~_GEN_1750 & ldq_21_bits_succeeded : ~_GEN_1610 & ldq_21_bits_succeeded;
  wire        _GEN_1899 = dis_ld_val_1 ? ~_GEN_1753 & ldq_22_bits_succeeded : ~_GEN_1611 & ldq_22_bits_succeeded;
  wire        _GEN_1900 = dis_ld_val_1 ? ~_GEN_1756 & ldq_23_bits_succeeded : ~_GEN_1612 & ldq_23_bits_succeeded;
  wire        _GEN_1901 = dis_ld_val_1 ? ~_GEN_1759 & ldq_24_bits_succeeded : ~_GEN_1613 & ldq_24_bits_succeeded;
  wire        _GEN_1902 = dis_ld_val_1 ? ~_GEN_1762 & ldq_25_bits_succeeded : ~_GEN_1614 & ldq_25_bits_succeeded;
  wire        _GEN_1903 = dis_ld_val_1 ? ~_GEN_1765 & ldq_26_bits_succeeded : ~_GEN_1615 & ldq_26_bits_succeeded;
  wire        _GEN_1904 = dis_ld_val_1 ? ~_GEN_1768 & ldq_27_bits_succeeded : ~_GEN_1616 & ldq_27_bits_succeeded;
  wire        _GEN_1905 = dis_ld_val_1 ? ~_GEN_1771 & ldq_28_bits_succeeded : ~_GEN_1617 & ldq_28_bits_succeeded;
  wire        _GEN_1906 = dis_ld_val_1 ? ~_GEN_1774 & ldq_29_bits_succeeded : ~_GEN_1618 & ldq_29_bits_succeeded;
  wire        _GEN_1907 = dis_ld_val_1 ? ~_GEN_1777 & ldq_30_bits_succeeded : ~_GEN_1619 & ldq_30_bits_succeeded;
  wire        _GEN_1908 = dis_ld_val_1 ? ~_GEN_1779 & ldq_31_bits_succeeded : ~_GEN_1620 & ldq_31_bits_succeeded;
  wire        _GEN_1909 = dis_ld_val_1 ? ~_GEN_1687 & ldq_0_bits_order_fail : ~_GEN_1589 & ldq_0_bits_order_fail;
  wire        _GEN_1910 = dis_ld_val_1 ? ~_GEN_1690 & ldq_1_bits_order_fail : ~_GEN_1590 & ldq_1_bits_order_fail;
  wire        _GEN_1911 = dis_ld_val_1 ? ~_GEN_1693 & ldq_2_bits_order_fail : ~_GEN_1591 & ldq_2_bits_order_fail;
  wire        _GEN_1912 = dis_ld_val_1 ? ~_GEN_1696 & ldq_3_bits_order_fail : ~_GEN_1592 & ldq_3_bits_order_fail;
  wire        _GEN_1913 = dis_ld_val_1 ? ~_GEN_1699 & ldq_4_bits_order_fail : ~_GEN_1593 & ldq_4_bits_order_fail;
  wire        _GEN_1914 = dis_ld_val_1 ? ~_GEN_1702 & ldq_5_bits_order_fail : ~_GEN_1594 & ldq_5_bits_order_fail;
  wire        _GEN_1915 = dis_ld_val_1 ? ~_GEN_1705 & ldq_6_bits_order_fail : ~_GEN_1595 & ldq_6_bits_order_fail;
  wire        _GEN_1916 = dis_ld_val_1 ? ~_GEN_1708 & ldq_7_bits_order_fail : ~_GEN_1596 & ldq_7_bits_order_fail;
  wire        _GEN_1917 = dis_ld_val_1 ? ~_GEN_1711 & ldq_8_bits_order_fail : ~_GEN_1597 & ldq_8_bits_order_fail;
  wire        _GEN_1918 = dis_ld_val_1 ? ~_GEN_1714 & ldq_9_bits_order_fail : ~_GEN_1598 & ldq_9_bits_order_fail;
  wire        _GEN_1919 = dis_ld_val_1 ? ~_GEN_1717 & ldq_10_bits_order_fail : ~_GEN_1599 & ldq_10_bits_order_fail;
  wire        _GEN_1920 = dis_ld_val_1 ? ~_GEN_1720 & ldq_11_bits_order_fail : ~_GEN_1600 & ldq_11_bits_order_fail;
  wire        _GEN_1921 = dis_ld_val_1 ? ~_GEN_1723 & ldq_12_bits_order_fail : ~_GEN_1601 & ldq_12_bits_order_fail;
  wire        _GEN_1922 = dis_ld_val_1 ? ~_GEN_1726 & ldq_13_bits_order_fail : ~_GEN_1602 & ldq_13_bits_order_fail;
  wire        _GEN_1923 = dis_ld_val_1 ? ~_GEN_1729 & ldq_14_bits_order_fail : ~_GEN_1603 & ldq_14_bits_order_fail;
  wire        _GEN_1924 = dis_ld_val_1 ? ~_GEN_1732 & ldq_15_bits_order_fail : ~_GEN_1604 & ldq_15_bits_order_fail;
  wire        _GEN_1925 = dis_ld_val_1 ? ~_GEN_1735 & ldq_16_bits_order_fail : ~_GEN_1605 & ldq_16_bits_order_fail;
  wire        _GEN_1926 = dis_ld_val_1 ? ~_GEN_1738 & ldq_17_bits_order_fail : ~_GEN_1606 & ldq_17_bits_order_fail;
  wire        _GEN_1927 = dis_ld_val_1 ? ~_GEN_1741 & ldq_18_bits_order_fail : ~_GEN_1607 & ldq_18_bits_order_fail;
  wire        _GEN_1928 = dis_ld_val_1 ? ~_GEN_1744 & ldq_19_bits_order_fail : ~_GEN_1608 & ldq_19_bits_order_fail;
  wire        _GEN_1929 = dis_ld_val_1 ? ~_GEN_1747 & ldq_20_bits_order_fail : ~_GEN_1609 & ldq_20_bits_order_fail;
  wire        _GEN_1930 = dis_ld_val_1 ? ~_GEN_1750 & ldq_21_bits_order_fail : ~_GEN_1610 & ldq_21_bits_order_fail;
  wire        _GEN_1931 = dis_ld_val_1 ? ~_GEN_1753 & ldq_22_bits_order_fail : ~_GEN_1611 & ldq_22_bits_order_fail;
  wire        _GEN_1932 = dis_ld_val_1 ? ~_GEN_1756 & ldq_23_bits_order_fail : ~_GEN_1612 & ldq_23_bits_order_fail;
  wire        _GEN_1933 = dis_ld_val_1 ? ~_GEN_1759 & ldq_24_bits_order_fail : ~_GEN_1613 & ldq_24_bits_order_fail;
  wire        _GEN_1934 = dis_ld_val_1 ? ~_GEN_1762 & ldq_25_bits_order_fail : ~_GEN_1614 & ldq_25_bits_order_fail;
  wire        _GEN_1935 = dis_ld_val_1 ? ~_GEN_1765 & ldq_26_bits_order_fail : ~_GEN_1615 & ldq_26_bits_order_fail;
  wire        _GEN_1936 = dis_ld_val_1 ? ~_GEN_1768 & ldq_27_bits_order_fail : ~_GEN_1616 & ldq_27_bits_order_fail;
  wire        _GEN_1937 = dis_ld_val_1 ? ~_GEN_1771 & ldq_28_bits_order_fail : ~_GEN_1617 & ldq_28_bits_order_fail;
  wire        _GEN_1938 = dis_ld_val_1 ? ~_GEN_1774 & ldq_29_bits_order_fail : ~_GEN_1618 & ldq_29_bits_order_fail;
  wire        _GEN_1939 = dis_ld_val_1 ? ~_GEN_1777 & ldq_30_bits_order_fail : ~_GEN_1619 & ldq_30_bits_order_fail;
  wire        _GEN_1940 = dis_ld_val_1 ? ~_GEN_1779 & ldq_31_bits_order_fail : ~_GEN_1620 & ldq_31_bits_order_fail;
  wire        _GEN_1941 = dis_ld_val_1 ? ~_GEN_1687 & ldq_0_bits_observed : ~_GEN_1589 & ldq_0_bits_observed;
  wire        _GEN_1942 = dis_ld_val_1 ? ~_GEN_1690 & ldq_1_bits_observed : ~_GEN_1590 & ldq_1_bits_observed;
  wire        _GEN_1943 = dis_ld_val_1 ? ~_GEN_1693 & ldq_2_bits_observed : ~_GEN_1591 & ldq_2_bits_observed;
  wire        _GEN_1944 = dis_ld_val_1 ? ~_GEN_1696 & ldq_3_bits_observed : ~_GEN_1592 & ldq_3_bits_observed;
  wire        _GEN_1945 = dis_ld_val_1 ? ~_GEN_1699 & ldq_4_bits_observed : ~_GEN_1593 & ldq_4_bits_observed;
  wire        _GEN_1946 = dis_ld_val_1 ? ~_GEN_1702 & ldq_5_bits_observed : ~_GEN_1594 & ldq_5_bits_observed;
  wire        _GEN_1947 = dis_ld_val_1 ? ~_GEN_1705 & ldq_6_bits_observed : ~_GEN_1595 & ldq_6_bits_observed;
  wire        _GEN_1948 = dis_ld_val_1 ? ~_GEN_1708 & ldq_7_bits_observed : ~_GEN_1596 & ldq_7_bits_observed;
  wire        _GEN_1949 = dis_ld_val_1 ? ~_GEN_1711 & ldq_8_bits_observed : ~_GEN_1597 & ldq_8_bits_observed;
  wire        _GEN_1950 = dis_ld_val_1 ? ~_GEN_1714 & ldq_9_bits_observed : ~_GEN_1598 & ldq_9_bits_observed;
  wire        _GEN_1951 = dis_ld_val_1 ? ~_GEN_1717 & ldq_10_bits_observed : ~_GEN_1599 & ldq_10_bits_observed;
  wire        _GEN_1952 = dis_ld_val_1 ? ~_GEN_1720 & ldq_11_bits_observed : ~_GEN_1600 & ldq_11_bits_observed;
  wire        _GEN_1953 = dis_ld_val_1 ? ~_GEN_1723 & ldq_12_bits_observed : ~_GEN_1601 & ldq_12_bits_observed;
  wire        _GEN_1954 = dis_ld_val_1 ? ~_GEN_1726 & ldq_13_bits_observed : ~_GEN_1602 & ldq_13_bits_observed;
  wire        _GEN_1955 = dis_ld_val_1 ? ~_GEN_1729 & ldq_14_bits_observed : ~_GEN_1603 & ldq_14_bits_observed;
  wire        _GEN_1956 = dis_ld_val_1 ? ~_GEN_1732 & ldq_15_bits_observed : ~_GEN_1604 & ldq_15_bits_observed;
  wire        _GEN_1957 = dis_ld_val_1 ? ~_GEN_1735 & ldq_16_bits_observed : ~_GEN_1605 & ldq_16_bits_observed;
  wire        _GEN_1958 = dis_ld_val_1 ? ~_GEN_1738 & ldq_17_bits_observed : ~_GEN_1606 & ldq_17_bits_observed;
  wire        _GEN_1959 = dis_ld_val_1 ? ~_GEN_1741 & ldq_18_bits_observed : ~_GEN_1607 & ldq_18_bits_observed;
  wire        _GEN_1960 = dis_ld_val_1 ? ~_GEN_1744 & ldq_19_bits_observed : ~_GEN_1608 & ldq_19_bits_observed;
  wire        _GEN_1961 = dis_ld_val_1 ? ~_GEN_1747 & ldq_20_bits_observed : ~_GEN_1609 & ldq_20_bits_observed;
  wire        _GEN_1962 = dis_ld_val_1 ? ~_GEN_1750 & ldq_21_bits_observed : ~_GEN_1610 & ldq_21_bits_observed;
  wire        _GEN_1963 = dis_ld_val_1 ? ~_GEN_1753 & ldq_22_bits_observed : ~_GEN_1611 & ldq_22_bits_observed;
  wire        _GEN_1964 = dis_ld_val_1 ? ~_GEN_1756 & ldq_23_bits_observed : ~_GEN_1612 & ldq_23_bits_observed;
  wire        _GEN_1965 = dis_ld_val_1 ? ~_GEN_1759 & ldq_24_bits_observed : ~_GEN_1613 & ldq_24_bits_observed;
  wire        _GEN_1966 = dis_ld_val_1 ? ~_GEN_1762 & ldq_25_bits_observed : ~_GEN_1614 & ldq_25_bits_observed;
  wire        _GEN_1967 = dis_ld_val_1 ? ~_GEN_1765 & ldq_26_bits_observed : ~_GEN_1615 & ldq_26_bits_observed;
  wire        _GEN_1968 = dis_ld_val_1 ? ~_GEN_1768 & ldq_27_bits_observed : ~_GEN_1616 & ldq_27_bits_observed;
  wire        _GEN_1969 = dis_ld_val_1 ? ~_GEN_1771 & ldq_28_bits_observed : ~_GEN_1617 & ldq_28_bits_observed;
  wire        _GEN_1970 = dis_ld_val_1 ? ~_GEN_1774 & ldq_29_bits_observed : ~_GEN_1618 & ldq_29_bits_observed;
  wire        _GEN_1971 = dis_ld_val_1 ? ~_GEN_1777 & ldq_30_bits_observed : ~_GEN_1619 & ldq_30_bits_observed;
  wire        _GEN_1972 = dis_ld_val_1 ? ~_GEN_1779 & ldq_31_bits_observed : ~_GEN_1620 & ldq_31_bits_observed;
  wire        _GEN_1973 = dis_ld_val_1 ? ~_GEN_1687 & ldq_0_bits_forward_std_val : ~_GEN_1589 & ldq_0_bits_forward_std_val;
  wire        _GEN_1974 = dis_ld_val_1 ? ~_GEN_1690 & ldq_1_bits_forward_std_val : ~_GEN_1590 & ldq_1_bits_forward_std_val;
  wire        _GEN_1975 = dis_ld_val_1 ? ~_GEN_1693 & ldq_2_bits_forward_std_val : ~_GEN_1591 & ldq_2_bits_forward_std_val;
  wire        _GEN_1976 = dis_ld_val_1 ? ~_GEN_1696 & ldq_3_bits_forward_std_val : ~_GEN_1592 & ldq_3_bits_forward_std_val;
  wire        _GEN_1977 = dis_ld_val_1 ? ~_GEN_1699 & ldq_4_bits_forward_std_val : ~_GEN_1593 & ldq_4_bits_forward_std_val;
  wire        _GEN_1978 = dis_ld_val_1 ? ~_GEN_1702 & ldq_5_bits_forward_std_val : ~_GEN_1594 & ldq_5_bits_forward_std_val;
  wire        _GEN_1979 = dis_ld_val_1 ? ~_GEN_1705 & ldq_6_bits_forward_std_val : ~_GEN_1595 & ldq_6_bits_forward_std_val;
  wire        _GEN_1980 = dis_ld_val_1 ? ~_GEN_1708 & ldq_7_bits_forward_std_val : ~_GEN_1596 & ldq_7_bits_forward_std_val;
  wire        _GEN_1981 = dis_ld_val_1 ? ~_GEN_1711 & ldq_8_bits_forward_std_val : ~_GEN_1597 & ldq_8_bits_forward_std_val;
  wire        _GEN_1982 = dis_ld_val_1 ? ~_GEN_1714 & ldq_9_bits_forward_std_val : ~_GEN_1598 & ldq_9_bits_forward_std_val;
  wire        _GEN_1983 = dis_ld_val_1 ? ~_GEN_1717 & ldq_10_bits_forward_std_val : ~_GEN_1599 & ldq_10_bits_forward_std_val;
  wire        _GEN_1984 = dis_ld_val_1 ? ~_GEN_1720 & ldq_11_bits_forward_std_val : ~_GEN_1600 & ldq_11_bits_forward_std_val;
  wire        _GEN_1985 = dis_ld_val_1 ? ~_GEN_1723 & ldq_12_bits_forward_std_val : ~_GEN_1601 & ldq_12_bits_forward_std_val;
  wire        _GEN_1986 = dis_ld_val_1 ? ~_GEN_1726 & ldq_13_bits_forward_std_val : ~_GEN_1602 & ldq_13_bits_forward_std_val;
  wire        _GEN_1987 = dis_ld_val_1 ? ~_GEN_1729 & ldq_14_bits_forward_std_val : ~_GEN_1603 & ldq_14_bits_forward_std_val;
  wire        _GEN_1988 = dis_ld_val_1 ? ~_GEN_1732 & ldq_15_bits_forward_std_val : ~_GEN_1604 & ldq_15_bits_forward_std_val;
  wire        _GEN_1989 = dis_ld_val_1 ? ~_GEN_1735 & ldq_16_bits_forward_std_val : ~_GEN_1605 & ldq_16_bits_forward_std_val;
  wire        _GEN_1990 = dis_ld_val_1 ? ~_GEN_1738 & ldq_17_bits_forward_std_val : ~_GEN_1606 & ldq_17_bits_forward_std_val;
  wire        _GEN_1991 = dis_ld_val_1 ? ~_GEN_1741 & ldq_18_bits_forward_std_val : ~_GEN_1607 & ldq_18_bits_forward_std_val;
  wire        _GEN_1992 = dis_ld_val_1 ? ~_GEN_1744 & ldq_19_bits_forward_std_val : ~_GEN_1608 & ldq_19_bits_forward_std_val;
  wire        _GEN_1993 = dis_ld_val_1 ? ~_GEN_1747 & ldq_20_bits_forward_std_val : ~_GEN_1609 & ldq_20_bits_forward_std_val;
  wire        _GEN_1994 = dis_ld_val_1 ? ~_GEN_1750 & ldq_21_bits_forward_std_val : ~_GEN_1610 & ldq_21_bits_forward_std_val;
  wire        _GEN_1995 = dis_ld_val_1 ? ~_GEN_1753 & ldq_22_bits_forward_std_val : ~_GEN_1611 & ldq_22_bits_forward_std_val;
  wire        _GEN_1996 = dis_ld_val_1 ? ~_GEN_1756 & ldq_23_bits_forward_std_val : ~_GEN_1612 & ldq_23_bits_forward_std_val;
  wire        _GEN_1997 = dis_ld_val_1 ? ~_GEN_1759 & ldq_24_bits_forward_std_val : ~_GEN_1613 & ldq_24_bits_forward_std_val;
  wire        _GEN_1998 = dis_ld_val_1 ? ~_GEN_1762 & ldq_25_bits_forward_std_val : ~_GEN_1614 & ldq_25_bits_forward_std_val;
  wire        _GEN_1999 = dis_ld_val_1 ? ~_GEN_1765 & ldq_26_bits_forward_std_val : ~_GEN_1615 & ldq_26_bits_forward_std_val;
  wire        _GEN_2000 = dis_ld_val_1 ? ~_GEN_1768 & ldq_27_bits_forward_std_val : ~_GEN_1616 & ldq_27_bits_forward_std_val;
  wire        _GEN_2001 = dis_ld_val_1 ? ~_GEN_1771 & ldq_28_bits_forward_std_val : ~_GEN_1617 & ldq_28_bits_forward_std_val;
  wire        _GEN_2002 = dis_ld_val_1 ? ~_GEN_1774 & ldq_29_bits_forward_std_val : ~_GEN_1618 & ldq_29_bits_forward_std_val;
  wire        _GEN_2003 = dis_ld_val_1 ? ~_GEN_1777 & ldq_30_bits_forward_std_val : ~_GEN_1619 & ldq_30_bits_forward_std_val;
  wire        _GEN_2004 = dis_ld_val_1 ? ~_GEN_1779 & ldq_31_bits_forward_std_val : ~_GEN_1620 & ldq_31_bits_forward_std_val;
  wire        _GEN_2005 = dis_st_val_1 & _GEN_6 == 5'h0;
  wire        _GEN_2006 = dis_st_val_1 & _GEN_6 == 5'h1;
  wire        _GEN_2007 = dis_st_val_1 & _GEN_6 == 5'h2;
  wire        _GEN_2008 = dis_st_val_1 & _GEN_6 == 5'h3;
  wire        _GEN_2009 = dis_st_val_1 & _GEN_6 == 5'h4;
  wire        _GEN_2010 = dis_st_val_1 & _GEN_6 == 5'h5;
  wire        _GEN_2011 = dis_st_val_1 & _GEN_6 == 5'h6;
  wire        _GEN_2012 = dis_st_val_1 & _GEN_6 == 5'h7;
  wire        _GEN_2013 = dis_st_val_1 & _GEN_6 == 5'h8;
  wire        _GEN_2014 = dis_st_val_1 & _GEN_6 == 5'h9;
  wire        _GEN_2015 = dis_st_val_1 & _GEN_6 == 5'hA;
  wire        _GEN_2016 = dis_st_val_1 & _GEN_6 == 5'hB;
  wire        _GEN_2017 = dis_st_val_1 & _GEN_6 == 5'hC;
  wire        _GEN_2018 = dis_st_val_1 & _GEN_6 == 5'hD;
  wire        _GEN_2019 = dis_st_val_1 & _GEN_6 == 5'hE;
  wire        _GEN_2020 = dis_st_val_1 & _GEN_6 == 5'hF;
  wire        _GEN_2021 = dis_st_val_1 & _GEN_6 == 5'h10;
  wire        _GEN_2022 = dis_st_val_1 & _GEN_6 == 5'h11;
  wire        _GEN_2023 = dis_st_val_1 & _GEN_6 == 5'h12;
  wire        _GEN_2024 = dis_st_val_1 & _GEN_6 == 5'h13;
  wire        _GEN_2025 = dis_st_val_1 & _GEN_6 == 5'h14;
  wire        _GEN_2026 = dis_st_val_1 & _GEN_6 == 5'h15;
  wire        _GEN_2027 = dis_st_val_1 & _GEN_6 == 5'h16;
  wire        _GEN_2028 = dis_st_val_1 & _GEN_6 == 5'h17;
  wire        _GEN_2029 = dis_st_val_1 & _GEN_6 == 5'h18;
  wire        _GEN_2030 = dis_st_val_1 & _GEN_6 == 5'h19;
  wire        _GEN_2031 = dis_st_val_1 & _GEN_6 == 5'h1A;
  wire        _GEN_2032 = dis_st_val_1 & _GEN_6 == 5'h1B;
  wire        _GEN_2033 = dis_st_val_1 & _GEN_6 == 5'h1C;
  wire        _GEN_2034 = dis_st_val_1 & _GEN_6 == 5'h1D;
  wire        _GEN_2035 = dis_st_val_1 & _GEN_6 == 5'h1E;
  wire        _GEN_2036 = dis_st_val_1 & (&_GEN_6);
  wire        _GEN_2037 = dis_ld_val_1 | ~_GEN_2005;
  wire        _GEN_2038 = dis_ld_val_1 | ~_GEN_2006;
  wire        _GEN_2039 = dis_ld_val_1 | ~_GEN_2007;
  wire        _GEN_2040 = dis_ld_val_1 | ~_GEN_2008;
  wire        _GEN_2041 = dis_ld_val_1 | ~_GEN_2009;
  wire        _GEN_2042 = dis_ld_val_1 | ~_GEN_2010;
  wire        _GEN_2043 = dis_ld_val_1 | ~_GEN_2011;
  wire        _GEN_2044 = dis_ld_val_1 | ~_GEN_2012;
  wire        _GEN_2045 = dis_ld_val_1 | ~_GEN_2013;
  wire        _GEN_2046 = dis_ld_val_1 | ~_GEN_2014;
  wire        _GEN_2047 = dis_ld_val_1 | ~_GEN_2015;
  wire        _GEN_2048 = dis_ld_val_1 | ~_GEN_2016;
  wire        _GEN_2049 = dis_ld_val_1 | ~_GEN_2017;
  wire        _GEN_2050 = dis_ld_val_1 | ~_GEN_2018;
  wire        _GEN_2051 = dis_ld_val_1 | ~_GEN_2019;
  wire        _GEN_2052 = dis_ld_val_1 | ~_GEN_2020;
  wire        _GEN_2053 = dis_ld_val_1 | ~_GEN_2021;
  wire        _GEN_2054 = dis_ld_val_1 | ~_GEN_2022;
  wire        _GEN_2055 = dis_ld_val_1 | ~_GEN_2023;
  wire        _GEN_2056 = dis_ld_val_1 | ~_GEN_2024;
  wire        _GEN_2057 = dis_ld_val_1 | ~_GEN_2025;
  wire        _GEN_2058 = dis_ld_val_1 | ~_GEN_2026;
  wire        _GEN_2059 = dis_ld_val_1 | ~_GEN_2027;
  wire        _GEN_2060 = dis_ld_val_1 | ~_GEN_2028;
  wire        _GEN_2061 = dis_ld_val_1 | ~_GEN_2029;
  wire        _GEN_2062 = dis_ld_val_1 | ~_GEN_2030;
  wire        _GEN_2063 = dis_ld_val_1 | ~_GEN_2031;
  wire        _GEN_2064 = dis_ld_val_1 | ~_GEN_2032;
  wire        _GEN_2065 = dis_ld_val_1 | ~_GEN_2033;
  wire        _GEN_2066 = dis_ld_val_1 | ~_GEN_2034;
  wire        _GEN_2067 = dis_ld_val_1 | ~_GEN_2035;
  wire        _GEN_2068 = dis_ld_val_1 | ~_GEN_2036;
  wire [31:0] _GEN_2069 = {32{dis_st_val_1}} & 32'h1 << _GEN_6 | _GEN_1685;
  wire        _GEN_2070 = dis_ld_val_2 & _GEN_9 == 5'h0;
  wire        _GEN_2071 = dis_ld_val_2 & _GEN_9 == 5'h1;
  wire        _GEN_2072 = dis_ld_val_2 & _GEN_9 == 5'h2;
  wire        _GEN_2073 = dis_ld_val_2 & _GEN_9 == 5'h3;
  wire        _GEN_2074 = dis_ld_val_2 & _GEN_9 == 5'h4;
  wire        _GEN_2075 = dis_ld_val_2 & _GEN_9 == 5'h5;
  wire        _GEN_2076 = dis_ld_val_2 & _GEN_9 == 5'h6;
  wire        _GEN_2077 = dis_ld_val_2 & _GEN_9 == 5'h7;
  wire        _GEN_2078 = dis_ld_val_2 & _GEN_9 == 5'h8;
  wire        _GEN_2079 = dis_ld_val_2 & _GEN_9 == 5'h9;
  wire        _GEN_2080 = dis_ld_val_2 & _GEN_9 == 5'hA;
  wire        _GEN_2081 = dis_ld_val_2 & _GEN_9 == 5'hB;
  wire        _GEN_2082 = dis_ld_val_2 & _GEN_9 == 5'hC;
  wire        _GEN_2083 = dis_ld_val_2 & _GEN_9 == 5'hD;
  wire        _GEN_2084 = dis_ld_val_2 & _GEN_9 == 5'hE;
  wire        _GEN_2085 = dis_ld_val_2 & _GEN_9 == 5'hF;
  wire        _GEN_2086 = dis_ld_val_2 & _GEN_9 == 5'h10;
  wire        _GEN_2087 = dis_ld_val_2 & _GEN_9 == 5'h11;
  wire        _GEN_2088 = dis_ld_val_2 & _GEN_9 == 5'h12;
  wire        _GEN_2089 = dis_ld_val_2 & _GEN_9 == 5'h13;
  wire        _GEN_2090 = dis_ld_val_2 & _GEN_9 == 5'h14;
  wire        _GEN_2091 = dis_ld_val_2 & _GEN_9 == 5'h15;
  wire        _GEN_2092 = dis_ld_val_2 & _GEN_9 == 5'h16;
  wire        _GEN_2093 = dis_ld_val_2 & _GEN_9 == 5'h17;
  wire        _GEN_2094 = dis_ld_val_2 & _GEN_9 == 5'h18;
  wire        _GEN_2095 = dis_ld_val_2 & _GEN_9 == 5'h19;
  wire        _GEN_2096 = dis_ld_val_2 & _GEN_9 == 5'h1A;
  wire        _GEN_2097 = dis_ld_val_2 & _GEN_9 == 5'h1B;
  wire        _GEN_2098 = dis_ld_val_2 & _GEN_9 == 5'h1C;
  wire        _GEN_2099 = dis_ld_val_2 & _GEN_9 == 5'h1D;
  wire        _GEN_2100 = dis_ld_val_2 & _GEN_9 == 5'h1E;
  wire        _GEN_2101 = dis_ld_val_2 & (&_GEN_9);
  wire        _GEN_2102 = dis_st_val_2 & _GEN_10 == 5'h0;
  wire        _GEN_2103 = dis_st_val_2 & _GEN_10 == 5'h1;
  wire        _GEN_2104 = dis_st_val_2 & _GEN_10 == 5'h2;
  wire        _GEN_2105 = dis_st_val_2 & _GEN_10 == 5'h3;
  wire        _GEN_2106 = dis_st_val_2 & _GEN_10 == 5'h4;
  wire        _GEN_2107 = dis_st_val_2 & _GEN_10 == 5'h5;
  wire        _GEN_2108 = dis_st_val_2 & _GEN_10 == 5'h6;
  wire        _GEN_2109 = dis_st_val_2 & _GEN_10 == 5'h7;
  wire        _GEN_2110 = dis_st_val_2 & _GEN_10 == 5'h8;
  wire        _GEN_2111 = dis_st_val_2 & _GEN_10 == 5'h9;
  wire        _GEN_2112 = dis_st_val_2 & _GEN_10 == 5'hA;
  wire        _GEN_2113 = dis_st_val_2 & _GEN_10 == 5'hB;
  wire        _GEN_2114 = dis_st_val_2 & _GEN_10 == 5'hC;
  wire        _GEN_2115 = dis_st_val_2 & _GEN_10 == 5'hD;
  wire        _GEN_2116 = dis_st_val_2 & _GEN_10 == 5'hE;
  wire        _GEN_2117 = dis_st_val_2 & _GEN_10 == 5'hF;
  wire        _GEN_2118 = dis_st_val_2 & _GEN_10 == 5'h10;
  wire        _GEN_2119 = dis_st_val_2 & _GEN_10 == 5'h11;
  wire        _GEN_2120 = dis_st_val_2 & _GEN_10 == 5'h12;
  wire        _GEN_2121 = dis_st_val_2 & _GEN_10 == 5'h13;
  wire        _GEN_2122 = dis_st_val_2 & _GEN_10 == 5'h14;
  wire        _GEN_2123 = dis_st_val_2 & _GEN_10 == 5'h15;
  wire        _GEN_2124 = dis_st_val_2 & _GEN_10 == 5'h16;
  wire        _GEN_2125 = dis_st_val_2 & _GEN_10 == 5'h17;
  wire        _GEN_2126 = dis_st_val_2 & _GEN_10 == 5'h18;
  wire        _GEN_2127 = dis_st_val_2 & _GEN_10 == 5'h19;
  wire        _GEN_2128 = dis_st_val_2 & _GEN_10 == 5'h1A;
  wire        _GEN_2129 = dis_st_val_2 & _GEN_10 == 5'h1B;
  wire        _GEN_2130 = dis_st_val_2 & _GEN_10 == 5'h1C;
  wire        _GEN_2131 = dis_st_val_2 & _GEN_10 == 5'h1D;
  wire        _GEN_2132 = dis_st_val_2 & _GEN_10 == 5'h1E;
  wire        _GEN_2133 = dis_st_val_2 & (&_GEN_10);
  wire        _GEN_2134 = dis_ld_val_2 | ~_GEN_2102;
  wire        _GEN_2135 = dis_ld_val_2 | ~_GEN_2103;
  wire        _GEN_2136 = dis_ld_val_2 | ~_GEN_2104;
  wire        _GEN_2137 = dis_ld_val_2 | ~_GEN_2105;
  wire        _GEN_2138 = dis_ld_val_2 | ~_GEN_2106;
  wire        _GEN_2139 = dis_ld_val_2 | ~_GEN_2107;
  wire        _GEN_2140 = dis_ld_val_2 | ~_GEN_2108;
  wire        _GEN_2141 = dis_ld_val_2 | ~_GEN_2109;
  wire        _GEN_2142 = dis_ld_val_2 | ~_GEN_2110;
  wire        _GEN_2143 = dis_ld_val_2 | ~_GEN_2111;
  wire        _GEN_2144 = dis_ld_val_2 | ~_GEN_2112;
  wire        _GEN_2145 = dis_ld_val_2 | ~_GEN_2113;
  wire        _GEN_2146 = dis_ld_val_2 | ~_GEN_2114;
  wire        _GEN_2147 = dis_ld_val_2 | ~_GEN_2115;
  wire        _GEN_2148 = dis_ld_val_2 | ~_GEN_2116;
  wire        _GEN_2149 = dis_ld_val_2 | ~_GEN_2117;
  wire        _GEN_2150 = dis_ld_val_2 | ~_GEN_2118;
  wire        _GEN_2151 = dis_ld_val_2 | ~_GEN_2119;
  wire        _GEN_2152 = dis_ld_val_2 | ~_GEN_2120;
  wire        _GEN_2153 = dis_ld_val_2 | ~_GEN_2121;
  wire        _GEN_2154 = dis_ld_val_2 | ~_GEN_2122;
  wire        _GEN_2155 = dis_ld_val_2 | ~_GEN_2123;
  wire        _GEN_2156 = dis_ld_val_2 | ~_GEN_2124;
  wire        _GEN_2157 = dis_ld_val_2 | ~_GEN_2125;
  wire        _GEN_2158 = dis_ld_val_2 | ~_GEN_2126;
  wire        _GEN_2159 = dis_ld_val_2 | ~_GEN_2127;
  wire        _GEN_2160 = dis_ld_val_2 | ~_GEN_2128;
  wire        _GEN_2161 = dis_ld_val_2 | ~_GEN_2129;
  wire        _GEN_2162 = dis_ld_val_2 | ~_GEN_2130;
  wire        _GEN_2163 = dis_ld_val_2 | ~_GEN_2131;
  wire        _GEN_2164 = dis_ld_val_2 | ~_GEN_2132;
  wire        _GEN_2165 = dis_ld_val_2 | ~_GEN_2133;
  wire [31:0] _GEN_2166 = {32{dis_st_val_2}} & 32'h1 << _GEN_10 | _GEN_2069;
  wire        _GEN_2167 = _GEN_13 == 5'h0;
  wire        _GEN_2168 = _GEN_2167 | _GEN_2070;
  wire        _GEN_2169 = dis_ld_val_3 ? _GEN_2168 | _GEN_1688 : _GEN_2070 | _GEN_1688;
  wire        _GEN_2170 = _GEN_13 == 5'h1;
  wire        _GEN_2171 = _GEN_2170 | _GEN_2071;
  wire        _GEN_2172 = dis_ld_val_3 ? _GEN_2171 | _GEN_1691 : _GEN_2071 | _GEN_1691;
  wire        _GEN_2173 = _GEN_13 == 5'h2;
  wire        _GEN_2174 = _GEN_2173 | _GEN_2072;
  wire        _GEN_2175 = dis_ld_val_3 ? _GEN_2174 | _GEN_1694 : _GEN_2072 | _GEN_1694;
  wire        _GEN_2176 = _GEN_13 == 5'h3;
  wire        _GEN_2177 = _GEN_2176 | _GEN_2073;
  wire        _GEN_2178 = dis_ld_val_3 ? _GEN_2177 | _GEN_1697 : _GEN_2073 | _GEN_1697;
  wire        _GEN_2179 = _GEN_13 == 5'h4;
  wire        _GEN_2180 = _GEN_2179 | _GEN_2074;
  wire        _GEN_2181 = dis_ld_val_3 ? _GEN_2180 | _GEN_1700 : _GEN_2074 | _GEN_1700;
  wire        _GEN_2182 = _GEN_13 == 5'h5;
  wire        _GEN_2183 = _GEN_2182 | _GEN_2075;
  wire        _GEN_2184 = dis_ld_val_3 ? _GEN_2183 | _GEN_1703 : _GEN_2075 | _GEN_1703;
  wire        _GEN_2185 = _GEN_13 == 5'h6;
  wire        _GEN_2186 = _GEN_2185 | _GEN_2076;
  wire        _GEN_2187 = dis_ld_val_3 ? _GEN_2186 | _GEN_1706 : _GEN_2076 | _GEN_1706;
  wire        _GEN_2188 = _GEN_13 == 5'h7;
  wire        _GEN_2189 = _GEN_2188 | _GEN_2077;
  wire        _GEN_2190 = dis_ld_val_3 ? _GEN_2189 | _GEN_1709 : _GEN_2077 | _GEN_1709;
  wire        _GEN_2191 = _GEN_13 == 5'h8;
  wire        _GEN_2192 = _GEN_2191 | _GEN_2078;
  wire        _GEN_2193 = dis_ld_val_3 ? _GEN_2192 | _GEN_1712 : _GEN_2078 | _GEN_1712;
  wire        _GEN_2194 = _GEN_13 == 5'h9;
  wire        _GEN_2195 = _GEN_2194 | _GEN_2079;
  wire        _GEN_2196 = dis_ld_val_3 ? _GEN_2195 | _GEN_1715 : _GEN_2079 | _GEN_1715;
  wire        _GEN_2197 = _GEN_13 == 5'hA;
  wire        _GEN_2198 = _GEN_2197 | _GEN_2080;
  wire        _GEN_2199 = dis_ld_val_3 ? _GEN_2198 | _GEN_1718 : _GEN_2080 | _GEN_1718;
  wire        _GEN_2200 = _GEN_13 == 5'hB;
  wire        _GEN_2201 = _GEN_2200 | _GEN_2081;
  wire        _GEN_2202 = dis_ld_val_3 ? _GEN_2201 | _GEN_1721 : _GEN_2081 | _GEN_1721;
  wire        _GEN_2203 = _GEN_13 == 5'hC;
  wire        _GEN_2204 = _GEN_2203 | _GEN_2082;
  wire        _GEN_2205 = dis_ld_val_3 ? _GEN_2204 | _GEN_1724 : _GEN_2082 | _GEN_1724;
  wire        _GEN_2206 = _GEN_13 == 5'hD;
  wire        _GEN_2207 = _GEN_2206 | _GEN_2083;
  wire        _GEN_2208 = dis_ld_val_3 ? _GEN_2207 | _GEN_1727 : _GEN_2083 | _GEN_1727;
  wire        _GEN_2209 = _GEN_13 == 5'hE;
  wire        _GEN_2210 = _GEN_2209 | _GEN_2084;
  wire        _GEN_2211 = dis_ld_val_3 ? _GEN_2210 | _GEN_1730 : _GEN_2084 | _GEN_1730;
  wire        _GEN_2212 = _GEN_13 == 5'hF;
  wire        _GEN_2213 = _GEN_2212 | _GEN_2085;
  wire        _GEN_2214 = dis_ld_val_3 ? _GEN_2213 | _GEN_1733 : _GEN_2085 | _GEN_1733;
  wire        _GEN_2215 = _GEN_13 == 5'h10;
  wire        _GEN_2216 = _GEN_2215 | _GEN_2086;
  wire        _GEN_2217 = dis_ld_val_3 ? _GEN_2216 | _GEN_1736 : _GEN_2086 | _GEN_1736;
  wire        _GEN_2218 = _GEN_13 == 5'h11;
  wire        _GEN_2219 = _GEN_2218 | _GEN_2087;
  wire        _GEN_2220 = dis_ld_val_3 ? _GEN_2219 | _GEN_1739 : _GEN_2087 | _GEN_1739;
  wire        _GEN_2221 = _GEN_13 == 5'h12;
  wire        _GEN_2222 = _GEN_2221 | _GEN_2088;
  wire        _GEN_2223 = dis_ld_val_3 ? _GEN_2222 | _GEN_1742 : _GEN_2088 | _GEN_1742;
  wire        _GEN_2224 = _GEN_13 == 5'h13;
  wire        _GEN_2225 = _GEN_2224 | _GEN_2089;
  wire        _GEN_2226 = dis_ld_val_3 ? _GEN_2225 | _GEN_1745 : _GEN_2089 | _GEN_1745;
  wire        _GEN_2227 = _GEN_13 == 5'h14;
  wire        _GEN_2228 = _GEN_2227 | _GEN_2090;
  wire        _GEN_2229 = dis_ld_val_3 ? _GEN_2228 | _GEN_1748 : _GEN_2090 | _GEN_1748;
  wire        _GEN_2230 = _GEN_13 == 5'h15;
  wire        _GEN_2231 = _GEN_2230 | _GEN_2091;
  wire        _GEN_2232 = dis_ld_val_3 ? _GEN_2231 | _GEN_1751 : _GEN_2091 | _GEN_1751;
  wire        _GEN_2233 = _GEN_13 == 5'h16;
  wire        _GEN_2234 = _GEN_2233 | _GEN_2092;
  wire        _GEN_2235 = dis_ld_val_3 ? _GEN_2234 | _GEN_1754 : _GEN_2092 | _GEN_1754;
  wire        _GEN_2236 = _GEN_13 == 5'h17;
  wire        _GEN_2237 = _GEN_2236 | _GEN_2093;
  wire        _GEN_2238 = dis_ld_val_3 ? _GEN_2237 | _GEN_1757 : _GEN_2093 | _GEN_1757;
  wire        _GEN_2239 = _GEN_13 == 5'h18;
  wire        _GEN_2240 = _GEN_2239 | _GEN_2094;
  wire        _GEN_2241 = dis_ld_val_3 ? _GEN_2240 | _GEN_1760 : _GEN_2094 | _GEN_1760;
  wire        _GEN_2242 = _GEN_13 == 5'h19;
  wire        _GEN_2243 = _GEN_2242 | _GEN_2095;
  wire        _GEN_2244 = dis_ld_val_3 ? _GEN_2243 | _GEN_1763 : _GEN_2095 | _GEN_1763;
  wire        _GEN_2245 = _GEN_13 == 5'h1A;
  wire        _GEN_2246 = _GEN_2245 | _GEN_2096;
  wire        _GEN_2247 = dis_ld_val_3 ? _GEN_2246 | _GEN_1766 : _GEN_2096 | _GEN_1766;
  wire        _GEN_2248 = _GEN_13 == 5'h1B;
  wire        _GEN_2249 = _GEN_2248 | _GEN_2097;
  wire        _GEN_2250 = dis_ld_val_3 ? _GEN_2249 | _GEN_1769 : _GEN_2097 | _GEN_1769;
  wire        _GEN_2251 = _GEN_13 == 5'h1C;
  wire        _GEN_2252 = _GEN_2251 | _GEN_2098;
  wire        _GEN_2253 = dis_ld_val_3 ? _GEN_2252 | _GEN_1772 : _GEN_2098 | _GEN_1772;
  wire        _GEN_2254 = _GEN_13 == 5'h1D;
  wire        _GEN_2255 = _GEN_2254 | _GEN_2099;
  wire        _GEN_2256 = dis_ld_val_3 ? _GEN_2255 | _GEN_1775 : _GEN_2099 | _GEN_1775;
  wire        _GEN_2257 = _GEN_13 == 5'h1E;
  wire        _GEN_2258 = _GEN_2257 | _GEN_2100;
  wire        _GEN_2259 = dis_ld_val_3 ? _GEN_2258 | _GEN_1778 : _GEN_2100 | _GEN_1778;
  wire        _GEN_2260 = (&_GEN_13) | _GEN_2101;
  wire        _GEN_2261 = dis_ld_val_3 ? _GEN_2260 | _GEN_1780 : _GEN_2101 | _GEN_1780;
  wire        _GEN_2262 = dis_ld_val_3 & _GEN_2167;
  wire        _GEN_2263 = _GEN_2262 ? io_core_dis_uops_3_bits_exception : _GEN_2070 ? io_core_dis_uops_2_bits_exception : _GEN_1781 ? io_core_dis_uops_1_bits_exception : _GEN_1589 ? io_core_dis_uops_0_bits_exception : ldq_0_bits_uop_exception;
  wire        _GEN_2264 = dis_ld_val_3 & _GEN_2170;
  wire        _GEN_2265 = _GEN_2264 ? io_core_dis_uops_3_bits_exception : _GEN_2071 ? io_core_dis_uops_2_bits_exception : _GEN_1782 ? io_core_dis_uops_1_bits_exception : _GEN_1590 ? io_core_dis_uops_0_bits_exception : ldq_1_bits_uop_exception;
  wire        _GEN_2266 = dis_ld_val_3 & _GEN_2173;
  wire        _GEN_2267 = _GEN_2266 ? io_core_dis_uops_3_bits_exception : _GEN_2072 ? io_core_dis_uops_2_bits_exception : _GEN_1783 ? io_core_dis_uops_1_bits_exception : _GEN_1591 ? io_core_dis_uops_0_bits_exception : ldq_2_bits_uop_exception;
  wire        _GEN_2268 = dis_ld_val_3 & _GEN_2176;
  wire        _GEN_2269 = _GEN_2268 ? io_core_dis_uops_3_bits_exception : _GEN_2073 ? io_core_dis_uops_2_bits_exception : _GEN_1784 ? io_core_dis_uops_1_bits_exception : _GEN_1592 ? io_core_dis_uops_0_bits_exception : ldq_3_bits_uop_exception;
  wire        _GEN_2270 = dis_ld_val_3 & _GEN_2179;
  wire        _GEN_2271 = _GEN_2270 ? io_core_dis_uops_3_bits_exception : _GEN_2074 ? io_core_dis_uops_2_bits_exception : _GEN_1785 ? io_core_dis_uops_1_bits_exception : _GEN_1593 ? io_core_dis_uops_0_bits_exception : ldq_4_bits_uop_exception;
  wire        _GEN_2272 = dis_ld_val_3 & _GEN_2182;
  wire        _GEN_2273 = _GEN_2272 ? io_core_dis_uops_3_bits_exception : _GEN_2075 ? io_core_dis_uops_2_bits_exception : _GEN_1786 ? io_core_dis_uops_1_bits_exception : _GEN_1594 ? io_core_dis_uops_0_bits_exception : ldq_5_bits_uop_exception;
  wire        _GEN_2274 = dis_ld_val_3 & _GEN_2185;
  wire        _GEN_2275 = _GEN_2274 ? io_core_dis_uops_3_bits_exception : _GEN_2076 ? io_core_dis_uops_2_bits_exception : _GEN_1787 ? io_core_dis_uops_1_bits_exception : _GEN_1595 ? io_core_dis_uops_0_bits_exception : ldq_6_bits_uop_exception;
  wire        _GEN_2276 = dis_ld_val_3 & _GEN_2188;
  wire        _GEN_2277 = _GEN_2276 ? io_core_dis_uops_3_bits_exception : _GEN_2077 ? io_core_dis_uops_2_bits_exception : _GEN_1788 ? io_core_dis_uops_1_bits_exception : _GEN_1596 ? io_core_dis_uops_0_bits_exception : ldq_7_bits_uop_exception;
  wire        _GEN_2278 = dis_ld_val_3 & _GEN_2191;
  wire        _GEN_2279 = _GEN_2278 ? io_core_dis_uops_3_bits_exception : _GEN_2078 ? io_core_dis_uops_2_bits_exception : _GEN_1789 ? io_core_dis_uops_1_bits_exception : _GEN_1597 ? io_core_dis_uops_0_bits_exception : ldq_8_bits_uop_exception;
  wire        _GEN_2280 = dis_ld_val_3 & _GEN_2194;
  wire        _GEN_2281 = _GEN_2280 ? io_core_dis_uops_3_bits_exception : _GEN_2079 ? io_core_dis_uops_2_bits_exception : _GEN_1790 ? io_core_dis_uops_1_bits_exception : _GEN_1598 ? io_core_dis_uops_0_bits_exception : ldq_9_bits_uop_exception;
  wire        _GEN_2282 = dis_ld_val_3 & _GEN_2197;
  wire        _GEN_2283 = _GEN_2282 ? io_core_dis_uops_3_bits_exception : _GEN_2080 ? io_core_dis_uops_2_bits_exception : _GEN_1791 ? io_core_dis_uops_1_bits_exception : _GEN_1599 ? io_core_dis_uops_0_bits_exception : ldq_10_bits_uop_exception;
  wire        _GEN_2284 = dis_ld_val_3 & _GEN_2200;
  wire        _GEN_2285 = _GEN_2284 ? io_core_dis_uops_3_bits_exception : _GEN_2081 ? io_core_dis_uops_2_bits_exception : _GEN_1792 ? io_core_dis_uops_1_bits_exception : _GEN_1600 ? io_core_dis_uops_0_bits_exception : ldq_11_bits_uop_exception;
  wire        _GEN_2286 = dis_ld_val_3 & _GEN_2203;
  wire        _GEN_2287 = _GEN_2286 ? io_core_dis_uops_3_bits_exception : _GEN_2082 ? io_core_dis_uops_2_bits_exception : _GEN_1793 ? io_core_dis_uops_1_bits_exception : _GEN_1601 ? io_core_dis_uops_0_bits_exception : ldq_12_bits_uop_exception;
  wire        _GEN_2288 = dis_ld_val_3 & _GEN_2206;
  wire        _GEN_2289 = _GEN_2288 ? io_core_dis_uops_3_bits_exception : _GEN_2083 ? io_core_dis_uops_2_bits_exception : _GEN_1794 ? io_core_dis_uops_1_bits_exception : _GEN_1602 ? io_core_dis_uops_0_bits_exception : ldq_13_bits_uop_exception;
  wire        _GEN_2290 = dis_ld_val_3 & _GEN_2209;
  wire        _GEN_2291 = _GEN_2290 ? io_core_dis_uops_3_bits_exception : _GEN_2084 ? io_core_dis_uops_2_bits_exception : _GEN_1795 ? io_core_dis_uops_1_bits_exception : _GEN_1603 ? io_core_dis_uops_0_bits_exception : ldq_14_bits_uop_exception;
  wire        _GEN_2292 = dis_ld_val_3 & _GEN_2212;
  wire        _GEN_2293 = _GEN_2292 ? io_core_dis_uops_3_bits_exception : _GEN_2085 ? io_core_dis_uops_2_bits_exception : _GEN_1796 ? io_core_dis_uops_1_bits_exception : _GEN_1604 ? io_core_dis_uops_0_bits_exception : ldq_15_bits_uop_exception;
  wire        _GEN_2294 = dis_ld_val_3 & _GEN_2215;
  wire        _GEN_2295 = _GEN_2294 ? io_core_dis_uops_3_bits_exception : _GEN_2086 ? io_core_dis_uops_2_bits_exception : _GEN_1797 ? io_core_dis_uops_1_bits_exception : _GEN_1605 ? io_core_dis_uops_0_bits_exception : ldq_16_bits_uop_exception;
  wire        _GEN_2296 = dis_ld_val_3 & _GEN_2218;
  wire        _GEN_2297 = _GEN_2296 ? io_core_dis_uops_3_bits_exception : _GEN_2087 ? io_core_dis_uops_2_bits_exception : _GEN_1798 ? io_core_dis_uops_1_bits_exception : _GEN_1606 ? io_core_dis_uops_0_bits_exception : ldq_17_bits_uop_exception;
  wire        _GEN_2298 = dis_ld_val_3 & _GEN_2221;
  wire        _GEN_2299 = _GEN_2298 ? io_core_dis_uops_3_bits_exception : _GEN_2088 ? io_core_dis_uops_2_bits_exception : _GEN_1799 ? io_core_dis_uops_1_bits_exception : _GEN_1607 ? io_core_dis_uops_0_bits_exception : ldq_18_bits_uop_exception;
  wire        _GEN_2300 = dis_ld_val_3 & _GEN_2224;
  wire        _GEN_2301 = _GEN_2300 ? io_core_dis_uops_3_bits_exception : _GEN_2089 ? io_core_dis_uops_2_bits_exception : _GEN_1800 ? io_core_dis_uops_1_bits_exception : _GEN_1608 ? io_core_dis_uops_0_bits_exception : ldq_19_bits_uop_exception;
  wire        _GEN_2302 = dis_ld_val_3 & _GEN_2227;
  wire        _GEN_2303 = _GEN_2302 ? io_core_dis_uops_3_bits_exception : _GEN_2090 ? io_core_dis_uops_2_bits_exception : _GEN_1801 ? io_core_dis_uops_1_bits_exception : _GEN_1609 ? io_core_dis_uops_0_bits_exception : ldq_20_bits_uop_exception;
  wire        _GEN_2304 = dis_ld_val_3 & _GEN_2230;
  wire        _GEN_2305 = _GEN_2304 ? io_core_dis_uops_3_bits_exception : _GEN_2091 ? io_core_dis_uops_2_bits_exception : _GEN_1802 ? io_core_dis_uops_1_bits_exception : _GEN_1610 ? io_core_dis_uops_0_bits_exception : ldq_21_bits_uop_exception;
  wire        _GEN_2306 = dis_ld_val_3 & _GEN_2233;
  wire        _GEN_2307 = _GEN_2306 ? io_core_dis_uops_3_bits_exception : _GEN_2092 ? io_core_dis_uops_2_bits_exception : _GEN_1803 ? io_core_dis_uops_1_bits_exception : _GEN_1611 ? io_core_dis_uops_0_bits_exception : ldq_22_bits_uop_exception;
  wire        _GEN_2308 = dis_ld_val_3 & _GEN_2236;
  wire        _GEN_2309 = _GEN_2308 ? io_core_dis_uops_3_bits_exception : _GEN_2093 ? io_core_dis_uops_2_bits_exception : _GEN_1804 ? io_core_dis_uops_1_bits_exception : _GEN_1612 ? io_core_dis_uops_0_bits_exception : ldq_23_bits_uop_exception;
  wire        _GEN_2310 = dis_ld_val_3 & _GEN_2239;
  wire        _GEN_2311 = _GEN_2310 ? io_core_dis_uops_3_bits_exception : _GEN_2094 ? io_core_dis_uops_2_bits_exception : _GEN_1805 ? io_core_dis_uops_1_bits_exception : _GEN_1613 ? io_core_dis_uops_0_bits_exception : ldq_24_bits_uop_exception;
  wire        _GEN_2312 = dis_ld_val_3 & _GEN_2242;
  wire        _GEN_2313 = _GEN_2312 ? io_core_dis_uops_3_bits_exception : _GEN_2095 ? io_core_dis_uops_2_bits_exception : _GEN_1806 ? io_core_dis_uops_1_bits_exception : _GEN_1614 ? io_core_dis_uops_0_bits_exception : ldq_25_bits_uop_exception;
  wire        _GEN_2314 = dis_ld_val_3 & _GEN_2245;
  wire        _GEN_2315 = _GEN_2314 ? io_core_dis_uops_3_bits_exception : _GEN_2096 ? io_core_dis_uops_2_bits_exception : _GEN_1807 ? io_core_dis_uops_1_bits_exception : _GEN_1615 ? io_core_dis_uops_0_bits_exception : ldq_26_bits_uop_exception;
  wire        _GEN_2316 = dis_ld_val_3 & _GEN_2248;
  wire        _GEN_2317 = _GEN_2316 ? io_core_dis_uops_3_bits_exception : _GEN_2097 ? io_core_dis_uops_2_bits_exception : _GEN_1808 ? io_core_dis_uops_1_bits_exception : _GEN_1616 ? io_core_dis_uops_0_bits_exception : ldq_27_bits_uop_exception;
  wire        _GEN_2318 = dis_ld_val_3 & _GEN_2251;
  wire        _GEN_2319 = _GEN_2318 ? io_core_dis_uops_3_bits_exception : _GEN_2098 ? io_core_dis_uops_2_bits_exception : _GEN_1809 ? io_core_dis_uops_1_bits_exception : _GEN_1617 ? io_core_dis_uops_0_bits_exception : ldq_28_bits_uop_exception;
  wire        _GEN_2320 = dis_ld_val_3 & _GEN_2254;
  wire        _GEN_2321 = _GEN_2320 ? io_core_dis_uops_3_bits_exception : _GEN_2099 ? io_core_dis_uops_2_bits_exception : _GEN_1810 ? io_core_dis_uops_1_bits_exception : _GEN_1618 ? io_core_dis_uops_0_bits_exception : ldq_29_bits_uop_exception;
  wire        _GEN_2322 = dis_ld_val_3 & _GEN_2257;
  wire        _GEN_2323 = _GEN_2322 ? io_core_dis_uops_3_bits_exception : _GEN_2100 ? io_core_dis_uops_2_bits_exception : _GEN_1811 ? io_core_dis_uops_1_bits_exception : _GEN_1619 ? io_core_dis_uops_0_bits_exception : ldq_30_bits_uop_exception;
  wire        _GEN_2324 = dis_ld_val_3 & (&_GEN_13);
  wire        _GEN_2325 = _GEN_2324 ? io_core_dis_uops_3_bits_exception : _GEN_2101 ? io_core_dis_uops_2_bits_exception : _GEN_1812 ? io_core_dis_uops_1_bits_exception : _GEN_1620 ? io_core_dis_uops_0_bits_exception : ldq_31_bits_uop_exception;
  wire        _GEN_2326 = dis_ld_val_3 ? ~_GEN_2168 & _GEN_1813 : ~_GEN_2070 & _GEN_1813;
  wire        _GEN_2327 = dis_ld_val_3 ? ~_GEN_2171 & _GEN_1814 : ~_GEN_2071 & _GEN_1814;
  wire        _GEN_2328 = dis_ld_val_3 ? ~_GEN_2174 & _GEN_1815 : ~_GEN_2072 & _GEN_1815;
  wire        _GEN_2329 = dis_ld_val_3 ? ~_GEN_2177 & _GEN_1816 : ~_GEN_2073 & _GEN_1816;
  wire        _GEN_2330 = dis_ld_val_3 ? ~_GEN_2180 & _GEN_1817 : ~_GEN_2074 & _GEN_1817;
  wire        _GEN_2331 = dis_ld_val_3 ? ~_GEN_2183 & _GEN_1818 : ~_GEN_2075 & _GEN_1818;
  wire        _GEN_2332 = dis_ld_val_3 ? ~_GEN_2186 & _GEN_1819 : ~_GEN_2076 & _GEN_1819;
  wire        _GEN_2333 = dis_ld_val_3 ? ~_GEN_2189 & _GEN_1820 : ~_GEN_2077 & _GEN_1820;
  wire        _GEN_2334 = dis_ld_val_3 ? ~_GEN_2192 & _GEN_1821 : ~_GEN_2078 & _GEN_1821;
  wire        _GEN_2335 = dis_ld_val_3 ? ~_GEN_2195 & _GEN_1822 : ~_GEN_2079 & _GEN_1822;
  wire        _GEN_2336 = dis_ld_val_3 ? ~_GEN_2198 & _GEN_1823 : ~_GEN_2080 & _GEN_1823;
  wire        _GEN_2337 = dis_ld_val_3 ? ~_GEN_2201 & _GEN_1824 : ~_GEN_2081 & _GEN_1824;
  wire        _GEN_2338 = dis_ld_val_3 ? ~_GEN_2204 & _GEN_1825 : ~_GEN_2082 & _GEN_1825;
  wire        _GEN_2339 = dis_ld_val_3 ? ~_GEN_2207 & _GEN_1826 : ~_GEN_2083 & _GEN_1826;
  wire        _GEN_2340 = dis_ld_val_3 ? ~_GEN_2210 & _GEN_1827 : ~_GEN_2084 & _GEN_1827;
  wire        _GEN_2341 = dis_ld_val_3 ? ~_GEN_2213 & _GEN_1828 : ~_GEN_2085 & _GEN_1828;
  wire        _GEN_2342 = dis_ld_val_3 ? ~_GEN_2216 & _GEN_1829 : ~_GEN_2086 & _GEN_1829;
  wire        _GEN_2343 = dis_ld_val_3 ? ~_GEN_2219 & _GEN_1830 : ~_GEN_2087 & _GEN_1830;
  wire        _GEN_2344 = dis_ld_val_3 ? ~_GEN_2222 & _GEN_1831 : ~_GEN_2088 & _GEN_1831;
  wire        _GEN_2345 = dis_ld_val_3 ? ~_GEN_2225 & _GEN_1832 : ~_GEN_2089 & _GEN_1832;
  wire        _GEN_2346 = dis_ld_val_3 ? ~_GEN_2228 & _GEN_1833 : ~_GEN_2090 & _GEN_1833;
  wire        _GEN_2347 = dis_ld_val_3 ? ~_GEN_2231 & _GEN_1834 : ~_GEN_2091 & _GEN_1834;
  wire        _GEN_2348 = dis_ld_val_3 ? ~_GEN_2234 & _GEN_1835 : ~_GEN_2092 & _GEN_1835;
  wire        _GEN_2349 = dis_ld_val_3 ? ~_GEN_2237 & _GEN_1836 : ~_GEN_2093 & _GEN_1836;
  wire        _GEN_2350 = dis_ld_val_3 ? ~_GEN_2240 & _GEN_1837 : ~_GEN_2094 & _GEN_1837;
  wire        _GEN_2351 = dis_ld_val_3 ? ~_GEN_2243 & _GEN_1838 : ~_GEN_2095 & _GEN_1838;
  wire        _GEN_2352 = dis_ld_val_3 ? ~_GEN_2246 & _GEN_1839 : ~_GEN_2096 & _GEN_1839;
  wire        _GEN_2353 = dis_ld_val_3 ? ~_GEN_2249 & _GEN_1840 : ~_GEN_2097 & _GEN_1840;
  wire        _GEN_2354 = dis_ld_val_3 ? ~_GEN_2252 & _GEN_1841 : ~_GEN_2098 & _GEN_1841;
  wire        _GEN_2355 = dis_ld_val_3 ? ~_GEN_2255 & _GEN_1842 : ~_GEN_2099 & _GEN_1842;
  wire        _GEN_2356 = dis_ld_val_3 ? ~_GEN_2258 & _GEN_1843 : ~_GEN_2100 & _GEN_1843;
  wire        _GEN_2357 = dis_ld_val_3 ? ~_GEN_2260 & _GEN_1844 : ~_GEN_2101 & _GEN_1844;
  wire        _GEN_2358 = dis_ld_val_3 ? ~_GEN_2168 & _GEN_1909 : ~_GEN_2070 & _GEN_1909;
  wire        _GEN_2359 = dis_ld_val_3 ? ~_GEN_2171 & _GEN_1910 : ~_GEN_2071 & _GEN_1910;
  wire        _GEN_2360 = dis_ld_val_3 ? ~_GEN_2174 & _GEN_1911 : ~_GEN_2072 & _GEN_1911;
  wire        _GEN_2361 = dis_ld_val_3 ? ~_GEN_2177 & _GEN_1912 : ~_GEN_2073 & _GEN_1912;
  wire        _GEN_2362 = dis_ld_val_3 ? ~_GEN_2180 & _GEN_1913 : ~_GEN_2074 & _GEN_1913;
  wire        _GEN_2363 = dis_ld_val_3 ? ~_GEN_2183 & _GEN_1914 : ~_GEN_2075 & _GEN_1914;
  wire        _GEN_2364 = dis_ld_val_3 ? ~_GEN_2186 & _GEN_1915 : ~_GEN_2076 & _GEN_1915;
  wire        _GEN_2365 = dis_ld_val_3 ? ~_GEN_2189 & _GEN_1916 : ~_GEN_2077 & _GEN_1916;
  wire        _GEN_2366 = dis_ld_val_3 ? ~_GEN_2192 & _GEN_1917 : ~_GEN_2078 & _GEN_1917;
  wire        _GEN_2367 = dis_ld_val_3 ? ~_GEN_2195 & _GEN_1918 : ~_GEN_2079 & _GEN_1918;
  wire        _GEN_2368 = dis_ld_val_3 ? ~_GEN_2198 & _GEN_1919 : ~_GEN_2080 & _GEN_1919;
  wire        _GEN_2369 = dis_ld_val_3 ? ~_GEN_2201 & _GEN_1920 : ~_GEN_2081 & _GEN_1920;
  wire        _GEN_2370 = dis_ld_val_3 ? ~_GEN_2204 & _GEN_1921 : ~_GEN_2082 & _GEN_1921;
  wire        _GEN_2371 = dis_ld_val_3 ? ~_GEN_2207 & _GEN_1922 : ~_GEN_2083 & _GEN_1922;
  wire        _GEN_2372 = dis_ld_val_3 ? ~_GEN_2210 & _GEN_1923 : ~_GEN_2084 & _GEN_1923;
  wire        _GEN_2373 = dis_ld_val_3 ? ~_GEN_2213 & _GEN_1924 : ~_GEN_2085 & _GEN_1924;
  wire        _GEN_2374 = dis_ld_val_3 ? ~_GEN_2216 & _GEN_1925 : ~_GEN_2086 & _GEN_1925;
  wire        _GEN_2375 = dis_ld_val_3 ? ~_GEN_2219 & _GEN_1926 : ~_GEN_2087 & _GEN_1926;
  wire        _GEN_2376 = dis_ld_val_3 ? ~_GEN_2222 & _GEN_1927 : ~_GEN_2088 & _GEN_1927;
  wire        _GEN_2377 = dis_ld_val_3 ? ~_GEN_2225 & _GEN_1928 : ~_GEN_2089 & _GEN_1928;
  wire        _GEN_2378 = dis_ld_val_3 ? ~_GEN_2228 & _GEN_1929 : ~_GEN_2090 & _GEN_1929;
  wire        _GEN_2379 = dis_ld_val_3 ? ~_GEN_2231 & _GEN_1930 : ~_GEN_2091 & _GEN_1930;
  wire        _GEN_2380 = dis_ld_val_3 ? ~_GEN_2234 & _GEN_1931 : ~_GEN_2092 & _GEN_1931;
  wire        _GEN_2381 = dis_ld_val_3 ? ~_GEN_2237 & _GEN_1932 : ~_GEN_2093 & _GEN_1932;
  wire        _GEN_2382 = dis_ld_val_3 ? ~_GEN_2240 & _GEN_1933 : ~_GEN_2094 & _GEN_1933;
  wire        _GEN_2383 = dis_ld_val_3 ? ~_GEN_2243 & _GEN_1934 : ~_GEN_2095 & _GEN_1934;
  wire        _GEN_2384 = dis_ld_val_3 ? ~_GEN_2246 & _GEN_1935 : ~_GEN_2096 & _GEN_1935;
  wire        _GEN_2385 = dis_ld_val_3 ? ~_GEN_2249 & _GEN_1936 : ~_GEN_2097 & _GEN_1936;
  wire        _GEN_2386 = dis_ld_val_3 ? ~_GEN_2252 & _GEN_1937 : ~_GEN_2098 & _GEN_1937;
  wire        _GEN_2387 = dis_ld_val_3 ? ~_GEN_2255 & _GEN_1938 : ~_GEN_2099 & _GEN_1938;
  wire        _GEN_2388 = dis_ld_val_3 ? ~_GEN_2258 & _GEN_1939 : ~_GEN_2100 & _GEN_1939;
  wire        _GEN_2389 = dis_ld_val_3 ? ~_GEN_2260 & _GEN_1940 : ~_GEN_2101 & _GEN_1940;
  wire        _GEN_2390 = dis_st_val_3 & _GEN_14 == 5'h0;
  wire        _GEN_2391 = ~dis_ld_val_3 & _GEN_2390 | ~dis_ld_val_2 & _GEN_2102 | ~dis_ld_val_1 & _GEN_2005 | ~dis_ld_val & _GEN_1621 | stq_0_valid;
  wire        _GEN_2392 = dis_st_val_3 & _GEN_14 == 5'h1;
  wire        _GEN_2393 = ~dis_ld_val_3 & _GEN_2392 | ~dis_ld_val_2 & _GEN_2103 | ~dis_ld_val_1 & _GEN_2006 | ~dis_ld_val & _GEN_1622 | stq_1_valid;
  wire        _GEN_2394 = dis_st_val_3 & _GEN_14 == 5'h2;
  wire        _GEN_2395 = ~dis_ld_val_3 & _GEN_2394 | ~dis_ld_val_2 & _GEN_2104 | ~dis_ld_val_1 & _GEN_2007 | ~dis_ld_val & _GEN_1623 | stq_2_valid;
  wire        _GEN_2396 = dis_st_val_3 & _GEN_14 == 5'h3;
  wire        _GEN_2397 = ~dis_ld_val_3 & _GEN_2396 | ~dis_ld_val_2 & _GEN_2105 | ~dis_ld_val_1 & _GEN_2008 | ~dis_ld_val & _GEN_1624 | stq_3_valid;
  wire        _GEN_2398 = dis_st_val_3 & _GEN_14 == 5'h4;
  wire        _GEN_2399 = ~dis_ld_val_3 & _GEN_2398 | ~dis_ld_val_2 & _GEN_2106 | ~dis_ld_val_1 & _GEN_2009 | ~dis_ld_val & _GEN_1625 | stq_4_valid;
  wire        _GEN_2400 = dis_st_val_3 & _GEN_14 == 5'h5;
  wire        _GEN_2401 = ~dis_ld_val_3 & _GEN_2400 | ~dis_ld_val_2 & _GEN_2107 | ~dis_ld_val_1 & _GEN_2010 | ~dis_ld_val & _GEN_1626 | stq_5_valid;
  wire        _GEN_2402 = dis_st_val_3 & _GEN_14 == 5'h6;
  wire        _GEN_2403 = ~dis_ld_val_3 & _GEN_2402 | ~dis_ld_val_2 & _GEN_2108 | ~dis_ld_val_1 & _GEN_2011 | ~dis_ld_val & _GEN_1627 | stq_6_valid;
  wire        _GEN_2404 = dis_st_val_3 & _GEN_14 == 5'h7;
  wire        _GEN_2405 = ~dis_ld_val_3 & _GEN_2404 | ~dis_ld_val_2 & _GEN_2109 | ~dis_ld_val_1 & _GEN_2012 | ~dis_ld_val & _GEN_1628 | stq_7_valid;
  wire        _GEN_2406 = dis_st_val_3 & _GEN_14 == 5'h8;
  wire        _GEN_2407 = ~dis_ld_val_3 & _GEN_2406 | ~dis_ld_val_2 & _GEN_2110 | ~dis_ld_val_1 & _GEN_2013 | ~dis_ld_val & _GEN_1629 | stq_8_valid;
  wire        _GEN_2408 = dis_st_val_3 & _GEN_14 == 5'h9;
  wire        _GEN_2409 = ~dis_ld_val_3 & _GEN_2408 | ~dis_ld_val_2 & _GEN_2111 | ~dis_ld_val_1 & _GEN_2014 | ~dis_ld_val & _GEN_1630 | stq_9_valid;
  wire        _GEN_2410 = dis_st_val_3 & _GEN_14 == 5'hA;
  wire        _GEN_2411 = ~dis_ld_val_3 & _GEN_2410 | ~dis_ld_val_2 & _GEN_2112 | ~dis_ld_val_1 & _GEN_2015 | ~dis_ld_val & _GEN_1631 | stq_10_valid;
  wire        _GEN_2412 = dis_st_val_3 & _GEN_14 == 5'hB;
  wire        _GEN_2413 = ~dis_ld_val_3 & _GEN_2412 | ~dis_ld_val_2 & _GEN_2113 | ~dis_ld_val_1 & _GEN_2016 | ~dis_ld_val & _GEN_1632 | stq_11_valid;
  wire        _GEN_2414 = dis_st_val_3 & _GEN_14 == 5'hC;
  wire        _GEN_2415 = ~dis_ld_val_3 & _GEN_2414 | ~dis_ld_val_2 & _GEN_2114 | ~dis_ld_val_1 & _GEN_2017 | ~dis_ld_val & _GEN_1633 | stq_12_valid;
  wire        _GEN_2416 = dis_st_val_3 & _GEN_14 == 5'hD;
  wire        _GEN_2417 = ~dis_ld_val_3 & _GEN_2416 | ~dis_ld_val_2 & _GEN_2115 | ~dis_ld_val_1 & _GEN_2018 | ~dis_ld_val & _GEN_1634 | stq_13_valid;
  wire        _GEN_2418 = dis_st_val_3 & _GEN_14 == 5'hE;
  wire        _GEN_2419 = ~dis_ld_val_3 & _GEN_2418 | ~dis_ld_val_2 & _GEN_2116 | ~dis_ld_val_1 & _GEN_2019 | ~dis_ld_val & _GEN_1635 | stq_14_valid;
  wire        _GEN_2420 = dis_st_val_3 & _GEN_14 == 5'hF;
  wire        _GEN_2421 = ~dis_ld_val_3 & _GEN_2420 | ~dis_ld_val_2 & _GEN_2117 | ~dis_ld_val_1 & _GEN_2020 | ~dis_ld_val & _GEN_1636 | stq_15_valid;
  wire        _GEN_2422 = dis_st_val_3 & _GEN_14 == 5'h10;
  wire        _GEN_2423 = ~dis_ld_val_3 & _GEN_2422 | ~dis_ld_val_2 & _GEN_2118 | ~dis_ld_val_1 & _GEN_2021 | ~dis_ld_val & _GEN_1637 | stq_16_valid;
  wire        _GEN_2424 = dis_st_val_3 & _GEN_14 == 5'h11;
  wire        _GEN_2425 = ~dis_ld_val_3 & _GEN_2424 | ~dis_ld_val_2 & _GEN_2119 | ~dis_ld_val_1 & _GEN_2022 | ~dis_ld_val & _GEN_1638 | stq_17_valid;
  wire        _GEN_2426 = dis_st_val_3 & _GEN_14 == 5'h12;
  wire        _GEN_2427 = ~dis_ld_val_3 & _GEN_2426 | ~dis_ld_val_2 & _GEN_2120 | ~dis_ld_val_1 & _GEN_2023 | ~dis_ld_val & _GEN_1639 | stq_18_valid;
  wire        _GEN_2428 = dis_st_val_3 & _GEN_14 == 5'h13;
  wire        _GEN_2429 = ~dis_ld_val_3 & _GEN_2428 | ~dis_ld_val_2 & _GEN_2121 | ~dis_ld_val_1 & _GEN_2024 | ~dis_ld_val & _GEN_1640 | stq_19_valid;
  wire        _GEN_2430 = dis_st_val_3 & _GEN_14 == 5'h14;
  wire        _GEN_2431 = ~dis_ld_val_3 & _GEN_2430 | ~dis_ld_val_2 & _GEN_2122 | ~dis_ld_val_1 & _GEN_2025 | ~dis_ld_val & _GEN_1641 | stq_20_valid;
  wire        _GEN_2432 = dis_st_val_3 & _GEN_14 == 5'h15;
  wire        _GEN_2433 = ~dis_ld_val_3 & _GEN_2432 | ~dis_ld_val_2 & _GEN_2123 | ~dis_ld_val_1 & _GEN_2026 | ~dis_ld_val & _GEN_1642 | stq_21_valid;
  wire        _GEN_2434 = dis_st_val_3 & _GEN_14 == 5'h16;
  wire        _GEN_2435 = ~dis_ld_val_3 & _GEN_2434 | ~dis_ld_val_2 & _GEN_2124 | ~dis_ld_val_1 & _GEN_2027 | ~dis_ld_val & _GEN_1643 | stq_22_valid;
  wire        _GEN_2436 = dis_st_val_3 & _GEN_14 == 5'h17;
  wire        _GEN_2437 = ~dis_ld_val_3 & _GEN_2436 | ~dis_ld_val_2 & _GEN_2125 | ~dis_ld_val_1 & _GEN_2028 | ~dis_ld_val & _GEN_1644 | stq_23_valid;
  wire        _GEN_2438 = dis_st_val_3 & _GEN_14 == 5'h18;
  wire        _GEN_2439 = ~dis_ld_val_3 & _GEN_2438 | ~dis_ld_val_2 & _GEN_2126 | ~dis_ld_val_1 & _GEN_2029 | ~dis_ld_val & _GEN_1645 | stq_24_valid;
  wire        _GEN_2440 = dis_st_val_3 & _GEN_14 == 5'h19;
  wire        _GEN_2441 = ~dis_ld_val_3 & _GEN_2440 | ~dis_ld_val_2 & _GEN_2127 | ~dis_ld_val_1 & _GEN_2030 | ~dis_ld_val & _GEN_1646 | stq_25_valid;
  wire        _GEN_2442 = dis_st_val_3 & _GEN_14 == 5'h1A;
  wire        _GEN_2443 = ~dis_ld_val_3 & _GEN_2442 | ~dis_ld_val_2 & _GEN_2128 | ~dis_ld_val_1 & _GEN_2031 | ~dis_ld_val & _GEN_1647 | stq_26_valid;
  wire        _GEN_2444 = dis_st_val_3 & _GEN_14 == 5'h1B;
  wire        _GEN_2445 = ~dis_ld_val_3 & _GEN_2444 | ~dis_ld_val_2 & _GEN_2129 | ~dis_ld_val_1 & _GEN_2032 | ~dis_ld_val & _GEN_1648 | stq_27_valid;
  wire        _GEN_2446 = dis_st_val_3 & _GEN_14 == 5'h1C;
  wire        _GEN_2447 = ~dis_ld_val_3 & _GEN_2446 | ~dis_ld_val_2 & _GEN_2130 | ~dis_ld_val_1 & _GEN_2033 | ~dis_ld_val & _GEN_1649 | stq_28_valid;
  wire        _GEN_2448 = dis_st_val_3 & _GEN_14 == 5'h1D;
  wire        _GEN_2449 = ~dis_ld_val_3 & _GEN_2448 | ~dis_ld_val_2 & _GEN_2131 | ~dis_ld_val_1 & _GEN_2034 | ~dis_ld_val & _GEN_1650 | stq_29_valid;
  wire        _GEN_2450 = dis_st_val_3 & _GEN_14 == 5'h1E;
  wire        _GEN_2451 = ~dis_ld_val_3 & _GEN_2450 | ~dis_ld_val_2 & _GEN_2132 | ~dis_ld_val_1 & _GEN_2035 | ~dis_ld_val & _GEN_1651 | stq_30_valid;
  wire        _GEN_2452 = dis_st_val_3 & (&_GEN_14);
  wire        _GEN_2453 = ~dis_ld_val_3 & _GEN_2452 | ~dis_ld_val_2 & _GEN_2133 | ~dis_ld_val_1 & _GEN_2036 | ~dis_ld_val & _GEN_1652 | stq_31_valid;
  wire        _GEN_2454 = dis_ld_val_3 | ~_GEN_2390;
  wire        _GEN_2455 = dis_ld_val_3 | ~_GEN_2392;
  wire        _GEN_2456 = dis_ld_val_3 | ~_GEN_2394;
  wire        _GEN_2457 = dis_ld_val_3 | ~_GEN_2396;
  wire        _GEN_2458 = dis_ld_val_3 | ~_GEN_2398;
  wire        _GEN_2459 = dis_ld_val_3 | ~_GEN_2400;
  wire        _GEN_2460 = dis_ld_val_3 | ~_GEN_2402;
  wire        _GEN_2461 = dis_ld_val_3 | ~_GEN_2404;
  wire        _GEN_2462 = dis_ld_val_3 | ~_GEN_2406;
  wire        _GEN_2463 = dis_ld_val_3 | ~_GEN_2408;
  wire        _GEN_2464 = dis_ld_val_3 | ~_GEN_2410;
  wire        _GEN_2465 = dis_ld_val_3 | ~_GEN_2412;
  wire        _GEN_2466 = dis_ld_val_3 | ~_GEN_2414;
  wire        _GEN_2467 = dis_ld_val_3 | ~_GEN_2416;
  wire        _GEN_2468 = dis_ld_val_3 | ~_GEN_2418;
  wire        _GEN_2469 = dis_ld_val_3 | ~_GEN_2420;
  wire        _GEN_2470 = dis_ld_val_3 | ~_GEN_2422;
  wire        _GEN_2471 = dis_ld_val_3 | ~_GEN_2424;
  wire        _GEN_2472 = dis_ld_val_3 | ~_GEN_2426;
  wire        _GEN_2473 = dis_ld_val_3 | ~_GEN_2428;
  wire        _GEN_2474 = dis_ld_val_3 | ~_GEN_2430;
  wire        _GEN_2475 = dis_ld_val_3 | ~_GEN_2432;
  wire        _GEN_2476 = dis_ld_val_3 | ~_GEN_2434;
  wire        _GEN_2477 = dis_ld_val_3 | ~_GEN_2436;
  wire        _GEN_2478 = dis_ld_val_3 | ~_GEN_2438;
  wire        _GEN_2479 = dis_ld_val_3 | ~_GEN_2440;
  wire        _GEN_2480 = dis_ld_val_3 | ~_GEN_2442;
  wire        _GEN_2481 = dis_ld_val_3 | ~_GEN_2444;
  wire        _GEN_2482 = dis_ld_val_3 | ~_GEN_2446;
  wire        _GEN_2483 = dis_ld_val_3 | ~_GEN_2448;
  wire        _GEN_2484 = dis_ld_val_3 | ~_GEN_2450;
  wire        _GEN_2485 = dis_ld_val_3 | ~_GEN_2452;
  wire        _GEN_2486 = _GEN_2454 & _GEN_2134 & _GEN_2037 & _GEN_1653 & stq_0_bits_data_valid;
  wire        _GEN_2487 = _GEN_2455 & _GEN_2135 & _GEN_2038 & _GEN_1654 & stq_1_bits_data_valid;
  wire        _GEN_2488 = _GEN_2456 & _GEN_2136 & _GEN_2039 & _GEN_1655 & stq_2_bits_data_valid;
  wire        _GEN_2489 = _GEN_2457 & _GEN_2137 & _GEN_2040 & _GEN_1656 & stq_3_bits_data_valid;
  wire        _GEN_2490 = _GEN_2458 & _GEN_2138 & _GEN_2041 & _GEN_1657 & stq_4_bits_data_valid;
  wire        _GEN_2491 = _GEN_2459 & _GEN_2139 & _GEN_2042 & _GEN_1658 & stq_5_bits_data_valid;
  wire        _GEN_2492 = _GEN_2460 & _GEN_2140 & _GEN_2043 & _GEN_1659 & stq_6_bits_data_valid;
  wire        _GEN_2493 = _GEN_2461 & _GEN_2141 & _GEN_2044 & _GEN_1660 & stq_7_bits_data_valid;
  wire        _GEN_2494 = _GEN_2462 & _GEN_2142 & _GEN_2045 & _GEN_1661 & stq_8_bits_data_valid;
  wire        _GEN_2495 = _GEN_2463 & _GEN_2143 & _GEN_2046 & _GEN_1662 & stq_9_bits_data_valid;
  wire        _GEN_2496 = _GEN_2464 & _GEN_2144 & _GEN_2047 & _GEN_1663 & stq_10_bits_data_valid;
  wire        _GEN_2497 = _GEN_2465 & _GEN_2145 & _GEN_2048 & _GEN_1664 & stq_11_bits_data_valid;
  wire        _GEN_2498 = _GEN_2466 & _GEN_2146 & _GEN_2049 & _GEN_1665 & stq_12_bits_data_valid;
  wire        _GEN_2499 = _GEN_2467 & _GEN_2147 & _GEN_2050 & _GEN_1666 & stq_13_bits_data_valid;
  wire        _GEN_2500 = _GEN_2468 & _GEN_2148 & _GEN_2051 & _GEN_1667 & stq_14_bits_data_valid;
  wire        _GEN_2501 = _GEN_2469 & _GEN_2149 & _GEN_2052 & _GEN_1668 & stq_15_bits_data_valid;
  wire        _GEN_2502 = _GEN_2470 & _GEN_2150 & _GEN_2053 & _GEN_1669 & stq_16_bits_data_valid;
  wire        _GEN_2503 = _GEN_2471 & _GEN_2151 & _GEN_2054 & _GEN_1670 & stq_17_bits_data_valid;
  wire        _GEN_2504 = _GEN_2472 & _GEN_2152 & _GEN_2055 & _GEN_1671 & stq_18_bits_data_valid;
  wire        _GEN_2505 = _GEN_2473 & _GEN_2153 & _GEN_2056 & _GEN_1672 & stq_19_bits_data_valid;
  wire        _GEN_2506 = _GEN_2474 & _GEN_2154 & _GEN_2057 & _GEN_1673 & stq_20_bits_data_valid;
  wire        _GEN_2507 = _GEN_2475 & _GEN_2155 & _GEN_2058 & _GEN_1674 & stq_21_bits_data_valid;
  wire        _GEN_2508 = _GEN_2476 & _GEN_2156 & _GEN_2059 & _GEN_1675 & stq_22_bits_data_valid;
  wire        _GEN_2509 = _GEN_2477 & _GEN_2157 & _GEN_2060 & _GEN_1676 & stq_23_bits_data_valid;
  wire        _GEN_2510 = _GEN_2478 & _GEN_2158 & _GEN_2061 & _GEN_1677 & stq_24_bits_data_valid;
  wire        _GEN_2511 = _GEN_2479 & _GEN_2159 & _GEN_2062 & _GEN_1678 & stq_25_bits_data_valid;
  wire        _GEN_2512 = _GEN_2480 & _GEN_2160 & _GEN_2063 & _GEN_1679 & stq_26_bits_data_valid;
  wire        _GEN_2513 = _GEN_2481 & _GEN_2161 & _GEN_2064 & _GEN_1680 & stq_27_bits_data_valid;
  wire        _GEN_2514 = _GEN_2482 & _GEN_2162 & _GEN_2065 & _GEN_1681 & stq_28_bits_data_valid;
  wire        _GEN_2515 = _GEN_2483 & _GEN_2163 & _GEN_2066 & _GEN_1682 & stq_29_bits_data_valid;
  wire        _GEN_2516 = _GEN_2484 & _GEN_2164 & _GEN_2067 & _GEN_1683 & stq_30_bits_data_valid;
  wire        _GEN_2517 = _GEN_2485 & _GEN_2165 & _GEN_2068 & _GEN_1684 & stq_31_bits_data_valid;
  wire        _GEN_2518 = _GEN_2454 & _GEN_2134 & _GEN_2037 & _GEN_1653 & stq_0_bits_committed;
  wire        _GEN_2519 = _GEN_2455 & _GEN_2135 & _GEN_2038 & _GEN_1654 & stq_1_bits_committed;
  wire        _GEN_2520 = _GEN_2456 & _GEN_2136 & _GEN_2039 & _GEN_1655 & stq_2_bits_committed;
  wire        _GEN_2521 = _GEN_2457 & _GEN_2137 & _GEN_2040 & _GEN_1656 & stq_3_bits_committed;
  wire        _GEN_2522 = _GEN_2458 & _GEN_2138 & _GEN_2041 & _GEN_1657 & stq_4_bits_committed;
  wire        _GEN_2523 = _GEN_2459 & _GEN_2139 & _GEN_2042 & _GEN_1658 & stq_5_bits_committed;
  wire        _GEN_2524 = _GEN_2460 & _GEN_2140 & _GEN_2043 & _GEN_1659 & stq_6_bits_committed;
  wire        _GEN_2525 = _GEN_2461 & _GEN_2141 & _GEN_2044 & _GEN_1660 & stq_7_bits_committed;
  wire        _GEN_2526 = _GEN_2462 & _GEN_2142 & _GEN_2045 & _GEN_1661 & stq_8_bits_committed;
  wire        _GEN_2527 = _GEN_2463 & _GEN_2143 & _GEN_2046 & _GEN_1662 & stq_9_bits_committed;
  wire        _GEN_2528 = _GEN_2464 & _GEN_2144 & _GEN_2047 & _GEN_1663 & stq_10_bits_committed;
  wire        _GEN_2529 = _GEN_2465 & _GEN_2145 & _GEN_2048 & _GEN_1664 & stq_11_bits_committed;
  wire        _GEN_2530 = _GEN_2466 & _GEN_2146 & _GEN_2049 & _GEN_1665 & stq_12_bits_committed;
  wire        _GEN_2531 = _GEN_2467 & _GEN_2147 & _GEN_2050 & _GEN_1666 & stq_13_bits_committed;
  wire        _GEN_2532 = _GEN_2468 & _GEN_2148 & _GEN_2051 & _GEN_1667 & stq_14_bits_committed;
  wire        _GEN_2533 = _GEN_2469 & _GEN_2149 & _GEN_2052 & _GEN_1668 & stq_15_bits_committed;
  wire        _GEN_2534 = _GEN_2470 & _GEN_2150 & _GEN_2053 & _GEN_1669 & stq_16_bits_committed;
  wire        _GEN_2535 = _GEN_2471 & _GEN_2151 & _GEN_2054 & _GEN_1670 & stq_17_bits_committed;
  wire        _GEN_2536 = _GEN_2472 & _GEN_2152 & _GEN_2055 & _GEN_1671 & stq_18_bits_committed;
  wire        _GEN_2537 = _GEN_2473 & _GEN_2153 & _GEN_2056 & _GEN_1672 & stq_19_bits_committed;
  wire        _GEN_2538 = _GEN_2474 & _GEN_2154 & _GEN_2057 & _GEN_1673 & stq_20_bits_committed;
  wire        _GEN_2539 = _GEN_2475 & _GEN_2155 & _GEN_2058 & _GEN_1674 & stq_21_bits_committed;
  wire        _GEN_2540 = _GEN_2476 & _GEN_2156 & _GEN_2059 & _GEN_1675 & stq_22_bits_committed;
  wire        _GEN_2541 = _GEN_2477 & _GEN_2157 & _GEN_2060 & _GEN_1676 & stq_23_bits_committed;
  wire        _GEN_2542 = _GEN_2478 & _GEN_2158 & _GEN_2061 & _GEN_1677 & stq_24_bits_committed;
  wire        _GEN_2543 = _GEN_2479 & _GEN_2159 & _GEN_2062 & _GEN_1678 & stq_25_bits_committed;
  wire        _GEN_2544 = _GEN_2480 & _GEN_2160 & _GEN_2063 & _GEN_1679 & stq_26_bits_committed;
  wire        _GEN_2545 = _GEN_2481 & _GEN_2161 & _GEN_2064 & _GEN_1680 & stq_27_bits_committed;
  wire        _GEN_2546 = _GEN_2482 & _GEN_2162 & _GEN_2065 & _GEN_1681 & stq_28_bits_committed;
  wire        _GEN_2547 = _GEN_2483 & _GEN_2163 & _GEN_2066 & _GEN_1682 & stq_29_bits_committed;
  wire        _GEN_2548 = _GEN_2484 & _GEN_2164 & _GEN_2067 & _GEN_1683 & stq_30_bits_committed;
  wire        _GEN_2549 = _GEN_2485 & _GEN_2165 & _GEN_2068 & _GEN_1684 & stq_31_bits_committed;
  wire        ldq_retry_idx_block = (will_fire_load_wakeup_1_will_fire ? _GEN_145 : will_fire_load_incoming_1_will_fire ? _GEN_178 : _GEN_240) | p1_block_load_mask_0;
  wire        _ldq_retry_idx_T_2 = ldq_0_bits_addr_valid & ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;
  wire        ldq_retry_idx_block_1 = (will_fire_load_wakeup_1_will_fire ? _GEN_146 : will_fire_load_incoming_1_will_fire ? _GEN_180 : _GEN_241) | p1_block_load_mask_1;
  wire        _ldq_retry_idx_T_5 = ldq_1_bits_addr_valid & ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;
  wire        ldq_retry_idx_block_2 = (will_fire_load_wakeup_1_will_fire ? _GEN_147 : will_fire_load_incoming_1_will_fire ? _GEN_182 : _GEN_242) | p1_block_load_mask_2;
  wire        _ldq_retry_idx_T_8 = ldq_2_bits_addr_valid & ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;
  wire        ldq_retry_idx_block_3 = (will_fire_load_wakeup_1_will_fire ? _GEN_148 : will_fire_load_incoming_1_will_fire ? _GEN_184 : _GEN_243) | p1_block_load_mask_3;
  wire        _ldq_retry_idx_T_11 = ldq_3_bits_addr_valid & ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;
  wire        ldq_retry_idx_block_4 = (will_fire_load_wakeup_1_will_fire ? _GEN_149 : will_fire_load_incoming_1_will_fire ? _GEN_186 : _GEN_244) | p1_block_load_mask_4;
  wire        _ldq_retry_idx_T_14 = ldq_4_bits_addr_valid & ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;
  wire        ldq_retry_idx_block_5 = (will_fire_load_wakeup_1_will_fire ? _GEN_150 : will_fire_load_incoming_1_will_fire ? _GEN_188 : _GEN_245) | p1_block_load_mask_5;
  wire        _ldq_retry_idx_T_17 = ldq_5_bits_addr_valid & ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;
  wire        ldq_retry_idx_block_6 = (will_fire_load_wakeup_1_will_fire ? _GEN_151 : will_fire_load_incoming_1_will_fire ? _GEN_190 : _GEN_246) | p1_block_load_mask_6;
  wire        _ldq_retry_idx_T_20 = ldq_6_bits_addr_valid & ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;
  wire        ldq_retry_idx_block_7 = (will_fire_load_wakeup_1_will_fire ? _GEN_152 : will_fire_load_incoming_1_will_fire ? _GEN_192 : _GEN_247) | p1_block_load_mask_7;
  wire        _ldq_retry_idx_T_23 = ldq_7_bits_addr_valid & ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;
  wire        ldq_retry_idx_block_8 = (will_fire_load_wakeup_1_will_fire ? _GEN_153 : will_fire_load_incoming_1_will_fire ? _GEN_194 : _GEN_248) | p1_block_load_mask_8;
  wire        _ldq_retry_idx_T_26 = ldq_8_bits_addr_valid & ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;
  wire        ldq_retry_idx_block_9 = (will_fire_load_wakeup_1_will_fire ? _GEN_154 : will_fire_load_incoming_1_will_fire ? _GEN_196 : _GEN_249) | p1_block_load_mask_9;
  wire        _ldq_retry_idx_T_29 = ldq_9_bits_addr_valid & ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;
  wire        ldq_retry_idx_block_10 = (will_fire_load_wakeup_1_will_fire ? _GEN_155 : will_fire_load_incoming_1_will_fire ? _GEN_198 : _GEN_250) | p1_block_load_mask_10;
  wire        _ldq_retry_idx_T_32 = ldq_10_bits_addr_valid & ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;
  wire        ldq_retry_idx_block_11 = (will_fire_load_wakeup_1_will_fire ? _GEN_156 : will_fire_load_incoming_1_will_fire ? _GEN_200 : _GEN_251) | p1_block_load_mask_11;
  wire        _ldq_retry_idx_T_35 = ldq_11_bits_addr_valid & ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;
  wire        ldq_retry_idx_block_12 = (will_fire_load_wakeup_1_will_fire ? _GEN_157 : will_fire_load_incoming_1_will_fire ? _GEN_202 : _GEN_252) | p1_block_load_mask_12;
  wire        _ldq_retry_idx_T_38 = ldq_12_bits_addr_valid & ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;
  wire        ldq_retry_idx_block_13 = (will_fire_load_wakeup_1_will_fire ? _GEN_158 : will_fire_load_incoming_1_will_fire ? _GEN_204 : _GEN_253) | p1_block_load_mask_13;
  wire        _ldq_retry_idx_T_41 = ldq_13_bits_addr_valid & ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;
  wire        ldq_retry_idx_block_14 = (will_fire_load_wakeup_1_will_fire ? _GEN_159 : will_fire_load_incoming_1_will_fire ? _GEN_206 : _GEN_254) | p1_block_load_mask_14;
  wire        _ldq_retry_idx_T_44 = ldq_14_bits_addr_valid & ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;
  wire        ldq_retry_idx_block_15 = (will_fire_load_wakeup_1_will_fire ? _GEN_160 : will_fire_load_incoming_1_will_fire ? _GEN_208 : _GEN_255) | p1_block_load_mask_15;
  wire        _ldq_retry_idx_T_47 = ldq_15_bits_addr_valid & ldq_15_bits_addr_is_virtual & ~ldq_retry_idx_block_15;
  wire        ldq_retry_idx_block_16 = (will_fire_load_wakeup_1_will_fire ? _GEN_161 : will_fire_load_incoming_1_will_fire ? _GEN_210 : _GEN_256) | p1_block_load_mask_16;
  wire        _ldq_retry_idx_T_50 = ldq_16_bits_addr_valid & ldq_16_bits_addr_is_virtual & ~ldq_retry_idx_block_16;
  wire        ldq_retry_idx_block_17 = (will_fire_load_wakeup_1_will_fire ? _GEN_162 : will_fire_load_incoming_1_will_fire ? _GEN_212 : _GEN_257) | p1_block_load_mask_17;
  wire        _ldq_retry_idx_T_53 = ldq_17_bits_addr_valid & ldq_17_bits_addr_is_virtual & ~ldq_retry_idx_block_17;
  wire        ldq_retry_idx_block_18 = (will_fire_load_wakeup_1_will_fire ? _GEN_163 : will_fire_load_incoming_1_will_fire ? _GEN_214 : _GEN_258) | p1_block_load_mask_18;
  wire        _ldq_retry_idx_T_56 = ldq_18_bits_addr_valid & ldq_18_bits_addr_is_virtual & ~ldq_retry_idx_block_18;
  wire        ldq_retry_idx_block_19 = (will_fire_load_wakeup_1_will_fire ? _GEN_164 : will_fire_load_incoming_1_will_fire ? _GEN_216 : _GEN_259) | p1_block_load_mask_19;
  wire        _ldq_retry_idx_T_59 = ldq_19_bits_addr_valid & ldq_19_bits_addr_is_virtual & ~ldq_retry_idx_block_19;
  wire        ldq_retry_idx_block_20 = (will_fire_load_wakeup_1_will_fire ? _GEN_165 : will_fire_load_incoming_1_will_fire ? _GEN_218 : _GEN_260) | p1_block_load_mask_20;
  wire        _ldq_retry_idx_T_62 = ldq_20_bits_addr_valid & ldq_20_bits_addr_is_virtual & ~ldq_retry_idx_block_20;
  wire        ldq_retry_idx_block_21 = (will_fire_load_wakeup_1_will_fire ? _GEN_166 : will_fire_load_incoming_1_will_fire ? _GEN_220 : _GEN_261) | p1_block_load_mask_21;
  wire        _ldq_retry_idx_T_65 = ldq_21_bits_addr_valid & ldq_21_bits_addr_is_virtual & ~ldq_retry_idx_block_21;
  wire        ldq_retry_idx_block_22 = (will_fire_load_wakeup_1_will_fire ? _GEN_167 : will_fire_load_incoming_1_will_fire ? _GEN_222 : _GEN_262) | p1_block_load_mask_22;
  wire        _ldq_retry_idx_T_68 = ldq_22_bits_addr_valid & ldq_22_bits_addr_is_virtual & ~ldq_retry_idx_block_22;
  wire        ldq_retry_idx_block_23 = (will_fire_load_wakeup_1_will_fire ? _GEN_168 : will_fire_load_incoming_1_will_fire ? _GEN_224 : _GEN_263) | p1_block_load_mask_23;
  wire        _ldq_retry_idx_T_71 = ldq_23_bits_addr_valid & ldq_23_bits_addr_is_virtual & ~ldq_retry_idx_block_23;
  wire        ldq_retry_idx_block_24 = (will_fire_load_wakeup_1_will_fire ? _GEN_169 : will_fire_load_incoming_1_will_fire ? _GEN_226 : _GEN_264) | p1_block_load_mask_24;
  wire        _ldq_retry_idx_T_74 = ldq_24_bits_addr_valid & ldq_24_bits_addr_is_virtual & ~ldq_retry_idx_block_24;
  wire        ldq_retry_idx_block_25 = (will_fire_load_wakeup_1_will_fire ? _GEN_170 : will_fire_load_incoming_1_will_fire ? _GEN_228 : _GEN_265) | p1_block_load_mask_25;
  wire        _ldq_retry_idx_T_77 = ldq_25_bits_addr_valid & ldq_25_bits_addr_is_virtual & ~ldq_retry_idx_block_25;
  wire        ldq_retry_idx_block_26 = (will_fire_load_wakeup_1_will_fire ? _GEN_171 : will_fire_load_incoming_1_will_fire ? _GEN_230 : _GEN_266) | p1_block_load_mask_26;
  wire        _ldq_retry_idx_T_80 = ldq_26_bits_addr_valid & ldq_26_bits_addr_is_virtual & ~ldq_retry_idx_block_26;
  wire        ldq_retry_idx_block_27 = (will_fire_load_wakeup_1_will_fire ? _GEN_172 : will_fire_load_incoming_1_will_fire ? _GEN_232 : _GEN_267) | p1_block_load_mask_27;
  wire        _ldq_retry_idx_T_83 = ldq_27_bits_addr_valid & ldq_27_bits_addr_is_virtual & ~ldq_retry_idx_block_27;
  wire        ldq_retry_idx_block_28 = (will_fire_load_wakeup_1_will_fire ? _GEN_173 : will_fire_load_incoming_1_will_fire ? _GEN_234 : _GEN_268) | p1_block_load_mask_28;
  wire        _ldq_retry_idx_T_86 = ldq_28_bits_addr_valid & ldq_28_bits_addr_is_virtual & ~ldq_retry_idx_block_28;
  wire        ldq_retry_idx_block_29 = (will_fire_load_wakeup_1_will_fire ? _GEN_174 : will_fire_load_incoming_1_will_fire ? _GEN_236 : _GEN_269) | p1_block_load_mask_29;
  wire        _ldq_retry_idx_T_89 = ldq_29_bits_addr_valid & ldq_29_bits_addr_is_virtual & ~ldq_retry_idx_block_29;
  wire        ldq_retry_idx_block_30 = (will_fire_load_wakeup_1_will_fire ? _GEN_175 : will_fire_load_incoming_1_will_fire ? _GEN_238 : _GEN_270) | p1_block_load_mask_30;
  wire        _ldq_retry_idx_T_92 = ldq_30_bits_addr_valid & ldq_30_bits_addr_is_virtual & ~ldq_retry_idx_block_30;
  wire        ldq_retry_idx_block_31 = (will_fire_load_wakeup_1_will_fire ? _GEN_176 : will_fire_load_incoming_1_will_fire ? _GEN_239 : _GEN_271) | p1_block_load_mask_31;
  wire        _stq_retry_idx_T = stq_0_bits_addr_valid & stq_0_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_1 = stq_1_bits_addr_valid & stq_1_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_2 = stq_2_bits_addr_valid & stq_2_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_3 = stq_3_bits_addr_valid & stq_3_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_4 = stq_4_bits_addr_valid & stq_4_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_5 = stq_5_bits_addr_valid & stq_5_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_6 = stq_6_bits_addr_valid & stq_6_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_7 = stq_7_bits_addr_valid & stq_7_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_8 = stq_8_bits_addr_valid & stq_8_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_9 = stq_9_bits_addr_valid & stq_9_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_10 = stq_10_bits_addr_valid & stq_10_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_11 = stq_11_bits_addr_valid & stq_11_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_12 = stq_12_bits_addr_valid & stq_12_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_13 = stq_13_bits_addr_valid & stq_13_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_14 = stq_14_bits_addr_valid & stq_14_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_15 = stq_15_bits_addr_valid & stq_15_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_16 = stq_16_bits_addr_valid & stq_16_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_17 = stq_17_bits_addr_valid & stq_17_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_18 = stq_18_bits_addr_valid & stq_18_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_19 = stq_19_bits_addr_valid & stq_19_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_20 = stq_20_bits_addr_valid & stq_20_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_21 = stq_21_bits_addr_valid & stq_21_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_22 = stq_22_bits_addr_valid & stq_22_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_23 = stq_23_bits_addr_valid & stq_23_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_24 = stq_24_bits_addr_valid & stq_24_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_25 = stq_25_bits_addr_valid & stq_25_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_26 = stq_26_bits_addr_valid & stq_26_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_27 = stq_27_bits_addr_valid & stq_27_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_28 = stq_28_bits_addr_valid & stq_28_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_29 = stq_29_bits_addr_valid & stq_29_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_30 = stq_30_bits_addr_valid & stq_30_bits_addr_is_virtual;
  wire        _ldq_wakeup_idx_T_7 = ldq_0_bits_addr_valid & ~ldq_0_bits_executed & ~ldq_0_bits_succeeded & ~ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;
  wire        _ldq_wakeup_idx_T_15 = ldq_1_bits_addr_valid & ~ldq_1_bits_executed & ~ldq_1_bits_succeeded & ~ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;
  wire        _ldq_wakeup_idx_T_23 = ldq_2_bits_addr_valid & ~ldq_2_bits_executed & ~ldq_2_bits_succeeded & ~ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;
  wire        _ldq_wakeup_idx_T_31 = ldq_3_bits_addr_valid & ~ldq_3_bits_executed & ~ldq_3_bits_succeeded & ~ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;
  wire        _ldq_wakeup_idx_T_39 = ldq_4_bits_addr_valid & ~ldq_4_bits_executed & ~ldq_4_bits_succeeded & ~ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;
  wire        _ldq_wakeup_idx_T_47 = ldq_5_bits_addr_valid & ~ldq_5_bits_executed & ~ldq_5_bits_succeeded & ~ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;
  wire        _ldq_wakeup_idx_T_55 = ldq_6_bits_addr_valid & ~ldq_6_bits_executed & ~ldq_6_bits_succeeded & ~ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;
  wire        _ldq_wakeup_idx_T_63 = ldq_7_bits_addr_valid & ~ldq_7_bits_executed & ~ldq_7_bits_succeeded & ~ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;
  wire        _ldq_wakeup_idx_T_71 = ldq_8_bits_addr_valid & ~ldq_8_bits_executed & ~ldq_8_bits_succeeded & ~ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;
  wire        _ldq_wakeup_idx_T_79 = ldq_9_bits_addr_valid & ~ldq_9_bits_executed & ~ldq_9_bits_succeeded & ~ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;
  wire        _ldq_wakeup_idx_T_87 = ldq_10_bits_addr_valid & ~ldq_10_bits_executed & ~ldq_10_bits_succeeded & ~ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;
  wire        _ldq_wakeup_idx_T_95 = ldq_11_bits_addr_valid & ~ldq_11_bits_executed & ~ldq_11_bits_succeeded & ~ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;
  wire        _ldq_wakeup_idx_T_103 = ldq_12_bits_addr_valid & ~ldq_12_bits_executed & ~ldq_12_bits_succeeded & ~ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;
  wire        _ldq_wakeup_idx_T_111 = ldq_13_bits_addr_valid & ~ldq_13_bits_executed & ~ldq_13_bits_succeeded & ~ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;
  wire        _ldq_wakeup_idx_T_119 = ldq_14_bits_addr_valid & ~ldq_14_bits_executed & ~ldq_14_bits_succeeded & ~ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;
  wire        _ldq_wakeup_idx_T_127 = ldq_15_bits_addr_valid & ~ldq_15_bits_executed & ~ldq_15_bits_succeeded & ~ldq_15_bits_addr_is_virtual & ~ldq_retry_idx_block_15;
  wire        _ldq_wakeup_idx_T_135 = ldq_16_bits_addr_valid & ~ldq_16_bits_executed & ~ldq_16_bits_succeeded & ~ldq_16_bits_addr_is_virtual & ~ldq_retry_idx_block_16;
  wire        _ldq_wakeup_idx_T_143 = ldq_17_bits_addr_valid & ~ldq_17_bits_executed & ~ldq_17_bits_succeeded & ~ldq_17_bits_addr_is_virtual & ~ldq_retry_idx_block_17;
  wire        _ldq_wakeup_idx_T_151 = ldq_18_bits_addr_valid & ~ldq_18_bits_executed & ~ldq_18_bits_succeeded & ~ldq_18_bits_addr_is_virtual & ~ldq_retry_idx_block_18;
  wire        _ldq_wakeup_idx_T_159 = ldq_19_bits_addr_valid & ~ldq_19_bits_executed & ~ldq_19_bits_succeeded & ~ldq_19_bits_addr_is_virtual & ~ldq_retry_idx_block_19;
  wire        _ldq_wakeup_idx_T_167 = ldq_20_bits_addr_valid & ~ldq_20_bits_executed & ~ldq_20_bits_succeeded & ~ldq_20_bits_addr_is_virtual & ~ldq_retry_idx_block_20;
  wire        _ldq_wakeup_idx_T_175 = ldq_21_bits_addr_valid & ~ldq_21_bits_executed & ~ldq_21_bits_succeeded & ~ldq_21_bits_addr_is_virtual & ~ldq_retry_idx_block_21;
  wire        _ldq_wakeup_idx_T_183 = ldq_22_bits_addr_valid & ~ldq_22_bits_executed & ~ldq_22_bits_succeeded & ~ldq_22_bits_addr_is_virtual & ~ldq_retry_idx_block_22;
  wire        _ldq_wakeup_idx_T_191 = ldq_23_bits_addr_valid & ~ldq_23_bits_executed & ~ldq_23_bits_succeeded & ~ldq_23_bits_addr_is_virtual & ~ldq_retry_idx_block_23;
  wire        _ldq_wakeup_idx_T_199 = ldq_24_bits_addr_valid & ~ldq_24_bits_executed & ~ldq_24_bits_succeeded & ~ldq_24_bits_addr_is_virtual & ~ldq_retry_idx_block_24;
  wire        _ldq_wakeup_idx_T_207 = ldq_25_bits_addr_valid & ~ldq_25_bits_executed & ~ldq_25_bits_succeeded & ~ldq_25_bits_addr_is_virtual & ~ldq_retry_idx_block_25;
  wire        _ldq_wakeup_idx_T_215 = ldq_26_bits_addr_valid & ~ldq_26_bits_executed & ~ldq_26_bits_succeeded & ~ldq_26_bits_addr_is_virtual & ~ldq_retry_idx_block_26;
  wire        _ldq_wakeup_idx_T_223 = ldq_27_bits_addr_valid & ~ldq_27_bits_executed & ~ldq_27_bits_succeeded & ~ldq_27_bits_addr_is_virtual & ~ldq_retry_idx_block_27;
  wire        _ldq_wakeup_idx_T_231 = ldq_28_bits_addr_valid & ~ldq_28_bits_executed & ~ldq_28_bits_succeeded & ~ldq_28_bits_addr_is_virtual & ~ldq_retry_idx_block_28;
  wire        _ldq_wakeup_idx_T_239 = ldq_29_bits_addr_valid & ~ldq_29_bits_executed & ~ldq_29_bits_succeeded & ~ldq_29_bits_addr_is_virtual & ~ldq_retry_idx_block_29;
  wire        _ldq_wakeup_idx_T_247 = ldq_30_bits_addr_valid & ~ldq_30_bits_executed & ~ldq_30_bits_succeeded & ~ldq_30_bits_addr_is_virtual & ~ldq_retry_idx_block_30;
  wire        ma_ld_0 = will_fire_load_incoming_0_will_fire & exe_req_0_bits_mxcpt_valid;
  wire        ma_ld_1 = will_fire_load_incoming_1_will_fire & exe_req_1_bits_mxcpt_valid;
  wire        ma_st_0 = _stq_idx_T & exe_req_0_bits_mxcpt_valid;
  wire        ma_st_1 = _stq_idx_T_1 & exe_req_1_bits_mxcpt_valid;
  wire        pf_ld_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_ld & _mem_xcpt_uops_WIRE_0_uses_ldq;
  wire        pf_ld_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_pf_ld & _mem_xcpt_uops_WIRE_1_uses_ldq;
  wire        pf_st_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_st & _mem_xcpt_uops_WIRE_0_uses_stq;
  wire        pf_st_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_pf_st & _mem_xcpt_uops_WIRE_1_uses_stq;
  wire        ae_ld_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_ae_ld & _mem_xcpt_uops_WIRE_0_uses_ldq;
  wire        ae_ld_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_ae_ld & _mem_xcpt_uops_WIRE_1_uses_ldq;
  wire        _GEN_2550 = mem_xcpt_valids_1 & (mem_xcpt_uops_1_rob_idx < mem_xcpt_uops_0_rob_idx ^ mem_xcpt_uops_1_rob_idx < io_core_rob_head_idx ^ mem_xcpt_uops_0_rob_idx < io_core_rob_head_idx | ~mem_xcpt_valids_0);
  wire [6:0]  mem_xcpt_uop_rob_idx = _GEN_2550 ? mem_xcpt_uops_1_rob_idx : mem_xcpt_uops_0_rob_idx;
  wire        _GEN_2551 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h0;
  wire        _GEN_2552 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h1;
  wire        _GEN_2553 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h2;
  wire        _GEN_2554 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h3;
  wire        _GEN_2555 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h4;
  wire        _GEN_2556 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h5;
  wire        _GEN_2557 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h6;
  wire        _GEN_2558 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h7;
  wire        _GEN_2559 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h8;
  wire        _GEN_2560 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h9;
  wire        _GEN_2561 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hA;
  wire        _GEN_2562 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hB;
  wire        _GEN_2563 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hC;
  wire        _GEN_2564 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hD;
  wire        _GEN_2565 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hE;
  wire        _GEN_2566 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'hF;
  wire        _GEN_2567 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h10;
  wire        _GEN_2568 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h11;
  wire        _GEN_2569 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h12;
  wire        _GEN_2570 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h13;
  wire        _GEN_2571 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h14;
  wire        _GEN_2572 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h15;
  wire        _GEN_2573 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h16;
  wire        _GEN_2574 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h17;
  wire        _GEN_2575 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h18;
  wire        _GEN_2576 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h19;
  wire        _GEN_2577 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h1A;
  wire        _GEN_2578 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h1B;
  wire        _GEN_2579 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h1C;
  wire        _GEN_2580 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h1D;
  wire        _GEN_2581 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_ldq_idx == 5'h1E;
  wire        _GEN_2582 = mem_xcpt_valids_0 & mem_xcpt_uops_0_uses_ldq & (&mem_xcpt_uops_0_ldq_idx);
  wire        dmem_req_fire_0 = dmem_req_0_valid & _dmem_req_fire_T_2;
  wire        _GEN_2583 = stq_execute_head == 5'h0;
  wire        _GEN_2584 = stq_execute_head == 5'h1;
  wire        _GEN_2585 = stq_execute_head == 5'h2;
  wire        _GEN_2586 = stq_execute_head == 5'h3;
  wire        _GEN_2587 = stq_execute_head == 5'h4;
  wire        _GEN_2588 = stq_execute_head == 5'h5;
  wire        _GEN_2589 = stq_execute_head == 5'h6;
  wire        _GEN_2590 = stq_execute_head == 5'h7;
  wire        _GEN_2591 = stq_execute_head == 5'h8;
  wire        _GEN_2592 = stq_execute_head == 5'h9;
  wire        _GEN_2593 = stq_execute_head == 5'hA;
  wire        _GEN_2594 = stq_execute_head == 5'hB;
  wire        _GEN_2595 = stq_execute_head == 5'hC;
  wire        _GEN_2596 = stq_execute_head == 5'hD;
  wire        _GEN_2597 = stq_execute_head == 5'hE;
  wire        _GEN_2598 = stq_execute_head == 5'hF;
  wire        _GEN_2599 = stq_execute_head == 5'h10;
  wire        _GEN_2600 = stq_execute_head == 5'h11;
  wire        _GEN_2601 = stq_execute_head == 5'h12;
  wire        _GEN_2602 = stq_execute_head == 5'h13;
  wire        _GEN_2603 = stq_execute_head == 5'h14;
  wire        _GEN_2604 = stq_execute_head == 5'h15;
  wire        _GEN_2605 = stq_execute_head == 5'h16;
  wire        _GEN_2606 = stq_execute_head == 5'h17;
  wire        _GEN_2607 = stq_execute_head == 5'h18;
  wire        _GEN_2608 = stq_execute_head == 5'h19;
  wire        _GEN_2609 = stq_execute_head == 5'h1A;
  wire        _GEN_2610 = stq_execute_head == 5'h1B;
  wire        _GEN_2611 = stq_execute_head == 5'h1C;
  wire        _GEN_2612 = stq_execute_head == 5'h1D;
  wire        _GEN_2613 = stq_execute_head == 5'h1E;
  wire        _GEN_2614 = will_fire_load_incoming_0_will_fire ? _GEN_50 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_81 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_19 & dmem_req_fire_0;
  wire        _GEN_2615 = will_fire_load_incoming_0_will_fire ? _GEN_51 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_83 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_20 & dmem_req_fire_0;
  wire        _GEN_2616 = will_fire_load_incoming_0_will_fire ? _GEN_52 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_85 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_21 & dmem_req_fire_0;
  wire        _GEN_2617 = will_fire_load_incoming_0_will_fire ? _GEN_53 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_87 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_22 & dmem_req_fire_0;
  wire        _GEN_2618 = will_fire_load_incoming_0_will_fire ? _GEN_54 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_89 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_23 & dmem_req_fire_0;
  wire        _GEN_2619 = will_fire_load_incoming_0_will_fire ? _GEN_55 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_91 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_24 & dmem_req_fire_0;
  wire        _GEN_2620 = will_fire_load_incoming_0_will_fire ? _GEN_56 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_93 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_25 & dmem_req_fire_0;
  wire        _GEN_2621 = will_fire_load_incoming_0_will_fire ? _GEN_57 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_95 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_26 & dmem_req_fire_0;
  wire        _GEN_2622 = will_fire_load_incoming_0_will_fire ? _GEN_58 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_97 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_27 & dmem_req_fire_0;
  wire        _GEN_2623 = will_fire_load_incoming_0_will_fire ? _GEN_59 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_99 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_28 & dmem_req_fire_0;
  wire        _GEN_2624 = will_fire_load_incoming_0_will_fire ? _GEN_60 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_101 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_29 & dmem_req_fire_0;
  wire        _GEN_2625 = will_fire_load_incoming_0_will_fire ? _GEN_61 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_103 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_30 & dmem_req_fire_0;
  wire        _GEN_2626 = will_fire_load_incoming_0_will_fire ? _GEN_62 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_105 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_31 & dmem_req_fire_0;
  wire        _GEN_2627 = will_fire_load_incoming_0_will_fire ? _GEN_63 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_107 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_32 & dmem_req_fire_0;
  wire        _GEN_2628 = will_fire_load_incoming_0_will_fire ? _GEN_64 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_109 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_33 & dmem_req_fire_0;
  wire        _GEN_2629 = will_fire_load_incoming_0_will_fire ? _GEN_65 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_111 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_34 & dmem_req_fire_0;
  wire        _GEN_2630 = will_fire_load_incoming_0_will_fire ? _GEN_66 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_113 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_35 & dmem_req_fire_0;
  wire        _GEN_2631 = will_fire_load_incoming_0_will_fire ? _GEN_67 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_115 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_36 & dmem_req_fire_0;
  wire        _GEN_2632 = will_fire_load_incoming_0_will_fire ? _GEN_68 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_117 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_37 & dmem_req_fire_0;
  wire        _GEN_2633 = will_fire_load_incoming_0_will_fire ? _GEN_69 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_119 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_38 & dmem_req_fire_0;
  wire        _GEN_2634 = will_fire_load_incoming_0_will_fire ? _GEN_70 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_121 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_39 & dmem_req_fire_0;
  wire        _GEN_2635 = will_fire_load_incoming_0_will_fire ? _GEN_71 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_123 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_40 & dmem_req_fire_0;
  wire        _GEN_2636 = will_fire_load_incoming_0_will_fire ? _GEN_72 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_125 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_41 & dmem_req_fire_0;
  wire        _GEN_2637 = will_fire_load_incoming_0_will_fire ? _GEN_73 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_127 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_42 & dmem_req_fire_0;
  wire        _GEN_2638 = will_fire_load_incoming_0_will_fire ? _GEN_74 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_129 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_43 & dmem_req_fire_0;
  wire        _GEN_2639 = will_fire_load_incoming_0_will_fire ? _GEN_75 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_131 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_44 & dmem_req_fire_0;
  wire        _GEN_2640 = will_fire_load_incoming_0_will_fire ? _GEN_76 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_133 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_45 & dmem_req_fire_0;
  wire        _GEN_2641 = will_fire_load_incoming_0_will_fire ? _GEN_77 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_135 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_46 & dmem_req_fire_0;
  wire        _GEN_2642 = will_fire_load_incoming_0_will_fire ? _GEN_78 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_137 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_47 & dmem_req_fire_0;
  wire        _GEN_2643 = will_fire_load_incoming_0_will_fire ? _GEN_79 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_139 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_48 & dmem_req_fire_0;
  wire        _GEN_2644 = will_fire_load_incoming_0_will_fire ? _GEN_80 & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? _GEN_141 & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & _GEN_49 & dmem_req_fire_0;
  wire        _GEN_2645 = will_fire_load_incoming_0_will_fire ? (&_mem_incoming_uop_WIRE_0_ldq_idx) & dmem_req_fire_0 : will_fire_load_retry_0_will_fire ? (&ldq_retry_idx) & dmem_req_fire_0 : ~will_fire_store_commit_0_will_fire & will_fire_load_wakeup_0_will_fire & (&ldq_wakeup_idx) & dmem_req_fire_0;
  wire [4:0]  ldq_idx = will_fire_load_incoming_0_will_fire ? _mem_incoming_uop_WIRE_0_ldq_idx : ldq_retry_idx;
  wire        _GEN_2646 = _GEN_275 & ldq_idx == 5'h0;
  wire        _GEN_2647 = _GEN_275 & ldq_idx == 5'h1;
  wire        _GEN_2648 = _GEN_275 & ldq_idx == 5'h2;
  wire        _GEN_2649 = _GEN_275 & ldq_idx == 5'h3;
  wire        _GEN_2650 = _GEN_275 & ldq_idx == 5'h4;
  wire        _GEN_2651 = _GEN_275 & ldq_idx == 5'h5;
  wire        _GEN_2652 = _GEN_275 & ldq_idx == 5'h6;
  wire        _GEN_2653 = _GEN_275 & ldq_idx == 5'h7;
  wire        _GEN_2654 = _GEN_275 & ldq_idx == 5'h8;
  wire        _GEN_2655 = _GEN_275 & ldq_idx == 5'h9;
  wire        _GEN_2656 = _GEN_275 & ldq_idx == 5'hA;
  wire        _GEN_2657 = _GEN_275 & ldq_idx == 5'hB;
  wire        _GEN_2658 = _GEN_275 & ldq_idx == 5'hC;
  wire        _GEN_2659 = _GEN_275 & ldq_idx == 5'hD;
  wire        _GEN_2660 = _GEN_275 & ldq_idx == 5'hE;
  wire        _GEN_2661 = _GEN_275 & ldq_idx == 5'hF;
  wire        _GEN_2662 = _GEN_275 & ldq_idx == 5'h10;
  wire        _GEN_2663 = _GEN_275 & ldq_idx == 5'h11;
  wire        _GEN_2664 = _GEN_275 & ldq_idx == 5'h12;
  wire        _GEN_2665 = _GEN_275 & ldq_idx == 5'h13;
  wire        _GEN_2666 = _GEN_275 & ldq_idx == 5'h14;
  wire        _GEN_2667 = _GEN_275 & ldq_idx == 5'h15;
  wire        _GEN_2668 = _GEN_275 & ldq_idx == 5'h16;
  wire        _GEN_2669 = _GEN_275 & ldq_idx == 5'h17;
  wire        _GEN_2670 = _GEN_275 & ldq_idx == 5'h18;
  wire        _GEN_2671 = _GEN_275 & ldq_idx == 5'h19;
  wire        _GEN_2672 = _GEN_275 & ldq_idx == 5'h1A;
  wire        _GEN_2673 = _GEN_275 & ldq_idx == 5'h1B;
  wire        _GEN_2674 = _GEN_275 & ldq_idx == 5'h1C;
  wire        _GEN_2675 = _GEN_275 & ldq_idx == 5'h1D;
  wire        _GEN_2676 = _GEN_275 & ldq_idx == 5'h1E;
  wire        _GEN_2677 = _GEN_275 & (&ldq_idx);
  wire        _ldq_bits_addr_is_uncacheable_T_1 = ~_dtlb_io_resp_0_cacheable & ~exe_tlb_miss_0;
  wire [4:0]  stq_idx = _stq_idx_T ? _mem_incoming_uop_WIRE_0_stq_idx : stq_retry_idx;
  wire        _GEN_2678 = _GEN_278 & stq_idx == 5'h0;
  wire        _GEN_2679 = _GEN_278 & stq_idx == 5'h1;
  wire        _GEN_2680 = _GEN_278 & stq_idx == 5'h2;
  wire        _GEN_2681 = _GEN_278 & stq_idx == 5'h3;
  wire        _GEN_2682 = _GEN_278 & stq_idx == 5'h4;
  wire        _GEN_2683 = _GEN_278 & stq_idx == 5'h5;
  wire        _GEN_2684 = _GEN_278 & stq_idx == 5'h6;
  wire        _GEN_2685 = _GEN_278 & stq_idx == 5'h7;
  wire        _GEN_2686 = _GEN_278 & stq_idx == 5'h8;
  wire        _GEN_2687 = _GEN_278 & stq_idx == 5'h9;
  wire        _GEN_2688 = _GEN_278 & stq_idx == 5'hA;
  wire        _GEN_2689 = _GEN_278 & stq_idx == 5'hB;
  wire        _GEN_2690 = _GEN_278 & stq_idx == 5'hC;
  wire        _GEN_2691 = _GEN_278 & stq_idx == 5'hD;
  wire        _GEN_2692 = _GEN_278 & stq_idx == 5'hE;
  wire        _GEN_2693 = _GEN_278 & stq_idx == 5'hF;
  wire        _GEN_2694 = _GEN_278 & stq_idx == 5'h10;
  wire        _GEN_2695 = _GEN_278 & stq_idx == 5'h11;
  wire        _GEN_2696 = _GEN_278 & stq_idx == 5'h12;
  wire        _GEN_2697 = _GEN_278 & stq_idx == 5'h13;
  wire        _GEN_2698 = _GEN_278 & stq_idx == 5'h14;
  wire        _GEN_2699 = _GEN_278 & stq_idx == 5'h15;
  wire        _GEN_2700 = _GEN_278 & stq_idx == 5'h16;
  wire        _GEN_2701 = _GEN_278 & stq_idx == 5'h17;
  wire        _GEN_2702 = _GEN_278 & stq_idx == 5'h18;
  wire        _GEN_2703 = _GEN_278 & stq_idx == 5'h19;
  wire        _GEN_2704 = _GEN_278 & stq_idx == 5'h1A;
  wire        _GEN_2705 = _GEN_278 & stq_idx == 5'h1B;
  wire        _GEN_2706 = _GEN_278 & stq_idx == 5'h1C;
  wire        _GEN_2707 = _GEN_278 & stq_idx == 5'h1D;
  wire        _GEN_2708 = _GEN_278 & stq_idx == 5'h1E;
  wire        _GEN_2709 = _GEN_278 & (&stq_idx);
  wire        _GEN_2710 = _GEN_279 & sidx == 5'h0;
  wire        _GEN_2711 = _GEN_279 & sidx == 5'h1;
  wire        _GEN_2712 = _GEN_279 & sidx == 5'h2;
  wire        _GEN_2713 = _GEN_279 & sidx == 5'h3;
  wire        _GEN_2714 = _GEN_279 & sidx == 5'h4;
  wire        _GEN_2715 = _GEN_279 & sidx == 5'h5;
  wire        _GEN_2716 = _GEN_279 & sidx == 5'h6;
  wire        _GEN_2717 = _GEN_279 & sidx == 5'h7;
  wire        _GEN_2718 = _GEN_279 & sidx == 5'h8;
  wire        _GEN_2719 = _GEN_279 & sidx == 5'h9;
  wire        _GEN_2720 = _GEN_279 & sidx == 5'hA;
  wire        _GEN_2721 = _GEN_279 & sidx == 5'hB;
  wire        _GEN_2722 = _GEN_279 & sidx == 5'hC;
  wire        _GEN_2723 = _GEN_279 & sidx == 5'hD;
  wire        _GEN_2724 = _GEN_279 & sidx == 5'hE;
  wire        _GEN_2725 = _GEN_279 & sidx == 5'hF;
  wire        _GEN_2726 = _GEN_279 & sidx == 5'h10;
  wire        _GEN_2727 = _GEN_279 & sidx == 5'h11;
  wire        _GEN_2728 = _GEN_279 & sidx == 5'h12;
  wire        _GEN_2729 = _GEN_279 & sidx == 5'h13;
  wire        _GEN_2730 = _GEN_279 & sidx == 5'h14;
  wire        _GEN_2731 = _GEN_279 & sidx == 5'h15;
  wire        _GEN_2732 = _GEN_279 & sidx == 5'h16;
  wire        _GEN_2733 = _GEN_279 & sidx == 5'h17;
  wire        _GEN_2734 = _GEN_279 & sidx == 5'h18;
  wire        _GEN_2735 = _GEN_279 & sidx == 5'h19;
  wire        _GEN_2736 = _GEN_279 & sidx == 5'h1A;
  wire        _GEN_2737 = _GEN_279 & sidx == 5'h1B;
  wire        _GEN_2738 = _GEN_279 & sidx == 5'h1C;
  wire        _GEN_2739 = _GEN_279 & sidx == 5'h1D;
  wire        _GEN_2740 = _GEN_279 & sidx == 5'h1E;
  wire        _GEN_2741 = _GEN_279 & (&sidx);
  wire [63:0] _stq_bits_data_bits_T_1 = _stq_bits_data_bits_T ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_data : io_core_exe_0_req_bits_data) : io_core_fp_stdata_bits_data;
  wire [4:0]  ldq_idx_1 = will_fire_load_incoming_1_will_fire ? _mem_incoming_uop_WIRE_1_ldq_idx : ldq_retry_idx;
  wire        _GEN_2742 = ldq_idx_1 == 5'h0;
  wire        _GEN_2743 = _GEN_281 ? _GEN_2742 | _GEN_2646 | _GEN_2326 : _GEN_2646 | _GEN_2326;
  wire        _GEN_2744 = ldq_idx_1 == 5'h1;
  wire        _GEN_2745 = _GEN_281 ? _GEN_2744 | _GEN_2647 | _GEN_2327 : _GEN_2647 | _GEN_2327;
  wire        _GEN_2746 = ldq_idx_1 == 5'h2;
  wire        _GEN_2747 = _GEN_281 ? _GEN_2746 | _GEN_2648 | _GEN_2328 : _GEN_2648 | _GEN_2328;
  wire        _GEN_2748 = ldq_idx_1 == 5'h3;
  wire        _GEN_2749 = _GEN_281 ? _GEN_2748 | _GEN_2649 | _GEN_2329 : _GEN_2649 | _GEN_2329;
  wire        _GEN_2750 = ldq_idx_1 == 5'h4;
  wire        _GEN_2751 = _GEN_281 ? _GEN_2750 | _GEN_2650 | _GEN_2330 : _GEN_2650 | _GEN_2330;
  wire        _GEN_2752 = ldq_idx_1 == 5'h5;
  wire        _GEN_2753 = _GEN_281 ? _GEN_2752 | _GEN_2651 | _GEN_2331 : _GEN_2651 | _GEN_2331;
  wire        _GEN_2754 = ldq_idx_1 == 5'h6;
  wire        _GEN_2755 = _GEN_281 ? _GEN_2754 | _GEN_2652 | _GEN_2332 : _GEN_2652 | _GEN_2332;
  wire        _GEN_2756 = ldq_idx_1 == 5'h7;
  wire        _GEN_2757 = _GEN_281 ? _GEN_2756 | _GEN_2653 | _GEN_2333 : _GEN_2653 | _GEN_2333;
  wire        _GEN_2758 = ldq_idx_1 == 5'h8;
  wire        _GEN_2759 = _GEN_281 ? _GEN_2758 | _GEN_2654 | _GEN_2334 : _GEN_2654 | _GEN_2334;
  wire        _GEN_2760 = ldq_idx_1 == 5'h9;
  wire        _GEN_2761 = _GEN_281 ? _GEN_2760 | _GEN_2655 | _GEN_2335 : _GEN_2655 | _GEN_2335;
  wire        _GEN_2762 = ldq_idx_1 == 5'hA;
  wire        _GEN_2763 = _GEN_281 ? _GEN_2762 | _GEN_2656 | _GEN_2336 : _GEN_2656 | _GEN_2336;
  wire        _GEN_2764 = ldq_idx_1 == 5'hB;
  wire        _GEN_2765 = _GEN_281 ? _GEN_2764 | _GEN_2657 | _GEN_2337 : _GEN_2657 | _GEN_2337;
  wire        _GEN_2766 = ldq_idx_1 == 5'hC;
  wire        _GEN_2767 = _GEN_281 ? _GEN_2766 | _GEN_2658 | _GEN_2338 : _GEN_2658 | _GEN_2338;
  wire        _GEN_2768 = ldq_idx_1 == 5'hD;
  wire        _GEN_2769 = _GEN_281 ? _GEN_2768 | _GEN_2659 | _GEN_2339 : _GEN_2659 | _GEN_2339;
  wire        _GEN_2770 = ldq_idx_1 == 5'hE;
  wire        _GEN_2771 = _GEN_281 ? _GEN_2770 | _GEN_2660 | _GEN_2340 : _GEN_2660 | _GEN_2340;
  wire        _GEN_2772 = ldq_idx_1 == 5'hF;
  wire        _GEN_2773 = _GEN_281 ? _GEN_2772 | _GEN_2661 | _GEN_2341 : _GEN_2661 | _GEN_2341;
  wire        _GEN_2774 = ldq_idx_1 == 5'h10;
  wire        _GEN_2775 = _GEN_281 ? _GEN_2774 | _GEN_2662 | _GEN_2342 : _GEN_2662 | _GEN_2342;
  wire        _GEN_2776 = ldq_idx_1 == 5'h11;
  wire        _GEN_2777 = _GEN_281 ? _GEN_2776 | _GEN_2663 | _GEN_2343 : _GEN_2663 | _GEN_2343;
  wire        _GEN_2778 = ldq_idx_1 == 5'h12;
  wire        _GEN_2779 = _GEN_281 ? _GEN_2778 | _GEN_2664 | _GEN_2344 : _GEN_2664 | _GEN_2344;
  wire        _GEN_2780 = ldq_idx_1 == 5'h13;
  wire        _GEN_2781 = _GEN_281 ? _GEN_2780 | _GEN_2665 | _GEN_2345 : _GEN_2665 | _GEN_2345;
  wire        _GEN_2782 = ldq_idx_1 == 5'h14;
  wire        _GEN_2783 = _GEN_281 ? _GEN_2782 | _GEN_2666 | _GEN_2346 : _GEN_2666 | _GEN_2346;
  wire        _GEN_2784 = ldq_idx_1 == 5'h15;
  wire        _GEN_2785 = _GEN_281 ? _GEN_2784 | _GEN_2667 | _GEN_2347 : _GEN_2667 | _GEN_2347;
  wire        _GEN_2786 = ldq_idx_1 == 5'h16;
  wire        _GEN_2787 = _GEN_281 ? _GEN_2786 | _GEN_2668 | _GEN_2348 : _GEN_2668 | _GEN_2348;
  wire        _GEN_2788 = ldq_idx_1 == 5'h17;
  wire        _GEN_2789 = _GEN_281 ? _GEN_2788 | _GEN_2669 | _GEN_2349 : _GEN_2669 | _GEN_2349;
  wire        _GEN_2790 = ldq_idx_1 == 5'h18;
  wire        _GEN_2791 = _GEN_281 ? _GEN_2790 | _GEN_2670 | _GEN_2350 : _GEN_2670 | _GEN_2350;
  wire        _GEN_2792 = ldq_idx_1 == 5'h19;
  wire        _GEN_2793 = _GEN_281 ? _GEN_2792 | _GEN_2671 | _GEN_2351 : _GEN_2671 | _GEN_2351;
  wire        _GEN_2794 = ldq_idx_1 == 5'h1A;
  wire        _GEN_2795 = _GEN_281 ? _GEN_2794 | _GEN_2672 | _GEN_2352 : _GEN_2672 | _GEN_2352;
  wire        _GEN_2796 = ldq_idx_1 == 5'h1B;
  wire        _GEN_2797 = _GEN_281 ? _GEN_2796 | _GEN_2673 | _GEN_2353 : _GEN_2673 | _GEN_2353;
  wire        _GEN_2798 = ldq_idx_1 == 5'h1C;
  wire        _GEN_2799 = _GEN_281 ? _GEN_2798 | _GEN_2674 | _GEN_2354 : _GEN_2674 | _GEN_2354;
  wire        _GEN_2800 = ldq_idx_1 == 5'h1D;
  wire        _GEN_2801 = _GEN_281 ? _GEN_2800 | _GEN_2675 | _GEN_2355 : _GEN_2675 | _GEN_2355;
  wire        _GEN_2802 = ldq_idx_1 == 5'h1E;
  wire        _GEN_2803 = _GEN_281 ? _GEN_2802 | _GEN_2676 | _GEN_2356 : _GEN_2676 | _GEN_2356;
  wire        _GEN_2804 = _GEN_281 ? (&ldq_idx_1) | _GEN_2677 | _GEN_2357 : _GEN_2677 | _GEN_2357;
  wire        _ldq_bits_addr_is_uncacheable_T_3 = ~_dtlb_io_resp_1_cacheable & ~exe_tlb_miss_1;
  wire [4:0]  stq_idx_1 = _stq_idx_T_1 ? _mem_incoming_uop_WIRE_1_stq_idx : stq_retry_idx;
  wire        _GEN_2805 = _GEN_283 & stq_idx_1 == 5'h0;
  wire        _GEN_2806 = _GEN_2805 ? ~pf_st_1 : _GEN_2678 ? ~pf_st_0 : _GEN_2454 & _GEN_2134 & _GEN_2037 & _GEN_1653 & stq_0_bits_addr_valid;
  wire        _GEN_2807 = _GEN_283 & stq_idx_1 == 5'h1;
  wire        _GEN_2808 = _GEN_2807 ? ~pf_st_1 : _GEN_2679 ? ~pf_st_0 : _GEN_2455 & _GEN_2135 & _GEN_2038 & _GEN_1654 & stq_1_bits_addr_valid;
  wire        _GEN_2809 = _GEN_283 & stq_idx_1 == 5'h2;
  wire        _GEN_2810 = _GEN_2809 ? ~pf_st_1 : _GEN_2680 ? ~pf_st_0 : _GEN_2456 & _GEN_2136 & _GEN_2039 & _GEN_1655 & stq_2_bits_addr_valid;
  wire        _GEN_2811 = _GEN_283 & stq_idx_1 == 5'h3;
  wire        _GEN_2812 = _GEN_2811 ? ~pf_st_1 : _GEN_2681 ? ~pf_st_0 : _GEN_2457 & _GEN_2137 & _GEN_2040 & _GEN_1656 & stq_3_bits_addr_valid;
  wire        _GEN_2813 = _GEN_283 & stq_idx_1 == 5'h4;
  wire        _GEN_2814 = _GEN_2813 ? ~pf_st_1 : _GEN_2682 ? ~pf_st_0 : _GEN_2458 & _GEN_2138 & _GEN_2041 & _GEN_1657 & stq_4_bits_addr_valid;
  wire        _GEN_2815 = _GEN_283 & stq_idx_1 == 5'h5;
  wire        _GEN_2816 = _GEN_2815 ? ~pf_st_1 : _GEN_2683 ? ~pf_st_0 : _GEN_2459 & _GEN_2139 & _GEN_2042 & _GEN_1658 & stq_5_bits_addr_valid;
  wire        _GEN_2817 = _GEN_283 & stq_idx_1 == 5'h6;
  wire        _GEN_2818 = _GEN_2817 ? ~pf_st_1 : _GEN_2684 ? ~pf_st_0 : _GEN_2460 & _GEN_2140 & _GEN_2043 & _GEN_1659 & stq_6_bits_addr_valid;
  wire        _GEN_2819 = _GEN_283 & stq_idx_1 == 5'h7;
  wire        _GEN_2820 = _GEN_2819 ? ~pf_st_1 : _GEN_2685 ? ~pf_st_0 : _GEN_2461 & _GEN_2141 & _GEN_2044 & _GEN_1660 & stq_7_bits_addr_valid;
  wire        _GEN_2821 = _GEN_283 & stq_idx_1 == 5'h8;
  wire        _GEN_2822 = _GEN_2821 ? ~pf_st_1 : _GEN_2686 ? ~pf_st_0 : _GEN_2462 & _GEN_2142 & _GEN_2045 & _GEN_1661 & stq_8_bits_addr_valid;
  wire        _GEN_2823 = _GEN_283 & stq_idx_1 == 5'h9;
  wire        _GEN_2824 = _GEN_2823 ? ~pf_st_1 : _GEN_2687 ? ~pf_st_0 : _GEN_2463 & _GEN_2143 & _GEN_2046 & _GEN_1662 & stq_9_bits_addr_valid;
  wire        _GEN_2825 = _GEN_283 & stq_idx_1 == 5'hA;
  wire        _GEN_2826 = _GEN_2825 ? ~pf_st_1 : _GEN_2688 ? ~pf_st_0 : _GEN_2464 & _GEN_2144 & _GEN_2047 & _GEN_1663 & stq_10_bits_addr_valid;
  wire        _GEN_2827 = _GEN_283 & stq_idx_1 == 5'hB;
  wire        _GEN_2828 = _GEN_2827 ? ~pf_st_1 : _GEN_2689 ? ~pf_st_0 : _GEN_2465 & _GEN_2145 & _GEN_2048 & _GEN_1664 & stq_11_bits_addr_valid;
  wire        _GEN_2829 = _GEN_283 & stq_idx_1 == 5'hC;
  wire        _GEN_2830 = _GEN_2829 ? ~pf_st_1 : _GEN_2690 ? ~pf_st_0 : _GEN_2466 & _GEN_2146 & _GEN_2049 & _GEN_1665 & stq_12_bits_addr_valid;
  wire        _GEN_2831 = _GEN_283 & stq_idx_1 == 5'hD;
  wire        _GEN_2832 = _GEN_2831 ? ~pf_st_1 : _GEN_2691 ? ~pf_st_0 : _GEN_2467 & _GEN_2147 & _GEN_2050 & _GEN_1666 & stq_13_bits_addr_valid;
  wire        _GEN_2833 = _GEN_283 & stq_idx_1 == 5'hE;
  wire        _GEN_2834 = _GEN_2833 ? ~pf_st_1 : _GEN_2692 ? ~pf_st_0 : _GEN_2468 & _GEN_2148 & _GEN_2051 & _GEN_1667 & stq_14_bits_addr_valid;
  wire        _GEN_2835 = _GEN_283 & stq_idx_1 == 5'hF;
  wire        _GEN_2836 = _GEN_2835 ? ~pf_st_1 : _GEN_2693 ? ~pf_st_0 : _GEN_2469 & _GEN_2149 & _GEN_2052 & _GEN_1668 & stq_15_bits_addr_valid;
  wire        _GEN_2837 = _GEN_283 & stq_idx_1 == 5'h10;
  wire        _GEN_2838 = _GEN_2837 ? ~pf_st_1 : _GEN_2694 ? ~pf_st_0 : _GEN_2470 & _GEN_2150 & _GEN_2053 & _GEN_1669 & stq_16_bits_addr_valid;
  wire        _GEN_2839 = _GEN_283 & stq_idx_1 == 5'h11;
  wire        _GEN_2840 = _GEN_2839 ? ~pf_st_1 : _GEN_2695 ? ~pf_st_0 : _GEN_2471 & _GEN_2151 & _GEN_2054 & _GEN_1670 & stq_17_bits_addr_valid;
  wire        _GEN_2841 = _GEN_283 & stq_idx_1 == 5'h12;
  wire        _GEN_2842 = _GEN_2841 ? ~pf_st_1 : _GEN_2696 ? ~pf_st_0 : _GEN_2472 & _GEN_2152 & _GEN_2055 & _GEN_1671 & stq_18_bits_addr_valid;
  wire        _GEN_2843 = _GEN_283 & stq_idx_1 == 5'h13;
  wire        _GEN_2844 = _GEN_2843 ? ~pf_st_1 : _GEN_2697 ? ~pf_st_0 : _GEN_2473 & _GEN_2153 & _GEN_2056 & _GEN_1672 & stq_19_bits_addr_valid;
  wire        _GEN_2845 = _GEN_283 & stq_idx_1 == 5'h14;
  wire        _GEN_2846 = _GEN_2845 ? ~pf_st_1 : _GEN_2698 ? ~pf_st_0 : _GEN_2474 & _GEN_2154 & _GEN_2057 & _GEN_1673 & stq_20_bits_addr_valid;
  wire        _GEN_2847 = _GEN_283 & stq_idx_1 == 5'h15;
  wire        _GEN_2848 = _GEN_2847 ? ~pf_st_1 : _GEN_2699 ? ~pf_st_0 : _GEN_2475 & _GEN_2155 & _GEN_2058 & _GEN_1674 & stq_21_bits_addr_valid;
  wire        _GEN_2849 = _GEN_283 & stq_idx_1 == 5'h16;
  wire        _GEN_2850 = _GEN_2849 ? ~pf_st_1 : _GEN_2700 ? ~pf_st_0 : _GEN_2476 & _GEN_2156 & _GEN_2059 & _GEN_1675 & stq_22_bits_addr_valid;
  wire        _GEN_2851 = _GEN_283 & stq_idx_1 == 5'h17;
  wire        _GEN_2852 = _GEN_2851 ? ~pf_st_1 : _GEN_2701 ? ~pf_st_0 : _GEN_2477 & _GEN_2157 & _GEN_2060 & _GEN_1676 & stq_23_bits_addr_valid;
  wire        _GEN_2853 = _GEN_283 & stq_idx_1 == 5'h18;
  wire        _GEN_2854 = _GEN_2853 ? ~pf_st_1 : _GEN_2702 ? ~pf_st_0 : _GEN_2478 & _GEN_2158 & _GEN_2061 & _GEN_1677 & stq_24_bits_addr_valid;
  wire        _GEN_2855 = _GEN_283 & stq_idx_1 == 5'h19;
  wire        _GEN_2856 = _GEN_2855 ? ~pf_st_1 : _GEN_2703 ? ~pf_st_0 : _GEN_2479 & _GEN_2159 & _GEN_2062 & _GEN_1678 & stq_25_bits_addr_valid;
  wire        _GEN_2857 = _GEN_283 & stq_idx_1 == 5'h1A;
  wire        _GEN_2858 = _GEN_2857 ? ~pf_st_1 : _GEN_2704 ? ~pf_st_0 : _GEN_2480 & _GEN_2160 & _GEN_2063 & _GEN_1679 & stq_26_bits_addr_valid;
  wire        _GEN_2859 = _GEN_283 & stq_idx_1 == 5'h1B;
  wire        _GEN_2860 = _GEN_2859 ? ~pf_st_1 : _GEN_2705 ? ~pf_st_0 : _GEN_2481 & _GEN_2161 & _GEN_2064 & _GEN_1680 & stq_27_bits_addr_valid;
  wire        _GEN_2861 = _GEN_283 & stq_idx_1 == 5'h1C;
  wire        _GEN_2862 = _GEN_2861 ? ~pf_st_1 : _GEN_2706 ? ~pf_st_0 : _GEN_2482 & _GEN_2162 & _GEN_2065 & _GEN_1681 & stq_28_bits_addr_valid;
  wire        _GEN_2863 = _GEN_283 & stq_idx_1 == 5'h1D;
  wire        _GEN_2864 = _GEN_2863 ? ~pf_st_1 : _GEN_2707 ? ~pf_st_0 : _GEN_2483 & _GEN_2163 & _GEN_2066 & _GEN_1682 & stq_29_bits_addr_valid;
  wire        _GEN_2865 = _GEN_283 & stq_idx_1 == 5'h1E;
  wire        _GEN_2866 = _GEN_2865 ? ~pf_st_1 : _GEN_2708 ? ~pf_st_0 : _GEN_2484 & _GEN_2164 & _GEN_2067 & _GEN_1683 & stq_30_bits_addr_valid;
  wire        _GEN_2867 = _GEN_283 & (&stq_idx_1);
  wire        _GEN_2868 = _GEN_2867 ? ~pf_st_1 : _GEN_2709 ? ~pf_st_0 : _GEN_2485 & _GEN_2165 & _GEN_2068 & _GEN_1684 & stq_31_bits_addr_valid;
  wire        _GEN_2869 = sidx_1 == 5'h0;
  wire        _GEN_2870 = _stq_bits_data_bits_T_2 ? _GEN_2869 | _GEN_2710 | _GEN_2486 : _GEN_2710 | _GEN_2486;
  wire        _GEN_2871 = sidx_1 == 5'h1;
  wire        _GEN_2872 = _stq_bits_data_bits_T_2 ? _GEN_2871 | _GEN_2711 | _GEN_2487 : _GEN_2711 | _GEN_2487;
  wire        _GEN_2873 = sidx_1 == 5'h2;
  wire        _GEN_2874 = _stq_bits_data_bits_T_2 ? _GEN_2873 | _GEN_2712 | _GEN_2488 : _GEN_2712 | _GEN_2488;
  wire        _GEN_2875 = sidx_1 == 5'h3;
  wire        _GEN_2876 = _stq_bits_data_bits_T_2 ? _GEN_2875 | _GEN_2713 | _GEN_2489 : _GEN_2713 | _GEN_2489;
  wire        _GEN_2877 = sidx_1 == 5'h4;
  wire        _GEN_2878 = _stq_bits_data_bits_T_2 ? _GEN_2877 | _GEN_2714 | _GEN_2490 : _GEN_2714 | _GEN_2490;
  wire        _GEN_2879 = sidx_1 == 5'h5;
  wire        _GEN_2880 = _stq_bits_data_bits_T_2 ? _GEN_2879 | _GEN_2715 | _GEN_2491 : _GEN_2715 | _GEN_2491;
  wire        _GEN_2881 = sidx_1 == 5'h6;
  wire        _GEN_2882 = _stq_bits_data_bits_T_2 ? _GEN_2881 | _GEN_2716 | _GEN_2492 : _GEN_2716 | _GEN_2492;
  wire        _GEN_2883 = sidx_1 == 5'h7;
  wire        _GEN_2884 = _stq_bits_data_bits_T_2 ? _GEN_2883 | _GEN_2717 | _GEN_2493 : _GEN_2717 | _GEN_2493;
  wire        _GEN_2885 = sidx_1 == 5'h8;
  wire        _GEN_2886 = _stq_bits_data_bits_T_2 ? _GEN_2885 | _GEN_2718 | _GEN_2494 : _GEN_2718 | _GEN_2494;
  wire        _GEN_2887 = sidx_1 == 5'h9;
  wire        _GEN_2888 = _stq_bits_data_bits_T_2 ? _GEN_2887 | _GEN_2719 | _GEN_2495 : _GEN_2719 | _GEN_2495;
  wire        _GEN_2889 = sidx_1 == 5'hA;
  wire        _GEN_2890 = _stq_bits_data_bits_T_2 ? _GEN_2889 | _GEN_2720 | _GEN_2496 : _GEN_2720 | _GEN_2496;
  wire        _GEN_2891 = sidx_1 == 5'hB;
  wire        _GEN_2892 = _stq_bits_data_bits_T_2 ? _GEN_2891 | _GEN_2721 | _GEN_2497 : _GEN_2721 | _GEN_2497;
  wire        _GEN_2893 = sidx_1 == 5'hC;
  wire        _GEN_2894 = _stq_bits_data_bits_T_2 ? _GEN_2893 | _GEN_2722 | _GEN_2498 : _GEN_2722 | _GEN_2498;
  wire        _GEN_2895 = sidx_1 == 5'hD;
  wire        _GEN_2896 = _stq_bits_data_bits_T_2 ? _GEN_2895 | _GEN_2723 | _GEN_2499 : _GEN_2723 | _GEN_2499;
  wire        _GEN_2897 = sidx_1 == 5'hE;
  wire        _GEN_2898 = _stq_bits_data_bits_T_2 ? _GEN_2897 | _GEN_2724 | _GEN_2500 : _GEN_2724 | _GEN_2500;
  wire        _GEN_2899 = sidx_1 == 5'hF;
  wire        _GEN_2900 = _stq_bits_data_bits_T_2 ? _GEN_2899 | _GEN_2725 | _GEN_2501 : _GEN_2725 | _GEN_2501;
  wire        _GEN_2901 = sidx_1 == 5'h10;
  wire        _GEN_2902 = _stq_bits_data_bits_T_2 ? _GEN_2901 | _GEN_2726 | _GEN_2502 : _GEN_2726 | _GEN_2502;
  wire        _GEN_2903 = sidx_1 == 5'h11;
  wire        _GEN_2904 = _stq_bits_data_bits_T_2 ? _GEN_2903 | _GEN_2727 | _GEN_2503 : _GEN_2727 | _GEN_2503;
  wire        _GEN_2905 = sidx_1 == 5'h12;
  wire        _GEN_2906 = _stq_bits_data_bits_T_2 ? _GEN_2905 | _GEN_2728 | _GEN_2504 : _GEN_2728 | _GEN_2504;
  wire        _GEN_2907 = sidx_1 == 5'h13;
  wire        _GEN_2908 = _stq_bits_data_bits_T_2 ? _GEN_2907 | _GEN_2729 | _GEN_2505 : _GEN_2729 | _GEN_2505;
  wire        _GEN_2909 = sidx_1 == 5'h14;
  wire        _GEN_2910 = _stq_bits_data_bits_T_2 ? _GEN_2909 | _GEN_2730 | _GEN_2506 : _GEN_2730 | _GEN_2506;
  wire        _GEN_2911 = sidx_1 == 5'h15;
  wire        _GEN_2912 = _stq_bits_data_bits_T_2 ? _GEN_2911 | _GEN_2731 | _GEN_2507 : _GEN_2731 | _GEN_2507;
  wire        _GEN_2913 = sidx_1 == 5'h16;
  wire        _GEN_2914 = _stq_bits_data_bits_T_2 ? _GEN_2913 | _GEN_2732 | _GEN_2508 : _GEN_2732 | _GEN_2508;
  wire        _GEN_2915 = sidx_1 == 5'h17;
  wire        _GEN_2916 = _stq_bits_data_bits_T_2 ? _GEN_2915 | _GEN_2733 | _GEN_2509 : _GEN_2733 | _GEN_2509;
  wire        _GEN_2917 = sidx_1 == 5'h18;
  wire        _GEN_2918 = _stq_bits_data_bits_T_2 ? _GEN_2917 | _GEN_2734 | _GEN_2510 : _GEN_2734 | _GEN_2510;
  wire        _GEN_2919 = sidx_1 == 5'h19;
  wire        _GEN_2920 = _stq_bits_data_bits_T_2 ? _GEN_2919 | _GEN_2735 | _GEN_2511 : _GEN_2735 | _GEN_2511;
  wire        _GEN_2921 = sidx_1 == 5'h1A;
  wire        _GEN_2922 = _stq_bits_data_bits_T_2 ? _GEN_2921 | _GEN_2736 | _GEN_2512 : _GEN_2736 | _GEN_2512;
  wire        _GEN_2923 = sidx_1 == 5'h1B;
  wire        _GEN_2924 = _stq_bits_data_bits_T_2 ? _GEN_2923 | _GEN_2737 | _GEN_2513 : _GEN_2737 | _GEN_2513;
  wire        _GEN_2925 = sidx_1 == 5'h1C;
  wire        _GEN_2926 = _stq_bits_data_bits_T_2 ? _GEN_2925 | _GEN_2738 | _GEN_2514 : _GEN_2738 | _GEN_2514;
  wire        _GEN_2927 = sidx_1 == 5'h1D;
  wire        _GEN_2928 = _stq_bits_data_bits_T_2 ? _GEN_2927 | _GEN_2739 | _GEN_2515 : _GEN_2739 | _GEN_2515;
  wire        _GEN_2929 = sidx_1 == 5'h1E;
  wire        _GEN_2930 = _stq_bits_data_bits_T_2 ? _GEN_2929 | _GEN_2740 | _GEN_2516 : _GEN_2740 | _GEN_2516;
  wire        _GEN_2931 = _stq_bits_data_bits_T_2 ? (&sidx_1) | _GEN_2741 | _GEN_2517 : _GEN_2741 | _GEN_2517;
  wire [63:0] _stq_bits_data_bits_T_3 = _stq_bits_data_bits_T_2 ? (_GEN_17 ? io_core_exe_1_req_bits_data : io_core_exe_0_req_bits_data) : io_core_fp_stdata_bits_data;
  wire        _fired_std_incoming_T = (io_core_brupdate_b1_mispredict_mask & exe_req_0_bits_uop_br_mask) == 20'h0;
  wire        _fired_std_incoming_T_2 = (io_core_brupdate_b1_mispredict_mask & exe_req_1_bits_uop_br_mask) == 20'h0;
  wire [19:0] _mem_ldq_retry_e_out_valid_T = io_core_brupdate_b1_mispredict_mask & casez_tmp_148;
  wire [19:0] _mem_stq_retry_e_out_valid_T = io_core_brupdate_b1_mispredict_mask & casez_tmp_234;
  wire [19:0] _mem_ldq_wakeup_e_out_valid_T = io_core_brupdate_b1_mispredict_mask & casez_tmp_318;
  wire        _GEN_2932 = _GEN_284 ? _GEN_2358 : _GEN_289 ? _GEN_290 | _GEN_2358 : _GEN_291 & searcher_is_older & _GEN_292 | _GEN_2358;
  wire        _GEN_2933 = _GEN_367 ? _GEN_2359 : _GEN_371 ? _GEN_372 | _GEN_2359 : _GEN_373 & searcher_is_older_2 & _GEN_374 | _GEN_2359;
  wire        _GEN_2934 = _GEN_390 ? _GEN_2360 : _GEN_394 ? _GEN_395 | _GEN_2360 : _GEN_396 & searcher_is_older_4 & _GEN_397 | _GEN_2360;
  wire        _GEN_2935 = _GEN_413 ? _GEN_2361 : _GEN_417 ? _GEN_418 | _GEN_2361 : _GEN_419 & searcher_is_older_6 & _GEN_420 | _GEN_2361;
  wire        _GEN_2936 = _GEN_436 ? _GEN_2362 : _GEN_440 ? _GEN_441 | _GEN_2362 : _GEN_442 & searcher_is_older_8 & _GEN_443 | _GEN_2362;
  wire        _GEN_2937 = _GEN_459 ? _GEN_2363 : _GEN_463 ? _GEN_464 | _GEN_2363 : _GEN_465 & searcher_is_older_10 & _GEN_466 | _GEN_2363;
  wire        _GEN_2938 = _GEN_482 ? _GEN_2364 : _GEN_486 ? _GEN_487 | _GEN_2364 : _GEN_488 & searcher_is_older_12 & _GEN_489 | _GEN_2364;
  wire        _GEN_2939 = _GEN_505 ? _GEN_2365 : _GEN_509 ? _GEN_510 | _GEN_2365 : _GEN_511 & searcher_is_older_14 & _GEN_512 | _GEN_2365;
  wire        _GEN_2940 = _GEN_528 ? _GEN_2366 : _GEN_532 ? _GEN_533 | _GEN_2366 : _GEN_534 & searcher_is_older_16 & _GEN_535 | _GEN_2366;
  wire        _GEN_2941 = _GEN_551 ? _GEN_2367 : _GEN_555 ? _GEN_556 | _GEN_2367 : _GEN_557 & searcher_is_older_18 & _GEN_558 | _GEN_2367;
  wire        _GEN_2942 = _GEN_574 ? _GEN_2368 : _GEN_578 ? _GEN_579 | _GEN_2368 : _GEN_580 & searcher_is_older_20 & _GEN_581 | _GEN_2368;
  wire        _GEN_2943 = _GEN_597 ? _GEN_2369 : _GEN_601 ? _GEN_602 | _GEN_2369 : _GEN_603 & searcher_is_older_22 & _GEN_604 | _GEN_2369;
  wire        _GEN_2944 = _GEN_620 ? _GEN_2370 : _GEN_624 ? _GEN_625 | _GEN_2370 : _GEN_626 & searcher_is_older_24 & _GEN_627 | _GEN_2370;
  wire        _GEN_2945 = _GEN_643 ? _GEN_2371 : _GEN_647 ? _GEN_648 | _GEN_2371 : _GEN_649 & searcher_is_older_26 & _GEN_650 | _GEN_2371;
  wire        _GEN_2946 = _GEN_666 ? _GEN_2372 : _GEN_670 ? _GEN_671 | _GEN_2372 : _GEN_672 & searcher_is_older_28 & _GEN_673 | _GEN_2372;
  wire        _GEN_2947 = _GEN_689 ? _GEN_2373 : _GEN_693 ? _GEN_694 | _GEN_2373 : _GEN_695 & searcher_is_older_30 & _GEN_696 | _GEN_2373;
  wire        _GEN_2948 = _GEN_712 ? _GEN_2374 : _GEN_716 ? _GEN_717 | _GEN_2374 : _GEN_718 & searcher_is_older_32 & _GEN_719 | _GEN_2374;
  wire        _GEN_2949 = _GEN_735 ? _GEN_2375 : _GEN_739 ? _GEN_740 | _GEN_2375 : _GEN_741 & searcher_is_older_34 & _GEN_742 | _GEN_2375;
  wire        _GEN_2950 = _GEN_758 ? _GEN_2376 : _GEN_762 ? _GEN_763 | _GEN_2376 : _GEN_764 & searcher_is_older_36 & _GEN_765 | _GEN_2376;
  wire        _GEN_2951 = _GEN_781 ? _GEN_2377 : _GEN_785 ? _GEN_786 | _GEN_2377 : _GEN_787 & searcher_is_older_38 & _GEN_788 | _GEN_2377;
  wire        _GEN_2952 = _GEN_804 ? _GEN_2378 : _GEN_808 ? _GEN_809 | _GEN_2378 : _GEN_810 & searcher_is_older_40 & _GEN_811 | _GEN_2378;
  wire        _GEN_2953 = _GEN_827 ? _GEN_2379 : _GEN_831 ? _GEN_832 | _GEN_2379 : _GEN_833 & searcher_is_older_42 & _GEN_834 | _GEN_2379;
  wire        _GEN_2954 = _GEN_850 ? _GEN_2380 : _GEN_854 ? _GEN_855 | _GEN_2380 : _GEN_856 & searcher_is_older_44 & _GEN_857 | _GEN_2380;
  wire        _GEN_2955 = _GEN_873 ? _GEN_2381 : _GEN_877 ? _GEN_878 | _GEN_2381 : _GEN_879 & searcher_is_older_46 & _GEN_880 | _GEN_2381;
  wire        _GEN_2956 = _GEN_896 ? _GEN_2382 : _GEN_900 ? _GEN_901 | _GEN_2382 : _GEN_902 & searcher_is_older_48 & _GEN_903 | _GEN_2382;
  wire        _GEN_2957 = _GEN_919 ? _GEN_2383 : _GEN_923 ? _GEN_924 | _GEN_2383 : _GEN_925 & searcher_is_older_50 & _GEN_926 | _GEN_2383;
  wire        _GEN_2958 = _GEN_942 ? _GEN_2384 : _GEN_946 ? _GEN_947 | _GEN_2384 : _GEN_948 & searcher_is_older_52 & _GEN_949 | _GEN_2384;
  wire        _GEN_2959 = _GEN_965 ? _GEN_2385 : _GEN_969 ? _GEN_970 | _GEN_2385 : _GEN_971 & searcher_is_older_54 & _GEN_972 | _GEN_2385;
  wire        _GEN_2960 = _GEN_988 ? _GEN_2386 : _GEN_992 ? _GEN_993 | _GEN_2386 : _GEN_994 & searcher_is_older_56 & _GEN_995 | _GEN_2386;
  wire        _GEN_2961 = _GEN_1011 ? _GEN_2387 : _GEN_1015 ? _GEN_1016 | _GEN_2387 : _GEN_1017 & searcher_is_older_58 & _GEN_1018 | _GEN_2387;
  wire        _GEN_2962 = _GEN_1034 ? _GEN_2388 : _GEN_1038 ? _GEN_1039 | _GEN_2388 : _GEN_1040 & searcher_is_older_60 & _GEN_1041 | _GEN_2388;
  wire        _GEN_2963 =
    (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & (&lcam_ldq_idx_1))) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & (&lcam_ldq_idx_0))) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & (&lcam_ldq_idx_1))) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & (&lcam_ldq_idx_0))) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & (&lcam_ldq_idx_1))) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & (&lcam_ldq_idx_0))) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & (&lcam_ldq_idx_1))) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & (&lcam_ldq_idx_0))) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & (&lcam_ldq_idx_1))) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & (&lcam_ldq_idx_0))) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & (&lcam_ldq_idx_1))) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & (&lcam_ldq_idx_0))) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & (&lcam_ldq_idx_1))) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & (&lcam_ldq_idx_0))) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & (&lcam_ldq_idx_1))) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & (&lcam_ldq_idx_0))) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & (&lcam_ldq_idx_1))) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & (&lcam_ldq_idx_0))) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & (&lcam_ldq_idx_1))) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & (&lcam_ldq_idx_0))) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & (&lcam_ldq_idx_1))) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & (&lcam_ldq_idx_0))) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & (&lcam_ldq_idx_1))) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & (&lcam_ldq_idx_0))) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & (&lcam_ldq_idx_1))) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & (&lcam_ldq_idx_0))) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & (&lcam_ldq_idx_1))) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & (&lcam_ldq_idx_0)))
    & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & (&lcam_ldq_idx_1))) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & (&lcam_ldq_idx_0))) & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & (&lcam_ldq_idx_1))) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & (&lcam_ldq_idx_0))) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & (&lcam_ldq_idx_1))) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & (&lcam_ldq_idx_0))) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & (&lcam_ldq_idx_1))) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & (&lcam_ldq_idx_0))) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & (&lcam_ldq_idx_1))) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & (&lcam_ldq_idx_0))) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & (&lcam_ldq_idx_1))) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & (&lcam_ldq_idx_0))) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & (&lcam_ldq_idx_1))) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & (&lcam_ldq_idx_0))) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & (&lcam_ldq_idx_1))) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & (&lcam_ldq_idx_0))) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & (&lcam_ldq_idx_1))) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & (&lcam_ldq_idx_0))) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & (&lcam_ldq_idx_1))) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & (&lcam_ldq_idx_0))) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & (&lcam_ldq_idx_1))) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & (&lcam_ldq_idx_0))) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & (&lcam_ldq_idx_1))) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & (&lcam_ldq_idx_0))) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & (&lcam_ldq_idx_1))) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & (&lcam_ldq_idx_0))) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & (&lcam_ldq_idx_1))) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & (&lcam_ldq_idx_0))) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & (&lcam_ldq_idx_1)))
    & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & (&lcam_ldq_idx_0))) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & (&lcam_ldq_idx_1))) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & (&lcam_ldq_idx_0))) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & (&lcam_ldq_idx_1))) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & (&lcam_ldq_idx_0))) & s1_executing_loads_31;
  wire        _GEN_2964 = _GEN_1057 ? _GEN_2389 : _GEN_1061 ? _GEN_1062 | _GEN_2389 : _GEN_1063 & searcher_is_older_62 & _GEN_1064 | _GEN_2389;
  wire        _GEN_2965 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & ~(|lcam_ldq_idx_1))) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & ~(|lcam_ldq_idx_0))) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & ~(|lcam_ldq_idx_1))) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & ~(|lcam_ldq_idx_0))) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & ~(|lcam_ldq_idx_1))) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & ~(|lcam_ldq_idx_0))) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & ~(|lcam_ldq_idx_1))) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & ~(|lcam_ldq_idx_0))) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & ~(|lcam_ldq_idx_1))) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & ~(|lcam_ldq_idx_0))) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & ~(|lcam_ldq_idx_1))) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & ~(|lcam_ldq_idx_0))) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & ~(|lcam_ldq_idx_1))) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & ~(|lcam_ldq_idx_0))) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & ~(|lcam_ldq_idx_1))) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & ~(|lcam_ldq_idx_0))) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & ~(|lcam_ldq_idx_1))) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & ~(|lcam_ldq_idx_0))) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & ~(|lcam_ldq_idx_1))) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & ~(|lcam_ldq_idx_0))) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & ~(|lcam_ldq_idx_1))) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & ~(|lcam_ldq_idx_0))) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & ~(|lcam_ldq_idx_1))) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & ~(|lcam_ldq_idx_0))) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & ~(|lcam_ldq_idx_1))) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & ~(|lcam_ldq_idx_0))) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & ~(|lcam_ldq_idx_1)))
    & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & ~(|lcam_ldq_idx_0))) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & ~(|lcam_ldq_idx_1))) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & ~(|lcam_ldq_idx_0))) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & ~(|lcam_ldq_idx_1)));
  wire        _GEN_2966 =
    (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & ~(|lcam_ldq_idx_0))) & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & ~(|lcam_ldq_idx_1))) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & ~(|lcam_ldq_idx_0))) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & ~(|lcam_ldq_idx_1))) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & ~(|lcam_ldq_idx_0))) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & ~(|lcam_ldq_idx_1))) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & ~(|lcam_ldq_idx_0))) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & ~(|lcam_ldq_idx_1))) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & ~(|lcam_ldq_idx_0))) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & ~(|lcam_ldq_idx_1))) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & ~(|lcam_ldq_idx_0))) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & ~(|lcam_ldq_idx_1))) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & ~(|lcam_ldq_idx_0))) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & ~(|lcam_ldq_idx_1))) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & ~(|lcam_ldq_idx_0))) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & ~(|lcam_ldq_idx_1))) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & ~(|lcam_ldq_idx_0))) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & ~(|lcam_ldq_idx_1))) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & ~(|lcam_ldq_idx_0))) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & ~(|lcam_ldq_idx_1))) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & ~(|lcam_ldq_idx_0))) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & ~(|lcam_ldq_idx_1))) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & ~(|lcam_ldq_idx_0))) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & ~(|lcam_ldq_idx_1))) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & ~(|lcam_ldq_idx_0))) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & ~(|lcam_ldq_idx_1))) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & ~(|lcam_ldq_idx_0))) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & ~(|lcam_ldq_idx_1)))
    & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & ~(|lcam_ldq_idx_0))) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & ~(|lcam_ldq_idx_1))) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & ~(|lcam_ldq_idx_0))) & s1_executing_loads_0;
  wire        _GEN_2967 = _GEN_2965 & _GEN_2966;
  wire        _GEN_2968 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_336)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_296)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_336)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_296)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_336)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_296)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_336)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_296)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_336)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_296)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_336)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_296)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_336)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_296)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_336)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_296)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_336)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_296)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_336)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_296)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_336)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_296)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_336)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_296)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_336)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_296)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_336)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_296)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_336)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_296)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_336)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_296))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_336)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_296)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_336)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_296)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_336)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_296)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_336)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_296)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_336)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_296)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_336)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_296)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_336)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_296)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_336)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_296)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_336)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_296)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_336)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_296)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_336)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_296)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_336)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_296)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_336)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_296)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_336)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_296)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_336)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_296)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_336)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_296)) & s1_executing_loads_1;
  wire        _GEN_2969 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_337)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_297)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_337)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_297)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_337)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_297)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_337)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_297)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_337)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_297)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_337)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_297)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_337)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_297)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_337)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_297)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_337)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_297)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_337)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_297)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_337)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_297)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_337)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_297)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_337)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_297)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_337)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_297)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_337)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_297)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_337)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_297))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_337)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_297)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_337)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_297)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_337)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_297)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_337)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_297)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_337)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_297)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_337)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_297)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_337)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_297)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_337)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_297)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_337)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_297)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_337)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_297)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_337)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_297)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_337)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_297)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_337)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_297)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_337)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_297)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_337)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_297)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_337)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_297)) & s1_executing_loads_2;
  wire        _GEN_2970 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_338)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_298)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_338)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_298)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_338)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_298)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_338)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_298)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_338)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_298)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_338)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_298)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_338)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_298)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_338)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_298)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_338)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_298)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_338)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_298)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_338)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_298)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_338)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_298)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_338)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_298)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_338)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_298)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_338)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_298)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_338)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_298))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_338)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_298)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_338)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_298)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_338)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_298)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_338)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_298)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_338)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_298)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_338)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_298)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_338)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_298)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_338)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_298)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_338)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_298)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_338)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_298)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_338)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_298)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_338)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_298)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_338)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_298)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_338)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_298)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_338)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_298)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_338)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_298)) & s1_executing_loads_3;
  wire        _GEN_2971 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_339)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_299)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_339)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_299)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_339)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_299)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_339)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_299)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_339)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_299)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_339)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_299)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_339)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_299)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_339)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_299)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_339)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_299)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_339)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_299)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_339)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_299)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_339)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_299)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_339)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_299)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_339)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_299)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_339)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_299)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_339)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_299))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_339)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_299)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_339)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_299)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_339)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_299)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_339)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_299)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_339)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_299)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_339)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_299)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_339)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_299)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_339)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_299)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_339)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_299)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_339)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_299)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_339)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_299)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_339)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_299)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_339)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_299)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_339)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_299)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_339)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_299)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_339)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_299)) & s1_executing_loads_4;
  wire        _GEN_2972 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_340)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_300)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_340)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_300)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_340)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_300)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_340)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_300)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_340)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_300)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_340)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_300)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_340)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_300)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_340)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_300)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_340)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_300)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_340)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_300)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_340)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_300)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_340)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_300)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_340)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_300)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_340)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_300)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_340)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_300)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_340)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_300))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_340)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_300)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_340)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_300)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_340)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_300)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_340)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_300)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_340)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_300)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_340)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_300)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_340)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_300)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_340)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_300)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_340)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_300)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_340)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_300)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_340)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_300)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_340)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_300)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_340)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_300)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_340)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_300)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_340)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_300)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_340)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_300)) & s1_executing_loads_5;
  wire        _GEN_2973 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_341)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_301)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_341)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_301)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_341)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_301)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_341)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_301)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_341)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_301)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_341)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_301)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_341)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_301)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_341)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_301)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_341)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_301)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_341)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_301)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_341)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_301)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_341)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_301)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_341)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_301)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_341)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_301)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_341)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_301)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_341)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_301))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_341)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_301)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_341)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_301)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_341)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_301)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_341)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_301)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_341)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_301)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_341)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_301)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_341)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_301)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_341)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_301)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_341)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_301)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_341)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_301)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_341)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_301)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_341)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_301)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_341)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_301)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_341)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_301)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_341)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_301)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_341)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_301)) & s1_executing_loads_6;
  wire        _GEN_2974 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_342)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_302)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_342)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_302)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_342)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_302)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_342)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_302)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_342)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_302)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_342)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_302)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_342)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_302)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_342)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_302)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_342)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_302)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_342)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_302)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_342)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_302)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_342)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_302)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_342)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_302)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_342)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_302)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_342)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_302)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_342)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_302))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_342)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_302)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_342)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_302)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_342)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_302)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_342)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_302)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_342)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_302)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_342)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_302)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_342)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_302)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_342)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_302)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_342)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_302)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_342)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_302)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_342)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_302)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_342)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_302)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_342)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_302)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_342)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_302)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_342)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_302)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_342)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_302)) & s1_executing_loads_7;
  wire        _GEN_2975 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_343)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_303)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_343)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_303)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_343)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_303)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_343)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_303)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_343)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_303)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_343)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_303)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_343)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_303)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_343)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_303)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_343)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_303)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_343)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_303)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_343)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_303)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_343)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_303)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_343)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_303)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_343)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_303)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_343)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_303)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_343)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_303))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_343)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_303)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_343)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_303)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_343)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_303)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_343)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_303)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_343)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_303)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_343)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_303)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_343)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_303)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_343)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_303)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_343)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_303)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_343)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_303)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_343)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_303)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_343)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_303)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_343)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_303)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_343)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_303)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_343)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_303)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_343)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_303)) & s1_executing_loads_8;
  wire        _GEN_2976 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_344)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_304)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_344)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_304)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_344)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_304)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_344)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_304)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_344)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_304)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_344)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_304)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_344)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_304)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_344)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_304)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_344)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_304)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_344)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_304)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_344)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_304)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_344)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_304)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_344)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_304)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_344)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_304)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_344)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_304)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_344)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_304))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_344)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_304)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_344)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_304)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_344)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_304)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_344)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_304)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_344)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_304)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_344)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_304)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_344)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_304)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_344)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_304)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_344)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_304)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_344)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_304)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_344)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_304)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_344)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_304)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_344)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_304)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_344)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_304)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_344)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_304)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_344)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_304)) & s1_executing_loads_9;
  wire        _GEN_2977 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_345)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_305)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_345)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_305)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_345)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_305)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_345)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_305)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_345)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_305)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_345)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_305)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_345)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_305)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_345)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_305)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_345)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_305)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_345)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_305)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_345)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_305)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_345)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_305)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_345)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_305)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_345)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_305)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_345)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_305)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_345)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_305))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_345)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_305)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_345)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_305)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_345)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_305)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_345)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_305)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_345)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_305)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_345)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_305)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_345)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_305)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_345)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_305)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_345)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_305)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_345)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_305)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_345)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_305)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_345)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_305)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_345)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_305)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_345)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_305)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_345)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_305)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_345)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_305)) & s1_executing_loads_10;
  wire        _GEN_2978 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_346)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_306)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_346)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_306)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_346)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_306)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_346)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_306)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_346)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_306)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_346)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_306)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_346)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_306)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_346)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_306)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_346)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_306)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_346)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_306)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_346)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_306)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_346)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_306)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_346)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_306)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_346)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_306)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_346)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_306)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_346)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_306))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_346)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_306)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_346)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_306)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_346)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_306)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_346)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_306)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_346)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_306)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_346)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_306)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_346)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_306)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_346)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_306)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_346)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_306)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_346)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_306)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_346)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_306)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_346)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_306)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_346)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_306)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_346)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_306)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_346)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_306)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_346)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_306)) & s1_executing_loads_11;
  wire        _GEN_2979 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_347)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_307)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_347)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_307)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_347)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_307)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_347)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_307)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_347)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_307)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_347)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_307)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_347)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_307)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_347)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_307)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_347)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_307)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_347)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_307)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_347)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_307)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_347)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_307)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_347)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_307)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_347)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_307)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_347)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_307)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_347)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_307))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_347)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_307)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_347)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_307)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_347)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_307)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_347)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_307)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_347)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_307)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_347)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_307)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_347)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_307)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_347)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_307)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_347)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_307)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_347)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_307)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_347)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_307)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_347)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_307)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_347)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_307)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_347)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_307)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_347)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_307)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_347)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_307)) & s1_executing_loads_12;
  wire        _GEN_2980 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_348)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_308)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_348)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_308)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_348)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_308)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_348)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_308)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_348)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_308)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_348)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_308)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_348)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_308)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_348)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_308)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_348)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_308)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_348)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_308)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_348)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_308)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_348)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_308)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_348)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_308)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_348)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_308)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_348)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_308)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_348)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_308))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_348)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_308)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_348)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_308)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_348)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_308)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_348)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_308)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_348)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_308)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_348)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_308)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_348)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_308)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_348)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_308)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_348)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_308)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_348)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_308)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_348)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_308)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_348)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_308)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_348)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_308)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_348)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_308)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_348)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_308)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_348)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_308)) & s1_executing_loads_13;
  wire        _GEN_2981 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_349)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_309)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_349)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_309)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_349)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_309)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_349)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_309)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_349)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_309)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_349)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_309)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_349)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_309)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_349)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_309)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_349)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_309)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_349)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_309)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_349)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_309)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_349)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_309)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_349)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_309)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_349)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_309)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_349)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_309)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_349)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_309))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_349)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_309)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_349)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_309)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_349)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_309)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_349)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_309)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_349)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_309)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_349)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_309)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_349)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_309)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_349)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_309)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_349)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_309)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_349)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_309)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_349)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_309)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_349)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_309)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_349)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_309)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_349)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_309)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_349)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_309)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_349)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_309)) & s1_executing_loads_14;
  wire        _GEN_2982 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_350)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_310)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_350)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_310)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_350)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_310)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_350)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_310)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_350)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_310)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_350)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_310)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_350)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_310)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_350)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_310)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_350)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_310)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_350)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_310)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_350)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_310)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_350)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_310)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_350)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_310)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_350)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_310)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_350)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_310)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_350)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_310))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_350)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_310)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_350)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_310)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_350)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_310)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_350)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_310)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_350)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_310)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_350)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_310)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_350)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_310)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_350)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_310)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_350)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_310)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_350)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_310)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_350)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_310)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_350)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_310)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_350)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_310)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_350)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_310)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_350)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_310)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_350)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_310)) & s1_executing_loads_15;
  wire        _GEN_2983 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_351)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_311)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_351)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_311)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_351)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_311)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_351)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_311)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_351)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_311)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_351)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_311)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_351)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_311)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_351)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_311)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_351)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_311)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_351)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_311)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_351)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_311)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_351)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_311)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_351)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_311)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_351)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_311)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_351)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_311)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_351)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_311))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_351)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_311)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_351)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_311)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_351)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_311)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_351)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_311)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_351)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_311)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_351)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_311)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_351)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_311)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_351)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_311)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_351)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_311)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_351)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_311)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_351)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_311)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_351)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_311)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_351)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_311)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_351)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_311)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_351)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_311)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_351)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_311)) & s1_executing_loads_16;
  wire        _GEN_2984 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_352)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_312)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_352)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_312)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_352)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_312)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_352)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_312)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_352)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_312)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_352)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_312)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_352)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_312)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_352)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_312)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_352)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_312)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_352)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_312)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_352)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_312)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_352)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_312)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_352)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_312)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_352)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_312)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_352)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_312)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_352)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_312))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_352)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_312)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_352)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_312)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_352)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_312)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_352)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_312)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_352)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_312)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_352)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_312)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_352)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_312)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_352)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_312)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_352)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_312)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_352)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_312)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_352)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_312)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_352)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_312)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_352)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_312)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_352)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_312)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_352)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_312)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_352)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_312)) & s1_executing_loads_17;
  wire        _GEN_2985 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_353)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_313)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_353)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_313)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_353)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_313)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_353)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_313)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_353)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_313)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_353)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_313)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_353)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_313)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_353)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_313)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_353)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_313)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_353)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_313)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_353)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_313)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_353)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_313)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_353)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_313)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_353)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_313)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_353)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_313)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_353)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_313))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_353)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_313)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_353)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_313)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_353)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_313)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_353)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_313)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_353)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_313)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_353)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_313)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_353)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_313)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_353)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_313)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_353)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_313)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_353)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_313)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_353)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_313)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_353)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_313)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_353)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_313)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_353)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_313)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_353)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_313)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_353)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_313)) & s1_executing_loads_18;
  wire        _GEN_2986 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_354)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_314)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_354)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_314)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_354)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_314)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_354)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_314)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_354)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_314)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_354)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_314)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_354)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_314)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_354)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_314)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_354)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_314)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_354)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_314)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_354)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_314)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_354)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_314)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_354)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_314)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_354)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_314)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_354)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_314)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_354)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_314))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_354)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_314)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_354)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_314)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_354)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_314)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_354)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_314)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_354)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_314)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_354)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_314)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_354)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_314)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_354)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_314)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_354)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_314)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_354)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_314)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_354)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_314)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_354)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_314)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_354)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_314)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_354)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_314)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_354)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_314)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_354)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_314)) & s1_executing_loads_19;
  wire        _GEN_2987 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_355)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_315)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_355)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_315)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_355)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_315)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_355)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_315)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_355)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_315)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_355)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_315)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_355)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_315)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_355)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_315)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_355)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_315)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_355)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_315)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_355)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_315)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_355)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_315)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_355)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_315)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_355)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_315)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_355)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_315)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_355)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_315))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_355)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_315)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_355)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_315)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_355)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_315)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_355)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_315)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_355)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_315)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_355)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_315)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_355)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_315)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_355)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_315)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_355)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_315)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_355)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_315)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_355)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_315)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_355)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_315)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_355)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_315)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_355)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_315)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_355)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_315)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_355)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_315)) & s1_executing_loads_20;
  wire        _GEN_2988 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_356)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_316)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_356)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_316)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_356)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_316)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_356)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_316)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_356)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_316)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_356)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_316)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_356)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_316)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_356)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_316)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_356)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_316)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_356)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_316)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_356)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_316)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_356)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_316)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_356)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_316)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_356)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_316)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_356)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_316)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_356)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_316))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_356)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_316)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_356)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_316)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_356)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_316)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_356)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_316)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_356)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_316)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_356)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_316)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_356)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_316)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_356)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_316)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_356)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_316)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_356)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_316)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_356)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_316)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_356)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_316)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_356)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_316)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_356)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_316)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_356)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_316)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_356)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_316)) & s1_executing_loads_21;
  wire        _GEN_2989 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_357)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_317)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_357)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_317)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_357)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_317)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_357)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_317)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_357)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_317)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_357)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_317)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_357)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_317)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_357)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_317)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_357)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_317)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_357)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_317)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_357)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_317)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_357)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_317)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_357)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_317)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_357)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_317)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_357)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_317)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_357)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_317))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_357)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_317)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_357)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_317)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_357)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_317)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_357)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_317)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_357)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_317)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_357)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_317)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_357)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_317)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_357)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_317)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_357)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_317)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_357)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_317)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_357)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_317)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_357)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_317)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_357)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_317)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_357)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_317)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_357)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_317)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_357)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_317)) & s1_executing_loads_22;
  wire        _GEN_2990 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_358)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_318)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_358)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_318)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_358)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_318)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_358)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_318)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_358)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_318)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_358)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_318)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_358)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_318)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_358)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_318)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_358)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_318)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_358)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_318)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_358)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_318)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_358)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_318)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_358)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_318)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_358)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_318)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_358)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_318)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_358)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_318))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_358)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_318)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_358)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_318)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_358)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_318)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_358)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_318)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_358)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_318)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_358)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_318)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_358)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_318)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_358)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_318)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_358)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_318)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_358)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_318)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_358)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_318)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_358)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_318)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_358)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_318)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_358)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_318)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_358)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_318)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_358)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_318)) & s1_executing_loads_23;
  wire        _GEN_2991 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_359)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_319)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_359)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_319)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_359)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_319)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_359)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_319)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_359)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_319)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_359)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_319)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_359)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_319)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_359)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_319)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_359)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_319)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_359)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_319)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_359)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_319)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_359)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_319)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_359)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_319)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_359)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_319)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_359)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_319)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_359)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_319))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_359)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_319)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_359)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_319)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_359)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_319)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_359)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_319)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_359)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_319)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_359)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_319)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_359)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_319)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_359)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_319)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_359)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_319)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_359)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_319)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_359)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_319)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_359)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_319)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_359)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_319)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_359)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_319)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_359)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_319)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_359)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_319)) & s1_executing_loads_24;
  wire        _GEN_2992 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_360)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_320)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_360)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_320)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_360)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_320)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_360)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_320)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_360)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_320)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_360)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_320)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_360)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_320)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_360)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_320)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_360)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_320)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_360)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_320)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_360)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_320)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_360)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_320)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_360)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_320)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_360)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_320)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_360)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_320)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_360)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_320))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_360)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_320)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_360)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_320)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_360)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_320)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_360)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_320)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_360)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_320)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_360)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_320)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_360)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_320)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_360)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_320)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_360)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_320)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_360)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_320)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_360)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_320)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_360)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_320)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_360)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_320)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_360)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_320)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_360)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_320)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_360)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_320)) & s1_executing_loads_25;
  wire        _GEN_2993 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_361)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_321)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_361)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_321)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_361)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_321)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_361)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_321)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_361)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_321)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_361)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_321)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_361)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_321)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_361)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_321)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_361)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_321)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_361)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_321)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_361)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_321)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_361)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_321)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_361)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_321)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_361)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_321)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_361)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_321)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_361)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_321))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_361)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_321)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_361)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_321)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_361)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_321)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_361)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_321)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_361)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_321)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_361)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_321)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_361)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_321)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_361)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_321)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_361)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_321)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_361)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_321)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_361)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_321)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_361)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_321)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_361)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_321)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_361)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_321)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_361)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_321)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_361)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_321)) & s1_executing_loads_26;
  wire        _GEN_2994 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_362)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_322)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_362)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_322)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_362)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_322)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_362)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_322)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_362)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_322)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_362)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_322)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_362)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_322)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_362)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_322)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_362)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_322)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_362)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_322)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_362)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_322)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_362)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_322)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_362)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_322)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_362)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_322)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_362)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_322)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_362)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_322))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_362)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_322)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_362)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_322)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_362)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_322)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_362)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_322)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_362)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_322)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_362)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_322)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_362)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_322)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_362)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_322)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_362)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_322)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_362)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_322)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_362)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_322)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_362)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_322)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_362)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_322)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_362)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_322)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_362)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_322)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_362)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_322)) & s1_executing_loads_27;
  wire        _GEN_2995 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_363)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_323)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_363)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_323)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_363)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_323)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_363)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_323)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_363)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_323)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_363)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_323)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_363)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_323)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_363)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_323)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_363)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_323)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_363)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_323)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_363)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_323)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_363)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_323)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_363)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_323)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_363)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_323)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_363)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_323)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_363)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_323))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_363)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_323)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_363)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_323)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_363)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_323)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_363)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_323)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_363)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_323)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_363)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_323)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_363)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_323)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_363)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_323)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_363)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_323)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_363)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_323)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_363)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_323)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_363)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_323)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_363)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_323)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_363)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_323)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_363)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_323)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_363)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_323)) & s1_executing_loads_28;
  wire        _GEN_2996 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_364)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_324)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_364)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_324)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_364)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_324)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_364)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_324)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_364)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_324)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_364)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_324)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_364)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_324)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_364)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_324)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_364)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_324)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_364)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_324)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_364)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_324)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_364)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_324)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_364)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_324)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_364)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_324)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_364)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_324)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_364)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_324))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_364)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_324)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_364)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_324)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_364)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_324)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_364)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_324)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_364)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_324)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_364)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_324)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_364)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_324)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_364)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_324)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_364)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_324)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_364)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_324)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_364)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_324)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_364)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_324)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_364)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_324)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_364)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_324)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_364)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_324)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_364)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_324)) & s1_executing_loads_29;
  wire        _GEN_2997 =
    (_GEN_1077 | ~_GEN_1074 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_1076 & _GEN_365)) & (_GEN_1067 | ~_GEN_1063 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_1066 & _GEN_325)) & (_GEN_1055 | ~_GEN_1051 | _GEN_1054 | ~(_GEN_1053 & _GEN_365)) & (_GEN_1045 | ~_GEN_1040 | _GEN_1044 | ~(_GEN_1043 & _GEN_325)) & (_GEN_1032 | ~_GEN_1028 | _GEN_1031 | ~(_GEN_1030 & _GEN_365)) & (_GEN_1022 | ~_GEN_1017 | _GEN_1021 | ~(_GEN_1020 & _GEN_325)) & (_GEN_1009 | ~_GEN_1005 | _GEN_1008 | ~(_GEN_1007 & _GEN_365)) & (_GEN_999 | ~_GEN_994 | _GEN_998 | ~(_GEN_997 & _GEN_325)) & (_GEN_986 | ~_GEN_982 | _GEN_985 | ~(_GEN_984 & _GEN_365)) & (_GEN_976 | ~_GEN_971 | _GEN_975 | ~(_GEN_974 & _GEN_325)) & (_GEN_963 | ~_GEN_959 | _GEN_962 | ~(_GEN_961 & _GEN_365)) & (_GEN_953 | ~_GEN_948 | _GEN_952 | ~(_GEN_951 & _GEN_325)) & (_GEN_940 | ~_GEN_936 | _GEN_939 | ~(_GEN_938 & _GEN_365)) & (_GEN_930 | ~_GEN_925 | _GEN_929 | ~(_GEN_928 & _GEN_325)) & (_GEN_917 | ~_GEN_913 | _GEN_916 | ~(_GEN_915 & _GEN_365)) & (_GEN_907 | ~_GEN_902 | _GEN_906 | ~(_GEN_905 & _GEN_325)) & (_GEN_894 | ~_GEN_890 | _GEN_893 | ~(_GEN_892 & _GEN_365)) & (_GEN_884 | ~_GEN_879 | _GEN_883 | ~(_GEN_882 & _GEN_325)) & (_GEN_871 | ~_GEN_867 | _GEN_870 | ~(_GEN_869 & _GEN_365)) & (_GEN_861 | ~_GEN_856 | _GEN_860 | ~(_GEN_859 & _GEN_325)) & (_GEN_848 | ~_GEN_844 | _GEN_847 | ~(_GEN_846 & _GEN_365)) & (_GEN_838 | ~_GEN_833 | _GEN_837 | ~(_GEN_836 & _GEN_325)) & (_GEN_825 | ~_GEN_821 | _GEN_824 | ~(_GEN_823 & _GEN_365)) & (_GEN_815 | ~_GEN_810 | _GEN_814 | ~(_GEN_813 & _GEN_325)) & (_GEN_802 | ~_GEN_798 | _GEN_801 | ~(_GEN_800 & _GEN_365)) & (_GEN_792 | ~_GEN_787 | _GEN_791 | ~(_GEN_790 & _GEN_325)) & (_GEN_779 | ~_GEN_775 | _GEN_778 | ~(_GEN_777 & _GEN_365)) & (_GEN_769 | ~_GEN_764 | _GEN_768 | ~(_GEN_767 & _GEN_325)) & (_GEN_756 | ~_GEN_752 | _GEN_755 | ~(_GEN_754 & _GEN_365)) & (_GEN_746 | ~_GEN_741 | _GEN_745 | ~(_GEN_744 & _GEN_325)) & (_GEN_733 | ~_GEN_729 | _GEN_732 | ~(_GEN_731 & _GEN_365)) & (_GEN_723 | ~_GEN_718 | _GEN_722 | ~(_GEN_721 & _GEN_325))
    & (_GEN_710 | ~_GEN_706 | _GEN_709 | ~(_GEN_708 & _GEN_365)) & (_GEN_700 | ~_GEN_695 | _GEN_699 | ~(_GEN_698 & _GEN_325)) & (_GEN_687 | ~_GEN_683 | _GEN_686 | ~(_GEN_685 & _GEN_365)) & (_GEN_677 | ~_GEN_672 | _GEN_676 | ~(_GEN_675 & _GEN_325)) & (_GEN_664 | ~_GEN_660 | _GEN_663 | ~(_GEN_662 & _GEN_365)) & (_GEN_654 | ~_GEN_649 | _GEN_653 | ~(_GEN_652 & _GEN_325)) & (_GEN_641 | ~_GEN_637 | _GEN_640 | ~(_GEN_639 & _GEN_365)) & (_GEN_631 | ~_GEN_626 | _GEN_630 | ~(_GEN_629 & _GEN_325)) & (_GEN_618 | ~_GEN_614 | _GEN_617 | ~(_GEN_616 & _GEN_365)) & (_GEN_608 | ~_GEN_603 | _GEN_607 | ~(_GEN_606 & _GEN_325)) & (_GEN_595 | ~_GEN_591 | _GEN_594 | ~(_GEN_593 & _GEN_365)) & (_GEN_585 | ~_GEN_580 | _GEN_584 | ~(_GEN_583 & _GEN_325)) & (_GEN_572 | ~_GEN_568 | _GEN_571 | ~(_GEN_570 & _GEN_365)) & (_GEN_562 | ~_GEN_557 | _GEN_561 | ~(_GEN_560 & _GEN_325)) & (_GEN_549 | ~_GEN_545 | _GEN_548 | ~(_GEN_547 & _GEN_365)) & (_GEN_539 | ~_GEN_534 | _GEN_538 | ~(_GEN_537 & _GEN_325)) & (_GEN_526 | ~_GEN_522 | _GEN_525 | ~(_GEN_524 & _GEN_365)) & (_GEN_516 | ~_GEN_511 | _GEN_515 | ~(_GEN_514 & _GEN_325)) & (_GEN_503 | ~_GEN_499 | _GEN_502 | ~(_GEN_501 & _GEN_365)) & (_GEN_493 | ~_GEN_488 | _GEN_492 | ~(_GEN_491 & _GEN_325)) & (_GEN_480 | ~_GEN_476 | _GEN_479 | ~(_GEN_478 & _GEN_365)) & (_GEN_470 | ~_GEN_465 | _GEN_469 | ~(_GEN_468 & _GEN_325)) & (_GEN_457 | ~_GEN_453 | _GEN_456 | ~(_GEN_455 & _GEN_365)) & (_GEN_447 | ~_GEN_442 | _GEN_446 | ~(_GEN_445 & _GEN_325)) & (_GEN_434 | ~_GEN_430 | _GEN_433 | ~(_GEN_432 & _GEN_365)) & (_GEN_424 | ~_GEN_419 | _GEN_423 | ~(_GEN_422 & _GEN_325)) & (_GEN_411 | ~_GEN_407 | _GEN_410 | ~(_GEN_409 & _GEN_365)) & (_GEN_401 | ~_GEN_396 | _GEN_400 | ~(_GEN_399 & _GEN_325)) & (_GEN_388 | ~_GEN_384 | _GEN_387 | ~(_GEN_386 & _GEN_365)) & (_GEN_378 | ~_GEN_373 | _GEN_377 | ~(_GEN_376 & _GEN_325)) & (_GEN_335 | ~_GEN_332 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_334 & _GEN_365)) & (_GEN_295 | ~_GEN_291 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_294 & _GEN_325)) & s1_executing_loads_30;
  wire        _GEN_2998 = _GEN_1082 | _GEN_1083;
  wire        _GEN_2999 = _GEN_1080 ? (_GEN_2998 ? (|lcam_ldq_idx_0) & _GEN_2967 : ~(_GEN_1084 & ~(|lcam_ldq_idx_0)) & _GEN_2967) : _GEN_2967;
  wire        _GEN_3000 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_296 & _GEN_2968 : ~(_GEN_1084 & _GEN_296) & _GEN_2968) : _GEN_2968;
  wire        _GEN_3001 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_297 & _GEN_2969 : ~(_GEN_1084 & _GEN_297) & _GEN_2969) : _GEN_2969;
  wire        _GEN_3002 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_298 & _GEN_2970 : ~(_GEN_1084 & _GEN_298) & _GEN_2970) : _GEN_2970;
  wire        _GEN_3003 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_299 & _GEN_2971 : ~(_GEN_1084 & _GEN_299) & _GEN_2971) : _GEN_2971;
  wire        _GEN_3004 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_300 & _GEN_2972 : ~(_GEN_1084 & _GEN_300) & _GEN_2972) : _GEN_2972;
  wire        _GEN_3005 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_301 & _GEN_2973 : ~(_GEN_1084 & _GEN_301) & _GEN_2973) : _GEN_2973;
  wire        _GEN_3006 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_302 & _GEN_2974 : ~(_GEN_1084 & _GEN_302) & _GEN_2974) : _GEN_2974;
  wire        _GEN_3007 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_303 & _GEN_2975 : ~(_GEN_1084 & _GEN_303) & _GEN_2975) : _GEN_2975;
  wire        _GEN_3008 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_304 & _GEN_2976 : ~(_GEN_1084 & _GEN_304) & _GEN_2976) : _GEN_2976;
  wire        _GEN_3009 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_305 & _GEN_2977 : ~(_GEN_1084 & _GEN_305) & _GEN_2977) : _GEN_2977;
  wire        _GEN_3010 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_306 & _GEN_2978 : ~(_GEN_1084 & _GEN_306) & _GEN_2978) : _GEN_2978;
  wire        _GEN_3011 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_307 & _GEN_2979 : ~(_GEN_1084 & _GEN_307) & _GEN_2979) : _GEN_2979;
  wire        _GEN_3012 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_308 & _GEN_2980 : ~(_GEN_1084 & _GEN_308) & _GEN_2980) : _GEN_2980;
  wire        _GEN_3013 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_309 & _GEN_2981 : ~(_GEN_1084 & _GEN_309) & _GEN_2981) : _GEN_2981;
  wire        _GEN_3014 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_310 & _GEN_2982 : ~(_GEN_1084 & _GEN_310) & _GEN_2982) : _GEN_2982;
  wire        _GEN_3015 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_311 & _GEN_2983 : ~(_GEN_1084 & _GEN_311) & _GEN_2983) : _GEN_2983;
  wire        _GEN_3016 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_312 & _GEN_2984 : ~(_GEN_1084 & _GEN_312) & _GEN_2984) : _GEN_2984;
  wire        _GEN_3017 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_313 & _GEN_2985 : ~(_GEN_1084 & _GEN_313) & _GEN_2985) : _GEN_2985;
  wire        _GEN_3018 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_314 & _GEN_2986 : ~(_GEN_1084 & _GEN_314) & _GEN_2986) : _GEN_2986;
  wire        _GEN_3019 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_315 & _GEN_2987 : ~(_GEN_1084 & _GEN_315) & _GEN_2987) : _GEN_2987;
  wire        _GEN_3020 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_316 & _GEN_2988 : ~(_GEN_1084 & _GEN_316) & _GEN_2988) : _GEN_2988;
  wire        _GEN_3021 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_317 & _GEN_2989 : ~(_GEN_1084 & _GEN_317) & _GEN_2989) : _GEN_2989;
  wire        _GEN_3022 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_318 & _GEN_2990 : ~(_GEN_1084 & _GEN_318) & _GEN_2990) : _GEN_2990;
  wire        _GEN_3023 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_319 & _GEN_2991 : ~(_GEN_1084 & _GEN_319) & _GEN_2991) : _GEN_2991;
  wire        _GEN_3024 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_320 & _GEN_2992 : ~(_GEN_1084 & _GEN_320) & _GEN_2992) : _GEN_2992;
  wire        _GEN_3025 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_321 & _GEN_2993 : ~(_GEN_1084 & _GEN_321) & _GEN_2993) : _GEN_2993;
  wire        _GEN_3026 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_322 & _GEN_2994 : ~(_GEN_1084 & _GEN_322) & _GEN_2994) : _GEN_2994;
  wire        _GEN_3027 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_323 & _GEN_2995 : ~(_GEN_1084 & _GEN_323) & _GEN_2995) : _GEN_2995;
  wire        _GEN_3028 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_324 & _GEN_2996 : ~(_GEN_1084 & _GEN_324) & _GEN_2996) : _GEN_2996;
  wire        _GEN_3029 = _GEN_1080 ? (_GEN_2998 ? ~_GEN_325 & _GEN_2997 : ~(_GEN_1084 & _GEN_325) & _GEN_2997) : _GEN_2997;
  wire        _GEN_3030 = _GEN_1080 ? (_GEN_2998 ? ~(&lcam_ldq_idx_0) & _GEN_2963 : ~(_GEN_1084 & (&lcam_ldq_idx_0)) & _GEN_2963) : _GEN_2963;
  wire        _GEN_3031 = _GEN_1088 | _GEN_1089;
  wire        _GEN_3032 = _GEN_1086 ? (_GEN_3031 ? (|lcam_ldq_idx_1) & _GEN_2999 : ~(_GEN_1084 & ~(|lcam_ldq_idx_1)) & _GEN_2999) : _GEN_2999;
  wire        _GEN_3033 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_336 & _GEN_3000 : ~(_GEN_1084 & _GEN_336) & _GEN_3000) : _GEN_3000;
  wire        _GEN_3034 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_337 & _GEN_3001 : ~(_GEN_1084 & _GEN_337) & _GEN_3001) : _GEN_3001;
  wire        _GEN_3035 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_338 & _GEN_3002 : ~(_GEN_1084 & _GEN_338) & _GEN_3002) : _GEN_3002;
  wire        _GEN_3036 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_339 & _GEN_3003 : ~(_GEN_1084 & _GEN_339) & _GEN_3003) : _GEN_3003;
  wire        _GEN_3037 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_340 & _GEN_3004 : ~(_GEN_1084 & _GEN_340) & _GEN_3004) : _GEN_3004;
  wire        _GEN_3038 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_341 & _GEN_3005 : ~(_GEN_1084 & _GEN_341) & _GEN_3005) : _GEN_3005;
  wire        _GEN_3039 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_342 & _GEN_3006 : ~(_GEN_1084 & _GEN_342) & _GEN_3006) : _GEN_3006;
  wire        _GEN_3040 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_343 & _GEN_3007 : ~(_GEN_1084 & _GEN_343) & _GEN_3007) : _GEN_3007;
  wire        _GEN_3041 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_344 & _GEN_3008 : ~(_GEN_1084 & _GEN_344) & _GEN_3008) : _GEN_3008;
  wire        _GEN_3042 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_345 & _GEN_3009 : ~(_GEN_1084 & _GEN_345) & _GEN_3009) : _GEN_3009;
  wire        _GEN_3043 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_346 & _GEN_3010 : ~(_GEN_1084 & _GEN_346) & _GEN_3010) : _GEN_3010;
  wire        _GEN_3044 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_347 & _GEN_3011 : ~(_GEN_1084 & _GEN_347) & _GEN_3011) : _GEN_3011;
  wire        _GEN_3045 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_348 & _GEN_3012 : ~(_GEN_1084 & _GEN_348) & _GEN_3012) : _GEN_3012;
  wire        _GEN_3046 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_349 & _GEN_3013 : ~(_GEN_1084 & _GEN_349) & _GEN_3013) : _GEN_3013;
  wire        _GEN_3047 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_350 & _GEN_3014 : ~(_GEN_1084 & _GEN_350) & _GEN_3014) : _GEN_3014;
  wire        _GEN_3048 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_351 & _GEN_3015 : ~(_GEN_1084 & _GEN_351) & _GEN_3015) : _GEN_3015;
  wire        _GEN_3049 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_352 & _GEN_3016 : ~(_GEN_1084 & _GEN_352) & _GEN_3016) : _GEN_3016;
  wire        _GEN_3050 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_353 & _GEN_3017 : ~(_GEN_1084 & _GEN_353) & _GEN_3017) : _GEN_3017;
  wire        _GEN_3051 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_354 & _GEN_3018 : ~(_GEN_1084 & _GEN_354) & _GEN_3018) : _GEN_3018;
  wire        _GEN_3052 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_355 & _GEN_3019 : ~(_GEN_1084 & _GEN_355) & _GEN_3019) : _GEN_3019;
  wire        _GEN_3053 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_356 & _GEN_3020 : ~(_GEN_1084 & _GEN_356) & _GEN_3020) : _GEN_3020;
  wire        _GEN_3054 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_357 & _GEN_3021 : ~(_GEN_1084 & _GEN_357) & _GEN_3021) : _GEN_3021;
  wire        _GEN_3055 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_358 & _GEN_3022 : ~(_GEN_1084 & _GEN_358) & _GEN_3022) : _GEN_3022;
  wire        _GEN_3056 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_359 & _GEN_3023 : ~(_GEN_1084 & _GEN_359) & _GEN_3023) : _GEN_3023;
  wire        _GEN_3057 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_360 & _GEN_3024 : ~(_GEN_1084 & _GEN_360) & _GEN_3024) : _GEN_3024;
  wire        _GEN_3058 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_361 & _GEN_3025 : ~(_GEN_1084 & _GEN_361) & _GEN_3025) : _GEN_3025;
  wire        _GEN_3059 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_362 & _GEN_3026 : ~(_GEN_1084 & _GEN_362) & _GEN_3026) : _GEN_3026;
  wire        _GEN_3060 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_363 & _GEN_3027 : ~(_GEN_1084 & _GEN_363) & _GEN_3027) : _GEN_3027;
  wire        _GEN_3061 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_364 & _GEN_3028 : ~(_GEN_1084 & _GEN_364) & _GEN_3028) : _GEN_3028;
  wire        _GEN_3062 = _GEN_1086 ? (_GEN_3031 ? ~_GEN_365 & _GEN_3029 : ~(_GEN_1084 & _GEN_365) & _GEN_3029) : _GEN_3029;
  wire        _GEN_3063 = _GEN_1086 ? (_GEN_3031 ? ~(&lcam_ldq_idx_1) & _GEN_3030 : ~(_GEN_1084 & (&lcam_ldq_idx_1)) & _GEN_3030) : _GEN_3030;
  wire        _GEN_3064 = _GEN_1093 | _GEN_1094;
  wire        _GEN_3065 = _GEN_1091 ? (_GEN_3064 ? (|lcam_ldq_idx_0) & _GEN_3032 : ~(_GEN_1095 & ~(|lcam_ldq_idx_0)) & _GEN_3032) : _GEN_3032;
  wire        _GEN_3066 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_296 & _GEN_3033 : ~(_GEN_1095 & _GEN_296) & _GEN_3033) : _GEN_3033;
  wire        _GEN_3067 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_297 & _GEN_3034 : ~(_GEN_1095 & _GEN_297) & _GEN_3034) : _GEN_3034;
  wire        _GEN_3068 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_298 & _GEN_3035 : ~(_GEN_1095 & _GEN_298) & _GEN_3035) : _GEN_3035;
  wire        _GEN_3069 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_299 & _GEN_3036 : ~(_GEN_1095 & _GEN_299) & _GEN_3036) : _GEN_3036;
  wire        _GEN_3070 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_300 & _GEN_3037 : ~(_GEN_1095 & _GEN_300) & _GEN_3037) : _GEN_3037;
  wire        _GEN_3071 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_301 & _GEN_3038 : ~(_GEN_1095 & _GEN_301) & _GEN_3038) : _GEN_3038;
  wire        _GEN_3072 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_302 & _GEN_3039 : ~(_GEN_1095 & _GEN_302) & _GEN_3039) : _GEN_3039;
  wire        _GEN_3073 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_303 & _GEN_3040 : ~(_GEN_1095 & _GEN_303) & _GEN_3040) : _GEN_3040;
  wire        _GEN_3074 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_304 & _GEN_3041 : ~(_GEN_1095 & _GEN_304) & _GEN_3041) : _GEN_3041;
  wire        _GEN_3075 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_305 & _GEN_3042 : ~(_GEN_1095 & _GEN_305) & _GEN_3042) : _GEN_3042;
  wire        _GEN_3076 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_306 & _GEN_3043 : ~(_GEN_1095 & _GEN_306) & _GEN_3043) : _GEN_3043;
  wire        _GEN_3077 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_307 & _GEN_3044 : ~(_GEN_1095 & _GEN_307) & _GEN_3044) : _GEN_3044;
  wire        _GEN_3078 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_308 & _GEN_3045 : ~(_GEN_1095 & _GEN_308) & _GEN_3045) : _GEN_3045;
  wire        _GEN_3079 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_309 & _GEN_3046 : ~(_GEN_1095 & _GEN_309) & _GEN_3046) : _GEN_3046;
  wire        _GEN_3080 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_310 & _GEN_3047 : ~(_GEN_1095 & _GEN_310) & _GEN_3047) : _GEN_3047;
  wire        _GEN_3081 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_311 & _GEN_3048 : ~(_GEN_1095 & _GEN_311) & _GEN_3048) : _GEN_3048;
  wire        _GEN_3082 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_312 & _GEN_3049 : ~(_GEN_1095 & _GEN_312) & _GEN_3049) : _GEN_3049;
  wire        _GEN_3083 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_313 & _GEN_3050 : ~(_GEN_1095 & _GEN_313) & _GEN_3050) : _GEN_3050;
  wire        _GEN_3084 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_314 & _GEN_3051 : ~(_GEN_1095 & _GEN_314) & _GEN_3051) : _GEN_3051;
  wire        _GEN_3085 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_315 & _GEN_3052 : ~(_GEN_1095 & _GEN_315) & _GEN_3052) : _GEN_3052;
  wire        _GEN_3086 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_316 & _GEN_3053 : ~(_GEN_1095 & _GEN_316) & _GEN_3053) : _GEN_3053;
  wire        _GEN_3087 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_317 & _GEN_3054 : ~(_GEN_1095 & _GEN_317) & _GEN_3054) : _GEN_3054;
  wire        _GEN_3088 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_318 & _GEN_3055 : ~(_GEN_1095 & _GEN_318) & _GEN_3055) : _GEN_3055;
  wire        _GEN_3089 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_319 & _GEN_3056 : ~(_GEN_1095 & _GEN_319) & _GEN_3056) : _GEN_3056;
  wire        _GEN_3090 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_320 & _GEN_3057 : ~(_GEN_1095 & _GEN_320) & _GEN_3057) : _GEN_3057;
  wire        _GEN_3091 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_321 & _GEN_3058 : ~(_GEN_1095 & _GEN_321) & _GEN_3058) : _GEN_3058;
  wire        _GEN_3092 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_322 & _GEN_3059 : ~(_GEN_1095 & _GEN_322) & _GEN_3059) : _GEN_3059;
  wire        _GEN_3093 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_323 & _GEN_3060 : ~(_GEN_1095 & _GEN_323) & _GEN_3060) : _GEN_3060;
  wire        _GEN_3094 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_324 & _GEN_3061 : ~(_GEN_1095 & _GEN_324) & _GEN_3061) : _GEN_3061;
  wire        _GEN_3095 = _GEN_1091 ? (_GEN_3064 ? ~_GEN_325 & _GEN_3062 : ~(_GEN_1095 & _GEN_325) & _GEN_3062) : _GEN_3062;
  wire        _GEN_3096 = _GEN_1091 ? (_GEN_3064 ? ~(&lcam_ldq_idx_0) & _GEN_3063 : ~(_GEN_1095 & (&lcam_ldq_idx_0)) & _GEN_3063) : _GEN_3063;
  wire        _GEN_3097 = _GEN_1099 | _GEN_1100;
  wire        _GEN_3098 = _GEN_1097 ? (_GEN_3097 ? (|lcam_ldq_idx_1) & _GEN_3065 : ~(_GEN_1095 & ~(|lcam_ldq_idx_1)) & _GEN_3065) : _GEN_3065;
  wire        _GEN_3099 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_336 & _GEN_3066 : ~(_GEN_1095 & _GEN_336) & _GEN_3066) : _GEN_3066;
  wire        _GEN_3100 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_337 & _GEN_3067 : ~(_GEN_1095 & _GEN_337) & _GEN_3067) : _GEN_3067;
  wire        _GEN_3101 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_338 & _GEN_3068 : ~(_GEN_1095 & _GEN_338) & _GEN_3068) : _GEN_3068;
  wire        _GEN_3102 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_339 & _GEN_3069 : ~(_GEN_1095 & _GEN_339) & _GEN_3069) : _GEN_3069;
  wire        _GEN_3103 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_340 & _GEN_3070 : ~(_GEN_1095 & _GEN_340) & _GEN_3070) : _GEN_3070;
  wire        _GEN_3104 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_341 & _GEN_3071 : ~(_GEN_1095 & _GEN_341) & _GEN_3071) : _GEN_3071;
  wire        _GEN_3105 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_342 & _GEN_3072 : ~(_GEN_1095 & _GEN_342) & _GEN_3072) : _GEN_3072;
  wire        _GEN_3106 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_343 & _GEN_3073 : ~(_GEN_1095 & _GEN_343) & _GEN_3073) : _GEN_3073;
  wire        _GEN_3107 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_344 & _GEN_3074 : ~(_GEN_1095 & _GEN_344) & _GEN_3074) : _GEN_3074;
  wire        _GEN_3108 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_345 & _GEN_3075 : ~(_GEN_1095 & _GEN_345) & _GEN_3075) : _GEN_3075;
  wire        _GEN_3109 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_346 & _GEN_3076 : ~(_GEN_1095 & _GEN_346) & _GEN_3076) : _GEN_3076;
  wire        _GEN_3110 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_347 & _GEN_3077 : ~(_GEN_1095 & _GEN_347) & _GEN_3077) : _GEN_3077;
  wire        _GEN_3111 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_348 & _GEN_3078 : ~(_GEN_1095 & _GEN_348) & _GEN_3078) : _GEN_3078;
  wire        _GEN_3112 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_349 & _GEN_3079 : ~(_GEN_1095 & _GEN_349) & _GEN_3079) : _GEN_3079;
  wire        _GEN_3113 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_350 & _GEN_3080 : ~(_GEN_1095 & _GEN_350) & _GEN_3080) : _GEN_3080;
  wire        _GEN_3114 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_351 & _GEN_3081 : ~(_GEN_1095 & _GEN_351) & _GEN_3081) : _GEN_3081;
  wire        _GEN_3115 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_352 & _GEN_3082 : ~(_GEN_1095 & _GEN_352) & _GEN_3082) : _GEN_3082;
  wire        _GEN_3116 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_353 & _GEN_3083 : ~(_GEN_1095 & _GEN_353) & _GEN_3083) : _GEN_3083;
  wire        _GEN_3117 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_354 & _GEN_3084 : ~(_GEN_1095 & _GEN_354) & _GEN_3084) : _GEN_3084;
  wire        _GEN_3118 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_355 & _GEN_3085 : ~(_GEN_1095 & _GEN_355) & _GEN_3085) : _GEN_3085;
  wire        _GEN_3119 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_356 & _GEN_3086 : ~(_GEN_1095 & _GEN_356) & _GEN_3086) : _GEN_3086;
  wire        _GEN_3120 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_357 & _GEN_3087 : ~(_GEN_1095 & _GEN_357) & _GEN_3087) : _GEN_3087;
  wire        _GEN_3121 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_358 & _GEN_3088 : ~(_GEN_1095 & _GEN_358) & _GEN_3088) : _GEN_3088;
  wire        _GEN_3122 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_359 & _GEN_3089 : ~(_GEN_1095 & _GEN_359) & _GEN_3089) : _GEN_3089;
  wire        _GEN_3123 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_360 & _GEN_3090 : ~(_GEN_1095 & _GEN_360) & _GEN_3090) : _GEN_3090;
  wire        _GEN_3124 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_361 & _GEN_3091 : ~(_GEN_1095 & _GEN_361) & _GEN_3091) : _GEN_3091;
  wire        _GEN_3125 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_362 & _GEN_3092 : ~(_GEN_1095 & _GEN_362) & _GEN_3092) : _GEN_3092;
  wire        _GEN_3126 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_363 & _GEN_3093 : ~(_GEN_1095 & _GEN_363) & _GEN_3093) : _GEN_3093;
  wire        _GEN_3127 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_364 & _GEN_3094 : ~(_GEN_1095 & _GEN_364) & _GEN_3094) : _GEN_3094;
  wire        _GEN_3128 = _GEN_1097 ? (_GEN_3097 ? ~_GEN_365 & _GEN_3095 : ~(_GEN_1095 & _GEN_365) & _GEN_3095) : _GEN_3095;
  wire        _GEN_3129 = _GEN_1097 ? (_GEN_3097 ? ~(&lcam_ldq_idx_1) & _GEN_3096 : ~(_GEN_1095 & (&lcam_ldq_idx_1)) & _GEN_3096) : _GEN_3096;
  wire        _GEN_3130 = _GEN_1104 | _GEN_1105;
  wire        _GEN_3131 = _GEN_1102 ? (_GEN_3130 ? (|lcam_ldq_idx_0) & _GEN_3098 : ~(_GEN_1106 & ~(|lcam_ldq_idx_0)) & _GEN_3098) : _GEN_3098;
  wire        _GEN_3132 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_296 & _GEN_3099 : ~(_GEN_1106 & _GEN_296) & _GEN_3099) : _GEN_3099;
  wire        _GEN_3133 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_297 & _GEN_3100 : ~(_GEN_1106 & _GEN_297) & _GEN_3100) : _GEN_3100;
  wire        _GEN_3134 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_298 & _GEN_3101 : ~(_GEN_1106 & _GEN_298) & _GEN_3101) : _GEN_3101;
  wire        _GEN_3135 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_299 & _GEN_3102 : ~(_GEN_1106 & _GEN_299) & _GEN_3102) : _GEN_3102;
  wire        _GEN_3136 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_300 & _GEN_3103 : ~(_GEN_1106 & _GEN_300) & _GEN_3103) : _GEN_3103;
  wire        _GEN_3137 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_301 & _GEN_3104 : ~(_GEN_1106 & _GEN_301) & _GEN_3104) : _GEN_3104;
  wire        _GEN_3138 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_302 & _GEN_3105 : ~(_GEN_1106 & _GEN_302) & _GEN_3105) : _GEN_3105;
  wire        _GEN_3139 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_303 & _GEN_3106 : ~(_GEN_1106 & _GEN_303) & _GEN_3106) : _GEN_3106;
  wire        _GEN_3140 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_304 & _GEN_3107 : ~(_GEN_1106 & _GEN_304) & _GEN_3107) : _GEN_3107;
  wire        _GEN_3141 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_305 & _GEN_3108 : ~(_GEN_1106 & _GEN_305) & _GEN_3108) : _GEN_3108;
  wire        _GEN_3142 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_306 & _GEN_3109 : ~(_GEN_1106 & _GEN_306) & _GEN_3109) : _GEN_3109;
  wire        _GEN_3143 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_307 & _GEN_3110 : ~(_GEN_1106 & _GEN_307) & _GEN_3110) : _GEN_3110;
  wire        _GEN_3144 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_308 & _GEN_3111 : ~(_GEN_1106 & _GEN_308) & _GEN_3111) : _GEN_3111;
  wire        _GEN_3145 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_309 & _GEN_3112 : ~(_GEN_1106 & _GEN_309) & _GEN_3112) : _GEN_3112;
  wire        _GEN_3146 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_310 & _GEN_3113 : ~(_GEN_1106 & _GEN_310) & _GEN_3113) : _GEN_3113;
  wire        _GEN_3147 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_311 & _GEN_3114 : ~(_GEN_1106 & _GEN_311) & _GEN_3114) : _GEN_3114;
  wire        _GEN_3148 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_312 & _GEN_3115 : ~(_GEN_1106 & _GEN_312) & _GEN_3115) : _GEN_3115;
  wire        _GEN_3149 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_313 & _GEN_3116 : ~(_GEN_1106 & _GEN_313) & _GEN_3116) : _GEN_3116;
  wire        _GEN_3150 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_314 & _GEN_3117 : ~(_GEN_1106 & _GEN_314) & _GEN_3117) : _GEN_3117;
  wire        _GEN_3151 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_315 & _GEN_3118 : ~(_GEN_1106 & _GEN_315) & _GEN_3118) : _GEN_3118;
  wire        _GEN_3152 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_316 & _GEN_3119 : ~(_GEN_1106 & _GEN_316) & _GEN_3119) : _GEN_3119;
  wire        _GEN_3153 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_317 & _GEN_3120 : ~(_GEN_1106 & _GEN_317) & _GEN_3120) : _GEN_3120;
  wire        _GEN_3154 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_318 & _GEN_3121 : ~(_GEN_1106 & _GEN_318) & _GEN_3121) : _GEN_3121;
  wire        _GEN_3155 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_319 & _GEN_3122 : ~(_GEN_1106 & _GEN_319) & _GEN_3122) : _GEN_3122;
  wire        _GEN_3156 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_320 & _GEN_3123 : ~(_GEN_1106 & _GEN_320) & _GEN_3123) : _GEN_3123;
  wire        _GEN_3157 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_321 & _GEN_3124 : ~(_GEN_1106 & _GEN_321) & _GEN_3124) : _GEN_3124;
  wire        _GEN_3158 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_322 & _GEN_3125 : ~(_GEN_1106 & _GEN_322) & _GEN_3125) : _GEN_3125;
  wire        _GEN_3159 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_323 & _GEN_3126 : ~(_GEN_1106 & _GEN_323) & _GEN_3126) : _GEN_3126;
  wire        _GEN_3160 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_324 & _GEN_3127 : ~(_GEN_1106 & _GEN_324) & _GEN_3127) : _GEN_3127;
  wire        _GEN_3161 = _GEN_1102 ? (_GEN_3130 ? ~_GEN_325 & _GEN_3128 : ~(_GEN_1106 & _GEN_325) & _GEN_3128) : _GEN_3128;
  wire        _GEN_3162 = _GEN_1102 ? (_GEN_3130 ? ~(&lcam_ldq_idx_0) & _GEN_3129 : ~(_GEN_1106 & (&lcam_ldq_idx_0)) & _GEN_3129) : _GEN_3129;
  wire        _GEN_3163 = _GEN_1110 | _GEN_1111;
  wire        _GEN_3164 = _GEN_1108 ? (_GEN_3163 ? (|lcam_ldq_idx_1) & _GEN_3131 : ~(_GEN_1106 & ~(|lcam_ldq_idx_1)) & _GEN_3131) : _GEN_3131;
  wire        _GEN_3165 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_336 & _GEN_3132 : ~(_GEN_1106 & _GEN_336) & _GEN_3132) : _GEN_3132;
  wire        _GEN_3166 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_337 & _GEN_3133 : ~(_GEN_1106 & _GEN_337) & _GEN_3133) : _GEN_3133;
  wire        _GEN_3167 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_338 & _GEN_3134 : ~(_GEN_1106 & _GEN_338) & _GEN_3134) : _GEN_3134;
  wire        _GEN_3168 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_339 & _GEN_3135 : ~(_GEN_1106 & _GEN_339) & _GEN_3135) : _GEN_3135;
  wire        _GEN_3169 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_340 & _GEN_3136 : ~(_GEN_1106 & _GEN_340) & _GEN_3136) : _GEN_3136;
  wire        _GEN_3170 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_341 & _GEN_3137 : ~(_GEN_1106 & _GEN_341) & _GEN_3137) : _GEN_3137;
  wire        _GEN_3171 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_342 & _GEN_3138 : ~(_GEN_1106 & _GEN_342) & _GEN_3138) : _GEN_3138;
  wire        _GEN_3172 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_343 & _GEN_3139 : ~(_GEN_1106 & _GEN_343) & _GEN_3139) : _GEN_3139;
  wire        _GEN_3173 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_344 & _GEN_3140 : ~(_GEN_1106 & _GEN_344) & _GEN_3140) : _GEN_3140;
  wire        _GEN_3174 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_345 & _GEN_3141 : ~(_GEN_1106 & _GEN_345) & _GEN_3141) : _GEN_3141;
  wire        _GEN_3175 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_346 & _GEN_3142 : ~(_GEN_1106 & _GEN_346) & _GEN_3142) : _GEN_3142;
  wire        _GEN_3176 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_347 & _GEN_3143 : ~(_GEN_1106 & _GEN_347) & _GEN_3143) : _GEN_3143;
  wire        _GEN_3177 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_348 & _GEN_3144 : ~(_GEN_1106 & _GEN_348) & _GEN_3144) : _GEN_3144;
  wire        _GEN_3178 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_349 & _GEN_3145 : ~(_GEN_1106 & _GEN_349) & _GEN_3145) : _GEN_3145;
  wire        _GEN_3179 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_350 & _GEN_3146 : ~(_GEN_1106 & _GEN_350) & _GEN_3146) : _GEN_3146;
  wire        _GEN_3180 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_351 & _GEN_3147 : ~(_GEN_1106 & _GEN_351) & _GEN_3147) : _GEN_3147;
  wire        _GEN_3181 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_352 & _GEN_3148 : ~(_GEN_1106 & _GEN_352) & _GEN_3148) : _GEN_3148;
  wire        _GEN_3182 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_353 & _GEN_3149 : ~(_GEN_1106 & _GEN_353) & _GEN_3149) : _GEN_3149;
  wire        _GEN_3183 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_354 & _GEN_3150 : ~(_GEN_1106 & _GEN_354) & _GEN_3150) : _GEN_3150;
  wire        _GEN_3184 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_355 & _GEN_3151 : ~(_GEN_1106 & _GEN_355) & _GEN_3151) : _GEN_3151;
  wire        _GEN_3185 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_356 & _GEN_3152 : ~(_GEN_1106 & _GEN_356) & _GEN_3152) : _GEN_3152;
  wire        _GEN_3186 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_357 & _GEN_3153 : ~(_GEN_1106 & _GEN_357) & _GEN_3153) : _GEN_3153;
  wire        _GEN_3187 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_358 & _GEN_3154 : ~(_GEN_1106 & _GEN_358) & _GEN_3154) : _GEN_3154;
  wire        _GEN_3188 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_359 & _GEN_3155 : ~(_GEN_1106 & _GEN_359) & _GEN_3155) : _GEN_3155;
  wire        _GEN_3189 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_360 & _GEN_3156 : ~(_GEN_1106 & _GEN_360) & _GEN_3156) : _GEN_3156;
  wire        _GEN_3190 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_361 & _GEN_3157 : ~(_GEN_1106 & _GEN_361) & _GEN_3157) : _GEN_3157;
  wire        _GEN_3191 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_362 & _GEN_3158 : ~(_GEN_1106 & _GEN_362) & _GEN_3158) : _GEN_3158;
  wire        _GEN_3192 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_363 & _GEN_3159 : ~(_GEN_1106 & _GEN_363) & _GEN_3159) : _GEN_3159;
  wire        _GEN_3193 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_364 & _GEN_3160 : ~(_GEN_1106 & _GEN_364) & _GEN_3160) : _GEN_3160;
  wire        _GEN_3194 = _GEN_1108 ? (_GEN_3163 ? ~_GEN_365 & _GEN_3161 : ~(_GEN_1106 & _GEN_365) & _GEN_3161) : _GEN_3161;
  wire        _GEN_3195 = _GEN_1108 ? (_GEN_3163 ? ~(&lcam_ldq_idx_1) & _GEN_3162 : ~(_GEN_1106 & (&lcam_ldq_idx_1)) & _GEN_3162) : _GEN_3162;
  wire        _GEN_3196 = _GEN_1115 | _GEN_1116;
  wire        _GEN_3197 = _GEN_1113 ? (_GEN_3196 ? (|lcam_ldq_idx_0) & _GEN_3164 : ~(_GEN_1117 & ~(|lcam_ldq_idx_0)) & _GEN_3164) : _GEN_3164;
  wire        _GEN_3198 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_296 & _GEN_3165 : ~(_GEN_1117 & _GEN_296) & _GEN_3165) : _GEN_3165;
  wire        _GEN_3199 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_297 & _GEN_3166 : ~(_GEN_1117 & _GEN_297) & _GEN_3166) : _GEN_3166;
  wire        _GEN_3200 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_298 & _GEN_3167 : ~(_GEN_1117 & _GEN_298) & _GEN_3167) : _GEN_3167;
  wire        _GEN_3201 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_299 & _GEN_3168 : ~(_GEN_1117 & _GEN_299) & _GEN_3168) : _GEN_3168;
  wire        _GEN_3202 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_300 & _GEN_3169 : ~(_GEN_1117 & _GEN_300) & _GEN_3169) : _GEN_3169;
  wire        _GEN_3203 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_301 & _GEN_3170 : ~(_GEN_1117 & _GEN_301) & _GEN_3170) : _GEN_3170;
  wire        _GEN_3204 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_302 & _GEN_3171 : ~(_GEN_1117 & _GEN_302) & _GEN_3171) : _GEN_3171;
  wire        _GEN_3205 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_303 & _GEN_3172 : ~(_GEN_1117 & _GEN_303) & _GEN_3172) : _GEN_3172;
  wire        _GEN_3206 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_304 & _GEN_3173 : ~(_GEN_1117 & _GEN_304) & _GEN_3173) : _GEN_3173;
  wire        _GEN_3207 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_305 & _GEN_3174 : ~(_GEN_1117 & _GEN_305) & _GEN_3174) : _GEN_3174;
  wire        _GEN_3208 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_306 & _GEN_3175 : ~(_GEN_1117 & _GEN_306) & _GEN_3175) : _GEN_3175;
  wire        _GEN_3209 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_307 & _GEN_3176 : ~(_GEN_1117 & _GEN_307) & _GEN_3176) : _GEN_3176;
  wire        _GEN_3210 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_308 & _GEN_3177 : ~(_GEN_1117 & _GEN_308) & _GEN_3177) : _GEN_3177;
  wire        _GEN_3211 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_309 & _GEN_3178 : ~(_GEN_1117 & _GEN_309) & _GEN_3178) : _GEN_3178;
  wire        _GEN_3212 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_310 & _GEN_3179 : ~(_GEN_1117 & _GEN_310) & _GEN_3179) : _GEN_3179;
  wire        _GEN_3213 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_311 & _GEN_3180 : ~(_GEN_1117 & _GEN_311) & _GEN_3180) : _GEN_3180;
  wire        _GEN_3214 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_312 & _GEN_3181 : ~(_GEN_1117 & _GEN_312) & _GEN_3181) : _GEN_3181;
  wire        _GEN_3215 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_313 & _GEN_3182 : ~(_GEN_1117 & _GEN_313) & _GEN_3182) : _GEN_3182;
  wire        _GEN_3216 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_314 & _GEN_3183 : ~(_GEN_1117 & _GEN_314) & _GEN_3183) : _GEN_3183;
  wire        _GEN_3217 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_315 & _GEN_3184 : ~(_GEN_1117 & _GEN_315) & _GEN_3184) : _GEN_3184;
  wire        _GEN_3218 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_316 & _GEN_3185 : ~(_GEN_1117 & _GEN_316) & _GEN_3185) : _GEN_3185;
  wire        _GEN_3219 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_317 & _GEN_3186 : ~(_GEN_1117 & _GEN_317) & _GEN_3186) : _GEN_3186;
  wire        _GEN_3220 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_318 & _GEN_3187 : ~(_GEN_1117 & _GEN_318) & _GEN_3187) : _GEN_3187;
  wire        _GEN_3221 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_319 & _GEN_3188 : ~(_GEN_1117 & _GEN_319) & _GEN_3188) : _GEN_3188;
  wire        _GEN_3222 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_320 & _GEN_3189 : ~(_GEN_1117 & _GEN_320) & _GEN_3189) : _GEN_3189;
  wire        _GEN_3223 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_321 & _GEN_3190 : ~(_GEN_1117 & _GEN_321) & _GEN_3190) : _GEN_3190;
  wire        _GEN_3224 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_322 & _GEN_3191 : ~(_GEN_1117 & _GEN_322) & _GEN_3191) : _GEN_3191;
  wire        _GEN_3225 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_323 & _GEN_3192 : ~(_GEN_1117 & _GEN_323) & _GEN_3192) : _GEN_3192;
  wire        _GEN_3226 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_324 & _GEN_3193 : ~(_GEN_1117 & _GEN_324) & _GEN_3193) : _GEN_3193;
  wire        _GEN_3227 = _GEN_1113 ? (_GEN_3196 ? ~_GEN_325 & _GEN_3194 : ~(_GEN_1117 & _GEN_325) & _GEN_3194) : _GEN_3194;
  wire        _GEN_3228 = _GEN_1113 ? (_GEN_3196 ? ~(&lcam_ldq_idx_0) & _GEN_3195 : ~(_GEN_1117 & (&lcam_ldq_idx_0)) & _GEN_3195) : _GEN_3195;
  wire        _GEN_3229 = _GEN_1121 | _GEN_1122;
  wire        _GEN_3230 = _GEN_1119 ? (_GEN_3229 ? (|lcam_ldq_idx_1) & _GEN_3197 : ~(_GEN_1117 & ~(|lcam_ldq_idx_1)) & _GEN_3197) : _GEN_3197;
  wire        _GEN_3231 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_336 & _GEN_3198 : ~(_GEN_1117 & _GEN_336) & _GEN_3198) : _GEN_3198;
  wire        _GEN_3232 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_337 & _GEN_3199 : ~(_GEN_1117 & _GEN_337) & _GEN_3199) : _GEN_3199;
  wire        _GEN_3233 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_338 & _GEN_3200 : ~(_GEN_1117 & _GEN_338) & _GEN_3200) : _GEN_3200;
  wire        _GEN_3234 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_339 & _GEN_3201 : ~(_GEN_1117 & _GEN_339) & _GEN_3201) : _GEN_3201;
  wire        _GEN_3235 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_340 & _GEN_3202 : ~(_GEN_1117 & _GEN_340) & _GEN_3202) : _GEN_3202;
  wire        _GEN_3236 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_341 & _GEN_3203 : ~(_GEN_1117 & _GEN_341) & _GEN_3203) : _GEN_3203;
  wire        _GEN_3237 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_342 & _GEN_3204 : ~(_GEN_1117 & _GEN_342) & _GEN_3204) : _GEN_3204;
  wire        _GEN_3238 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_343 & _GEN_3205 : ~(_GEN_1117 & _GEN_343) & _GEN_3205) : _GEN_3205;
  wire        _GEN_3239 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_344 & _GEN_3206 : ~(_GEN_1117 & _GEN_344) & _GEN_3206) : _GEN_3206;
  wire        _GEN_3240 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_345 & _GEN_3207 : ~(_GEN_1117 & _GEN_345) & _GEN_3207) : _GEN_3207;
  wire        _GEN_3241 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_346 & _GEN_3208 : ~(_GEN_1117 & _GEN_346) & _GEN_3208) : _GEN_3208;
  wire        _GEN_3242 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_347 & _GEN_3209 : ~(_GEN_1117 & _GEN_347) & _GEN_3209) : _GEN_3209;
  wire        _GEN_3243 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_348 & _GEN_3210 : ~(_GEN_1117 & _GEN_348) & _GEN_3210) : _GEN_3210;
  wire        _GEN_3244 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_349 & _GEN_3211 : ~(_GEN_1117 & _GEN_349) & _GEN_3211) : _GEN_3211;
  wire        _GEN_3245 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_350 & _GEN_3212 : ~(_GEN_1117 & _GEN_350) & _GEN_3212) : _GEN_3212;
  wire        _GEN_3246 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_351 & _GEN_3213 : ~(_GEN_1117 & _GEN_351) & _GEN_3213) : _GEN_3213;
  wire        _GEN_3247 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_352 & _GEN_3214 : ~(_GEN_1117 & _GEN_352) & _GEN_3214) : _GEN_3214;
  wire        _GEN_3248 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_353 & _GEN_3215 : ~(_GEN_1117 & _GEN_353) & _GEN_3215) : _GEN_3215;
  wire        _GEN_3249 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_354 & _GEN_3216 : ~(_GEN_1117 & _GEN_354) & _GEN_3216) : _GEN_3216;
  wire        _GEN_3250 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_355 & _GEN_3217 : ~(_GEN_1117 & _GEN_355) & _GEN_3217) : _GEN_3217;
  wire        _GEN_3251 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_356 & _GEN_3218 : ~(_GEN_1117 & _GEN_356) & _GEN_3218) : _GEN_3218;
  wire        _GEN_3252 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_357 & _GEN_3219 : ~(_GEN_1117 & _GEN_357) & _GEN_3219) : _GEN_3219;
  wire        _GEN_3253 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_358 & _GEN_3220 : ~(_GEN_1117 & _GEN_358) & _GEN_3220) : _GEN_3220;
  wire        _GEN_3254 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_359 & _GEN_3221 : ~(_GEN_1117 & _GEN_359) & _GEN_3221) : _GEN_3221;
  wire        _GEN_3255 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_360 & _GEN_3222 : ~(_GEN_1117 & _GEN_360) & _GEN_3222) : _GEN_3222;
  wire        _GEN_3256 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_361 & _GEN_3223 : ~(_GEN_1117 & _GEN_361) & _GEN_3223) : _GEN_3223;
  wire        _GEN_3257 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_362 & _GEN_3224 : ~(_GEN_1117 & _GEN_362) & _GEN_3224) : _GEN_3224;
  wire        _GEN_3258 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_363 & _GEN_3225 : ~(_GEN_1117 & _GEN_363) & _GEN_3225) : _GEN_3225;
  wire        _GEN_3259 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_364 & _GEN_3226 : ~(_GEN_1117 & _GEN_364) & _GEN_3226) : _GEN_3226;
  wire        _GEN_3260 = _GEN_1119 ? (_GEN_3229 ? ~_GEN_365 & _GEN_3227 : ~(_GEN_1117 & _GEN_365) & _GEN_3227) : _GEN_3227;
  wire        _GEN_3261 = _GEN_1119 ? (_GEN_3229 ? ~(&lcam_ldq_idx_1) & _GEN_3228 : ~(_GEN_1117 & (&lcam_ldq_idx_1)) & _GEN_3228) : _GEN_3228;
  wire        _GEN_3262 = _GEN_1126 | _GEN_1127;
  wire        _GEN_3263 = _GEN_1124 ? (_GEN_3262 ? (|lcam_ldq_idx_0) & _GEN_3230 : ~(_GEN_1128 & ~(|lcam_ldq_idx_0)) & _GEN_3230) : _GEN_3230;
  wire        _GEN_3264 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_296 & _GEN_3231 : ~(_GEN_1128 & _GEN_296) & _GEN_3231) : _GEN_3231;
  wire        _GEN_3265 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_297 & _GEN_3232 : ~(_GEN_1128 & _GEN_297) & _GEN_3232) : _GEN_3232;
  wire        _GEN_3266 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_298 & _GEN_3233 : ~(_GEN_1128 & _GEN_298) & _GEN_3233) : _GEN_3233;
  wire        _GEN_3267 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_299 & _GEN_3234 : ~(_GEN_1128 & _GEN_299) & _GEN_3234) : _GEN_3234;
  wire        _GEN_3268 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_300 & _GEN_3235 : ~(_GEN_1128 & _GEN_300) & _GEN_3235) : _GEN_3235;
  wire        _GEN_3269 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_301 & _GEN_3236 : ~(_GEN_1128 & _GEN_301) & _GEN_3236) : _GEN_3236;
  wire        _GEN_3270 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_302 & _GEN_3237 : ~(_GEN_1128 & _GEN_302) & _GEN_3237) : _GEN_3237;
  wire        _GEN_3271 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_303 & _GEN_3238 : ~(_GEN_1128 & _GEN_303) & _GEN_3238) : _GEN_3238;
  wire        _GEN_3272 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_304 & _GEN_3239 : ~(_GEN_1128 & _GEN_304) & _GEN_3239) : _GEN_3239;
  wire        _GEN_3273 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_305 & _GEN_3240 : ~(_GEN_1128 & _GEN_305) & _GEN_3240) : _GEN_3240;
  wire        _GEN_3274 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_306 & _GEN_3241 : ~(_GEN_1128 & _GEN_306) & _GEN_3241) : _GEN_3241;
  wire        _GEN_3275 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_307 & _GEN_3242 : ~(_GEN_1128 & _GEN_307) & _GEN_3242) : _GEN_3242;
  wire        _GEN_3276 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_308 & _GEN_3243 : ~(_GEN_1128 & _GEN_308) & _GEN_3243) : _GEN_3243;
  wire        _GEN_3277 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_309 & _GEN_3244 : ~(_GEN_1128 & _GEN_309) & _GEN_3244) : _GEN_3244;
  wire        _GEN_3278 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_310 & _GEN_3245 : ~(_GEN_1128 & _GEN_310) & _GEN_3245) : _GEN_3245;
  wire        _GEN_3279 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_311 & _GEN_3246 : ~(_GEN_1128 & _GEN_311) & _GEN_3246) : _GEN_3246;
  wire        _GEN_3280 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_312 & _GEN_3247 : ~(_GEN_1128 & _GEN_312) & _GEN_3247) : _GEN_3247;
  wire        _GEN_3281 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_313 & _GEN_3248 : ~(_GEN_1128 & _GEN_313) & _GEN_3248) : _GEN_3248;
  wire        _GEN_3282 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_314 & _GEN_3249 : ~(_GEN_1128 & _GEN_314) & _GEN_3249) : _GEN_3249;
  wire        _GEN_3283 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_315 & _GEN_3250 : ~(_GEN_1128 & _GEN_315) & _GEN_3250) : _GEN_3250;
  wire        _GEN_3284 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_316 & _GEN_3251 : ~(_GEN_1128 & _GEN_316) & _GEN_3251) : _GEN_3251;
  wire        _GEN_3285 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_317 & _GEN_3252 : ~(_GEN_1128 & _GEN_317) & _GEN_3252) : _GEN_3252;
  wire        _GEN_3286 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_318 & _GEN_3253 : ~(_GEN_1128 & _GEN_318) & _GEN_3253) : _GEN_3253;
  wire        _GEN_3287 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_319 & _GEN_3254 : ~(_GEN_1128 & _GEN_319) & _GEN_3254) : _GEN_3254;
  wire        _GEN_3288 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_320 & _GEN_3255 : ~(_GEN_1128 & _GEN_320) & _GEN_3255) : _GEN_3255;
  wire        _GEN_3289 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_321 & _GEN_3256 : ~(_GEN_1128 & _GEN_321) & _GEN_3256) : _GEN_3256;
  wire        _GEN_3290 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_322 & _GEN_3257 : ~(_GEN_1128 & _GEN_322) & _GEN_3257) : _GEN_3257;
  wire        _GEN_3291 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_323 & _GEN_3258 : ~(_GEN_1128 & _GEN_323) & _GEN_3258) : _GEN_3258;
  wire        _GEN_3292 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_324 & _GEN_3259 : ~(_GEN_1128 & _GEN_324) & _GEN_3259) : _GEN_3259;
  wire        _GEN_3293 = _GEN_1124 ? (_GEN_3262 ? ~_GEN_325 & _GEN_3260 : ~(_GEN_1128 & _GEN_325) & _GEN_3260) : _GEN_3260;
  wire        _GEN_3294 = _GEN_1124 ? (_GEN_3262 ? ~(&lcam_ldq_idx_0) & _GEN_3261 : ~(_GEN_1128 & (&lcam_ldq_idx_0)) & _GEN_3261) : _GEN_3261;
  wire        _GEN_3295 = _GEN_1132 | _GEN_1133;
  wire        _GEN_3296 = _GEN_1130 ? (_GEN_3295 ? (|lcam_ldq_idx_1) & _GEN_3263 : ~(_GEN_1128 & ~(|lcam_ldq_idx_1)) & _GEN_3263) : _GEN_3263;
  wire        _GEN_3297 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_336 & _GEN_3264 : ~(_GEN_1128 & _GEN_336) & _GEN_3264) : _GEN_3264;
  wire        _GEN_3298 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_337 & _GEN_3265 : ~(_GEN_1128 & _GEN_337) & _GEN_3265) : _GEN_3265;
  wire        _GEN_3299 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_338 & _GEN_3266 : ~(_GEN_1128 & _GEN_338) & _GEN_3266) : _GEN_3266;
  wire        _GEN_3300 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_339 & _GEN_3267 : ~(_GEN_1128 & _GEN_339) & _GEN_3267) : _GEN_3267;
  wire        _GEN_3301 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_340 & _GEN_3268 : ~(_GEN_1128 & _GEN_340) & _GEN_3268) : _GEN_3268;
  wire        _GEN_3302 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_341 & _GEN_3269 : ~(_GEN_1128 & _GEN_341) & _GEN_3269) : _GEN_3269;
  wire        _GEN_3303 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_342 & _GEN_3270 : ~(_GEN_1128 & _GEN_342) & _GEN_3270) : _GEN_3270;
  wire        _GEN_3304 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_343 & _GEN_3271 : ~(_GEN_1128 & _GEN_343) & _GEN_3271) : _GEN_3271;
  wire        _GEN_3305 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_344 & _GEN_3272 : ~(_GEN_1128 & _GEN_344) & _GEN_3272) : _GEN_3272;
  wire        _GEN_3306 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_345 & _GEN_3273 : ~(_GEN_1128 & _GEN_345) & _GEN_3273) : _GEN_3273;
  wire        _GEN_3307 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_346 & _GEN_3274 : ~(_GEN_1128 & _GEN_346) & _GEN_3274) : _GEN_3274;
  wire        _GEN_3308 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_347 & _GEN_3275 : ~(_GEN_1128 & _GEN_347) & _GEN_3275) : _GEN_3275;
  wire        _GEN_3309 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_348 & _GEN_3276 : ~(_GEN_1128 & _GEN_348) & _GEN_3276) : _GEN_3276;
  wire        _GEN_3310 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_349 & _GEN_3277 : ~(_GEN_1128 & _GEN_349) & _GEN_3277) : _GEN_3277;
  wire        _GEN_3311 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_350 & _GEN_3278 : ~(_GEN_1128 & _GEN_350) & _GEN_3278) : _GEN_3278;
  wire        _GEN_3312 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_351 & _GEN_3279 : ~(_GEN_1128 & _GEN_351) & _GEN_3279) : _GEN_3279;
  wire        _GEN_3313 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_352 & _GEN_3280 : ~(_GEN_1128 & _GEN_352) & _GEN_3280) : _GEN_3280;
  wire        _GEN_3314 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_353 & _GEN_3281 : ~(_GEN_1128 & _GEN_353) & _GEN_3281) : _GEN_3281;
  wire        _GEN_3315 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_354 & _GEN_3282 : ~(_GEN_1128 & _GEN_354) & _GEN_3282) : _GEN_3282;
  wire        _GEN_3316 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_355 & _GEN_3283 : ~(_GEN_1128 & _GEN_355) & _GEN_3283) : _GEN_3283;
  wire        _GEN_3317 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_356 & _GEN_3284 : ~(_GEN_1128 & _GEN_356) & _GEN_3284) : _GEN_3284;
  wire        _GEN_3318 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_357 & _GEN_3285 : ~(_GEN_1128 & _GEN_357) & _GEN_3285) : _GEN_3285;
  wire        _GEN_3319 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_358 & _GEN_3286 : ~(_GEN_1128 & _GEN_358) & _GEN_3286) : _GEN_3286;
  wire        _GEN_3320 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_359 & _GEN_3287 : ~(_GEN_1128 & _GEN_359) & _GEN_3287) : _GEN_3287;
  wire        _GEN_3321 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_360 & _GEN_3288 : ~(_GEN_1128 & _GEN_360) & _GEN_3288) : _GEN_3288;
  wire        _GEN_3322 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_361 & _GEN_3289 : ~(_GEN_1128 & _GEN_361) & _GEN_3289) : _GEN_3289;
  wire        _GEN_3323 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_362 & _GEN_3290 : ~(_GEN_1128 & _GEN_362) & _GEN_3290) : _GEN_3290;
  wire        _GEN_3324 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_363 & _GEN_3291 : ~(_GEN_1128 & _GEN_363) & _GEN_3291) : _GEN_3291;
  wire        _GEN_3325 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_364 & _GEN_3292 : ~(_GEN_1128 & _GEN_364) & _GEN_3292) : _GEN_3292;
  wire        _GEN_3326 = _GEN_1130 ? (_GEN_3295 ? ~_GEN_365 & _GEN_3293 : ~(_GEN_1128 & _GEN_365) & _GEN_3293) : _GEN_3293;
  wire        _GEN_3327 = _GEN_1130 ? (_GEN_3295 ? ~(&lcam_ldq_idx_1) & _GEN_3294 : ~(_GEN_1128 & (&lcam_ldq_idx_1)) & _GEN_3294) : _GEN_3294;
  wire        _GEN_3328 = _GEN_1137 | _GEN_1138;
  wire        _GEN_3329 = _GEN_1135 ? (_GEN_3328 ? (|lcam_ldq_idx_0) & _GEN_3296 : ~(_GEN_1139 & ~(|lcam_ldq_idx_0)) & _GEN_3296) : _GEN_3296;
  wire        _GEN_3330 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_296 & _GEN_3297 : ~(_GEN_1139 & _GEN_296) & _GEN_3297) : _GEN_3297;
  wire        _GEN_3331 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_297 & _GEN_3298 : ~(_GEN_1139 & _GEN_297) & _GEN_3298) : _GEN_3298;
  wire        _GEN_3332 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_298 & _GEN_3299 : ~(_GEN_1139 & _GEN_298) & _GEN_3299) : _GEN_3299;
  wire        _GEN_3333 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_299 & _GEN_3300 : ~(_GEN_1139 & _GEN_299) & _GEN_3300) : _GEN_3300;
  wire        _GEN_3334 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_300 & _GEN_3301 : ~(_GEN_1139 & _GEN_300) & _GEN_3301) : _GEN_3301;
  wire        _GEN_3335 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_301 & _GEN_3302 : ~(_GEN_1139 & _GEN_301) & _GEN_3302) : _GEN_3302;
  wire        _GEN_3336 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_302 & _GEN_3303 : ~(_GEN_1139 & _GEN_302) & _GEN_3303) : _GEN_3303;
  wire        _GEN_3337 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_303 & _GEN_3304 : ~(_GEN_1139 & _GEN_303) & _GEN_3304) : _GEN_3304;
  wire        _GEN_3338 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_304 & _GEN_3305 : ~(_GEN_1139 & _GEN_304) & _GEN_3305) : _GEN_3305;
  wire        _GEN_3339 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_305 & _GEN_3306 : ~(_GEN_1139 & _GEN_305) & _GEN_3306) : _GEN_3306;
  wire        _GEN_3340 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_306 & _GEN_3307 : ~(_GEN_1139 & _GEN_306) & _GEN_3307) : _GEN_3307;
  wire        _GEN_3341 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_307 & _GEN_3308 : ~(_GEN_1139 & _GEN_307) & _GEN_3308) : _GEN_3308;
  wire        _GEN_3342 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_308 & _GEN_3309 : ~(_GEN_1139 & _GEN_308) & _GEN_3309) : _GEN_3309;
  wire        _GEN_3343 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_309 & _GEN_3310 : ~(_GEN_1139 & _GEN_309) & _GEN_3310) : _GEN_3310;
  wire        _GEN_3344 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_310 & _GEN_3311 : ~(_GEN_1139 & _GEN_310) & _GEN_3311) : _GEN_3311;
  wire        _GEN_3345 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_311 & _GEN_3312 : ~(_GEN_1139 & _GEN_311) & _GEN_3312) : _GEN_3312;
  wire        _GEN_3346 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_312 & _GEN_3313 : ~(_GEN_1139 & _GEN_312) & _GEN_3313) : _GEN_3313;
  wire        _GEN_3347 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_313 & _GEN_3314 : ~(_GEN_1139 & _GEN_313) & _GEN_3314) : _GEN_3314;
  wire        _GEN_3348 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_314 & _GEN_3315 : ~(_GEN_1139 & _GEN_314) & _GEN_3315) : _GEN_3315;
  wire        _GEN_3349 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_315 & _GEN_3316 : ~(_GEN_1139 & _GEN_315) & _GEN_3316) : _GEN_3316;
  wire        _GEN_3350 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_316 & _GEN_3317 : ~(_GEN_1139 & _GEN_316) & _GEN_3317) : _GEN_3317;
  wire        _GEN_3351 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_317 & _GEN_3318 : ~(_GEN_1139 & _GEN_317) & _GEN_3318) : _GEN_3318;
  wire        _GEN_3352 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_318 & _GEN_3319 : ~(_GEN_1139 & _GEN_318) & _GEN_3319) : _GEN_3319;
  wire        _GEN_3353 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_319 & _GEN_3320 : ~(_GEN_1139 & _GEN_319) & _GEN_3320) : _GEN_3320;
  wire        _GEN_3354 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_320 & _GEN_3321 : ~(_GEN_1139 & _GEN_320) & _GEN_3321) : _GEN_3321;
  wire        _GEN_3355 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_321 & _GEN_3322 : ~(_GEN_1139 & _GEN_321) & _GEN_3322) : _GEN_3322;
  wire        _GEN_3356 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_322 & _GEN_3323 : ~(_GEN_1139 & _GEN_322) & _GEN_3323) : _GEN_3323;
  wire        _GEN_3357 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_323 & _GEN_3324 : ~(_GEN_1139 & _GEN_323) & _GEN_3324) : _GEN_3324;
  wire        _GEN_3358 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_324 & _GEN_3325 : ~(_GEN_1139 & _GEN_324) & _GEN_3325) : _GEN_3325;
  wire        _GEN_3359 = _GEN_1135 ? (_GEN_3328 ? ~_GEN_325 & _GEN_3326 : ~(_GEN_1139 & _GEN_325) & _GEN_3326) : _GEN_3326;
  wire        _GEN_3360 = _GEN_1135 ? (_GEN_3328 ? ~(&lcam_ldq_idx_0) & _GEN_3327 : ~(_GEN_1139 & (&lcam_ldq_idx_0)) & _GEN_3327) : _GEN_3327;
  wire        _GEN_3361 = _GEN_1143 | _GEN_1144;
  wire        _GEN_3362 = _GEN_1141 ? (_GEN_3361 ? (|lcam_ldq_idx_1) & _GEN_3329 : ~(_GEN_1139 & ~(|lcam_ldq_idx_1)) & _GEN_3329) : _GEN_3329;
  wire        _GEN_3363 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_336 & _GEN_3330 : ~(_GEN_1139 & _GEN_336) & _GEN_3330) : _GEN_3330;
  wire        _GEN_3364 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_337 & _GEN_3331 : ~(_GEN_1139 & _GEN_337) & _GEN_3331) : _GEN_3331;
  wire        _GEN_3365 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_338 & _GEN_3332 : ~(_GEN_1139 & _GEN_338) & _GEN_3332) : _GEN_3332;
  wire        _GEN_3366 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_339 & _GEN_3333 : ~(_GEN_1139 & _GEN_339) & _GEN_3333) : _GEN_3333;
  wire        _GEN_3367 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_340 & _GEN_3334 : ~(_GEN_1139 & _GEN_340) & _GEN_3334) : _GEN_3334;
  wire        _GEN_3368 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_341 & _GEN_3335 : ~(_GEN_1139 & _GEN_341) & _GEN_3335) : _GEN_3335;
  wire        _GEN_3369 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_342 & _GEN_3336 : ~(_GEN_1139 & _GEN_342) & _GEN_3336) : _GEN_3336;
  wire        _GEN_3370 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_343 & _GEN_3337 : ~(_GEN_1139 & _GEN_343) & _GEN_3337) : _GEN_3337;
  wire        _GEN_3371 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_344 & _GEN_3338 : ~(_GEN_1139 & _GEN_344) & _GEN_3338) : _GEN_3338;
  wire        _GEN_3372 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_345 & _GEN_3339 : ~(_GEN_1139 & _GEN_345) & _GEN_3339) : _GEN_3339;
  wire        _GEN_3373 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_346 & _GEN_3340 : ~(_GEN_1139 & _GEN_346) & _GEN_3340) : _GEN_3340;
  wire        _GEN_3374 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_347 & _GEN_3341 : ~(_GEN_1139 & _GEN_347) & _GEN_3341) : _GEN_3341;
  wire        _GEN_3375 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_348 & _GEN_3342 : ~(_GEN_1139 & _GEN_348) & _GEN_3342) : _GEN_3342;
  wire        _GEN_3376 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_349 & _GEN_3343 : ~(_GEN_1139 & _GEN_349) & _GEN_3343) : _GEN_3343;
  wire        _GEN_3377 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_350 & _GEN_3344 : ~(_GEN_1139 & _GEN_350) & _GEN_3344) : _GEN_3344;
  wire        _GEN_3378 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_351 & _GEN_3345 : ~(_GEN_1139 & _GEN_351) & _GEN_3345) : _GEN_3345;
  wire        _GEN_3379 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_352 & _GEN_3346 : ~(_GEN_1139 & _GEN_352) & _GEN_3346) : _GEN_3346;
  wire        _GEN_3380 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_353 & _GEN_3347 : ~(_GEN_1139 & _GEN_353) & _GEN_3347) : _GEN_3347;
  wire        _GEN_3381 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_354 & _GEN_3348 : ~(_GEN_1139 & _GEN_354) & _GEN_3348) : _GEN_3348;
  wire        _GEN_3382 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_355 & _GEN_3349 : ~(_GEN_1139 & _GEN_355) & _GEN_3349) : _GEN_3349;
  wire        _GEN_3383 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_356 & _GEN_3350 : ~(_GEN_1139 & _GEN_356) & _GEN_3350) : _GEN_3350;
  wire        _GEN_3384 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_357 & _GEN_3351 : ~(_GEN_1139 & _GEN_357) & _GEN_3351) : _GEN_3351;
  wire        _GEN_3385 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_358 & _GEN_3352 : ~(_GEN_1139 & _GEN_358) & _GEN_3352) : _GEN_3352;
  wire        _GEN_3386 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_359 & _GEN_3353 : ~(_GEN_1139 & _GEN_359) & _GEN_3353) : _GEN_3353;
  wire        _GEN_3387 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_360 & _GEN_3354 : ~(_GEN_1139 & _GEN_360) & _GEN_3354) : _GEN_3354;
  wire        _GEN_3388 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_361 & _GEN_3355 : ~(_GEN_1139 & _GEN_361) & _GEN_3355) : _GEN_3355;
  wire        _GEN_3389 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_362 & _GEN_3356 : ~(_GEN_1139 & _GEN_362) & _GEN_3356) : _GEN_3356;
  wire        _GEN_3390 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_363 & _GEN_3357 : ~(_GEN_1139 & _GEN_363) & _GEN_3357) : _GEN_3357;
  wire        _GEN_3391 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_364 & _GEN_3358 : ~(_GEN_1139 & _GEN_364) & _GEN_3358) : _GEN_3358;
  wire        _GEN_3392 = _GEN_1141 ? (_GEN_3361 ? ~_GEN_365 & _GEN_3359 : ~(_GEN_1139 & _GEN_365) & _GEN_3359) : _GEN_3359;
  wire        _GEN_3393 = _GEN_1141 ? (_GEN_3361 ? ~(&lcam_ldq_idx_1) & _GEN_3360 : ~(_GEN_1139 & (&lcam_ldq_idx_1)) & _GEN_3360) : _GEN_3360;
  wire        _GEN_3394 = _GEN_1148 | _GEN_1149;
  wire        _GEN_3395 = _GEN_1146 ? (_GEN_3394 ? (|lcam_ldq_idx_0) & _GEN_3362 : ~(_GEN_1150 & ~(|lcam_ldq_idx_0)) & _GEN_3362) : _GEN_3362;
  wire        _GEN_3396 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_296 & _GEN_3363 : ~(_GEN_1150 & _GEN_296) & _GEN_3363) : _GEN_3363;
  wire        _GEN_3397 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_297 & _GEN_3364 : ~(_GEN_1150 & _GEN_297) & _GEN_3364) : _GEN_3364;
  wire        _GEN_3398 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_298 & _GEN_3365 : ~(_GEN_1150 & _GEN_298) & _GEN_3365) : _GEN_3365;
  wire        _GEN_3399 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_299 & _GEN_3366 : ~(_GEN_1150 & _GEN_299) & _GEN_3366) : _GEN_3366;
  wire        _GEN_3400 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_300 & _GEN_3367 : ~(_GEN_1150 & _GEN_300) & _GEN_3367) : _GEN_3367;
  wire        _GEN_3401 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_301 & _GEN_3368 : ~(_GEN_1150 & _GEN_301) & _GEN_3368) : _GEN_3368;
  wire        _GEN_3402 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_302 & _GEN_3369 : ~(_GEN_1150 & _GEN_302) & _GEN_3369) : _GEN_3369;
  wire        _GEN_3403 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_303 & _GEN_3370 : ~(_GEN_1150 & _GEN_303) & _GEN_3370) : _GEN_3370;
  wire        _GEN_3404 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_304 & _GEN_3371 : ~(_GEN_1150 & _GEN_304) & _GEN_3371) : _GEN_3371;
  wire        _GEN_3405 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_305 & _GEN_3372 : ~(_GEN_1150 & _GEN_305) & _GEN_3372) : _GEN_3372;
  wire        _GEN_3406 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_306 & _GEN_3373 : ~(_GEN_1150 & _GEN_306) & _GEN_3373) : _GEN_3373;
  wire        _GEN_3407 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_307 & _GEN_3374 : ~(_GEN_1150 & _GEN_307) & _GEN_3374) : _GEN_3374;
  wire        _GEN_3408 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_308 & _GEN_3375 : ~(_GEN_1150 & _GEN_308) & _GEN_3375) : _GEN_3375;
  wire        _GEN_3409 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_309 & _GEN_3376 : ~(_GEN_1150 & _GEN_309) & _GEN_3376) : _GEN_3376;
  wire        _GEN_3410 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_310 & _GEN_3377 : ~(_GEN_1150 & _GEN_310) & _GEN_3377) : _GEN_3377;
  wire        _GEN_3411 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_311 & _GEN_3378 : ~(_GEN_1150 & _GEN_311) & _GEN_3378) : _GEN_3378;
  wire        _GEN_3412 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_312 & _GEN_3379 : ~(_GEN_1150 & _GEN_312) & _GEN_3379) : _GEN_3379;
  wire        _GEN_3413 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_313 & _GEN_3380 : ~(_GEN_1150 & _GEN_313) & _GEN_3380) : _GEN_3380;
  wire        _GEN_3414 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_314 & _GEN_3381 : ~(_GEN_1150 & _GEN_314) & _GEN_3381) : _GEN_3381;
  wire        _GEN_3415 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_315 & _GEN_3382 : ~(_GEN_1150 & _GEN_315) & _GEN_3382) : _GEN_3382;
  wire        _GEN_3416 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_316 & _GEN_3383 : ~(_GEN_1150 & _GEN_316) & _GEN_3383) : _GEN_3383;
  wire        _GEN_3417 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_317 & _GEN_3384 : ~(_GEN_1150 & _GEN_317) & _GEN_3384) : _GEN_3384;
  wire        _GEN_3418 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_318 & _GEN_3385 : ~(_GEN_1150 & _GEN_318) & _GEN_3385) : _GEN_3385;
  wire        _GEN_3419 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_319 & _GEN_3386 : ~(_GEN_1150 & _GEN_319) & _GEN_3386) : _GEN_3386;
  wire        _GEN_3420 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_320 & _GEN_3387 : ~(_GEN_1150 & _GEN_320) & _GEN_3387) : _GEN_3387;
  wire        _GEN_3421 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_321 & _GEN_3388 : ~(_GEN_1150 & _GEN_321) & _GEN_3388) : _GEN_3388;
  wire        _GEN_3422 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_322 & _GEN_3389 : ~(_GEN_1150 & _GEN_322) & _GEN_3389) : _GEN_3389;
  wire        _GEN_3423 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_323 & _GEN_3390 : ~(_GEN_1150 & _GEN_323) & _GEN_3390) : _GEN_3390;
  wire        _GEN_3424 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_324 & _GEN_3391 : ~(_GEN_1150 & _GEN_324) & _GEN_3391) : _GEN_3391;
  wire        _GEN_3425 = _GEN_1146 ? (_GEN_3394 ? ~_GEN_325 & _GEN_3392 : ~(_GEN_1150 & _GEN_325) & _GEN_3392) : _GEN_3392;
  wire        _GEN_3426 = _GEN_1146 ? (_GEN_3394 ? ~(&lcam_ldq_idx_0) & _GEN_3393 : ~(_GEN_1150 & (&lcam_ldq_idx_0)) & _GEN_3393) : _GEN_3393;
  wire        _GEN_3427 = _GEN_1154 | _GEN_1155;
  wire        _GEN_3428 = _GEN_1152 ? (_GEN_3427 ? (|lcam_ldq_idx_1) & _GEN_3395 : ~(_GEN_1150 & ~(|lcam_ldq_idx_1)) & _GEN_3395) : _GEN_3395;
  wire        _GEN_3429 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_336 & _GEN_3396 : ~(_GEN_1150 & _GEN_336) & _GEN_3396) : _GEN_3396;
  wire        _GEN_3430 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_337 & _GEN_3397 : ~(_GEN_1150 & _GEN_337) & _GEN_3397) : _GEN_3397;
  wire        _GEN_3431 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_338 & _GEN_3398 : ~(_GEN_1150 & _GEN_338) & _GEN_3398) : _GEN_3398;
  wire        _GEN_3432 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_339 & _GEN_3399 : ~(_GEN_1150 & _GEN_339) & _GEN_3399) : _GEN_3399;
  wire        _GEN_3433 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_340 & _GEN_3400 : ~(_GEN_1150 & _GEN_340) & _GEN_3400) : _GEN_3400;
  wire        _GEN_3434 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_341 & _GEN_3401 : ~(_GEN_1150 & _GEN_341) & _GEN_3401) : _GEN_3401;
  wire        _GEN_3435 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_342 & _GEN_3402 : ~(_GEN_1150 & _GEN_342) & _GEN_3402) : _GEN_3402;
  wire        _GEN_3436 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_343 & _GEN_3403 : ~(_GEN_1150 & _GEN_343) & _GEN_3403) : _GEN_3403;
  wire        _GEN_3437 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_344 & _GEN_3404 : ~(_GEN_1150 & _GEN_344) & _GEN_3404) : _GEN_3404;
  wire        _GEN_3438 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_345 & _GEN_3405 : ~(_GEN_1150 & _GEN_345) & _GEN_3405) : _GEN_3405;
  wire        _GEN_3439 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_346 & _GEN_3406 : ~(_GEN_1150 & _GEN_346) & _GEN_3406) : _GEN_3406;
  wire        _GEN_3440 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_347 & _GEN_3407 : ~(_GEN_1150 & _GEN_347) & _GEN_3407) : _GEN_3407;
  wire        _GEN_3441 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_348 & _GEN_3408 : ~(_GEN_1150 & _GEN_348) & _GEN_3408) : _GEN_3408;
  wire        _GEN_3442 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_349 & _GEN_3409 : ~(_GEN_1150 & _GEN_349) & _GEN_3409) : _GEN_3409;
  wire        _GEN_3443 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_350 & _GEN_3410 : ~(_GEN_1150 & _GEN_350) & _GEN_3410) : _GEN_3410;
  wire        _GEN_3444 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_351 & _GEN_3411 : ~(_GEN_1150 & _GEN_351) & _GEN_3411) : _GEN_3411;
  wire        _GEN_3445 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_352 & _GEN_3412 : ~(_GEN_1150 & _GEN_352) & _GEN_3412) : _GEN_3412;
  wire        _GEN_3446 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_353 & _GEN_3413 : ~(_GEN_1150 & _GEN_353) & _GEN_3413) : _GEN_3413;
  wire        _GEN_3447 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_354 & _GEN_3414 : ~(_GEN_1150 & _GEN_354) & _GEN_3414) : _GEN_3414;
  wire        _GEN_3448 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_355 & _GEN_3415 : ~(_GEN_1150 & _GEN_355) & _GEN_3415) : _GEN_3415;
  wire        _GEN_3449 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_356 & _GEN_3416 : ~(_GEN_1150 & _GEN_356) & _GEN_3416) : _GEN_3416;
  wire        _GEN_3450 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_357 & _GEN_3417 : ~(_GEN_1150 & _GEN_357) & _GEN_3417) : _GEN_3417;
  wire        _GEN_3451 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_358 & _GEN_3418 : ~(_GEN_1150 & _GEN_358) & _GEN_3418) : _GEN_3418;
  wire        _GEN_3452 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_359 & _GEN_3419 : ~(_GEN_1150 & _GEN_359) & _GEN_3419) : _GEN_3419;
  wire        _GEN_3453 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_360 & _GEN_3420 : ~(_GEN_1150 & _GEN_360) & _GEN_3420) : _GEN_3420;
  wire        _GEN_3454 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_361 & _GEN_3421 : ~(_GEN_1150 & _GEN_361) & _GEN_3421) : _GEN_3421;
  wire        _GEN_3455 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_362 & _GEN_3422 : ~(_GEN_1150 & _GEN_362) & _GEN_3422) : _GEN_3422;
  wire        _GEN_3456 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_363 & _GEN_3423 : ~(_GEN_1150 & _GEN_363) & _GEN_3423) : _GEN_3423;
  wire        _GEN_3457 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_364 & _GEN_3424 : ~(_GEN_1150 & _GEN_364) & _GEN_3424) : _GEN_3424;
  wire        _GEN_3458 = _GEN_1152 ? (_GEN_3427 ? ~_GEN_365 & _GEN_3425 : ~(_GEN_1150 & _GEN_365) & _GEN_3425) : _GEN_3425;
  wire        _GEN_3459 = _GEN_1152 ? (_GEN_3427 ? ~(&lcam_ldq_idx_1) & _GEN_3426 : ~(_GEN_1150 & (&lcam_ldq_idx_1)) & _GEN_3426) : _GEN_3426;
  wire        _GEN_3460 = _GEN_1159 | _GEN_1160;
  wire        _GEN_3461 = _GEN_1157 ? (_GEN_3460 ? (|lcam_ldq_idx_0) & _GEN_3428 : ~(_GEN_1161 & ~(|lcam_ldq_idx_0)) & _GEN_3428) : _GEN_3428;
  wire        _GEN_3462 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_296 & _GEN_3429 : ~(_GEN_1161 & _GEN_296) & _GEN_3429) : _GEN_3429;
  wire        _GEN_3463 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_297 & _GEN_3430 : ~(_GEN_1161 & _GEN_297) & _GEN_3430) : _GEN_3430;
  wire        _GEN_3464 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_298 & _GEN_3431 : ~(_GEN_1161 & _GEN_298) & _GEN_3431) : _GEN_3431;
  wire        _GEN_3465 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_299 & _GEN_3432 : ~(_GEN_1161 & _GEN_299) & _GEN_3432) : _GEN_3432;
  wire        _GEN_3466 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_300 & _GEN_3433 : ~(_GEN_1161 & _GEN_300) & _GEN_3433) : _GEN_3433;
  wire        _GEN_3467 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_301 & _GEN_3434 : ~(_GEN_1161 & _GEN_301) & _GEN_3434) : _GEN_3434;
  wire        _GEN_3468 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_302 & _GEN_3435 : ~(_GEN_1161 & _GEN_302) & _GEN_3435) : _GEN_3435;
  wire        _GEN_3469 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_303 & _GEN_3436 : ~(_GEN_1161 & _GEN_303) & _GEN_3436) : _GEN_3436;
  wire        _GEN_3470 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_304 & _GEN_3437 : ~(_GEN_1161 & _GEN_304) & _GEN_3437) : _GEN_3437;
  wire        _GEN_3471 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_305 & _GEN_3438 : ~(_GEN_1161 & _GEN_305) & _GEN_3438) : _GEN_3438;
  wire        _GEN_3472 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_306 & _GEN_3439 : ~(_GEN_1161 & _GEN_306) & _GEN_3439) : _GEN_3439;
  wire        _GEN_3473 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_307 & _GEN_3440 : ~(_GEN_1161 & _GEN_307) & _GEN_3440) : _GEN_3440;
  wire        _GEN_3474 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_308 & _GEN_3441 : ~(_GEN_1161 & _GEN_308) & _GEN_3441) : _GEN_3441;
  wire        _GEN_3475 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_309 & _GEN_3442 : ~(_GEN_1161 & _GEN_309) & _GEN_3442) : _GEN_3442;
  wire        _GEN_3476 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_310 & _GEN_3443 : ~(_GEN_1161 & _GEN_310) & _GEN_3443) : _GEN_3443;
  wire        _GEN_3477 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_311 & _GEN_3444 : ~(_GEN_1161 & _GEN_311) & _GEN_3444) : _GEN_3444;
  wire        _GEN_3478 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_312 & _GEN_3445 : ~(_GEN_1161 & _GEN_312) & _GEN_3445) : _GEN_3445;
  wire        _GEN_3479 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_313 & _GEN_3446 : ~(_GEN_1161 & _GEN_313) & _GEN_3446) : _GEN_3446;
  wire        _GEN_3480 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_314 & _GEN_3447 : ~(_GEN_1161 & _GEN_314) & _GEN_3447) : _GEN_3447;
  wire        _GEN_3481 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_315 & _GEN_3448 : ~(_GEN_1161 & _GEN_315) & _GEN_3448) : _GEN_3448;
  wire        _GEN_3482 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_316 & _GEN_3449 : ~(_GEN_1161 & _GEN_316) & _GEN_3449) : _GEN_3449;
  wire        _GEN_3483 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_317 & _GEN_3450 : ~(_GEN_1161 & _GEN_317) & _GEN_3450) : _GEN_3450;
  wire        _GEN_3484 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_318 & _GEN_3451 : ~(_GEN_1161 & _GEN_318) & _GEN_3451) : _GEN_3451;
  wire        _GEN_3485 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_319 & _GEN_3452 : ~(_GEN_1161 & _GEN_319) & _GEN_3452) : _GEN_3452;
  wire        _GEN_3486 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_320 & _GEN_3453 : ~(_GEN_1161 & _GEN_320) & _GEN_3453) : _GEN_3453;
  wire        _GEN_3487 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_321 & _GEN_3454 : ~(_GEN_1161 & _GEN_321) & _GEN_3454) : _GEN_3454;
  wire        _GEN_3488 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_322 & _GEN_3455 : ~(_GEN_1161 & _GEN_322) & _GEN_3455) : _GEN_3455;
  wire        _GEN_3489 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_323 & _GEN_3456 : ~(_GEN_1161 & _GEN_323) & _GEN_3456) : _GEN_3456;
  wire        _GEN_3490 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_324 & _GEN_3457 : ~(_GEN_1161 & _GEN_324) & _GEN_3457) : _GEN_3457;
  wire        _GEN_3491 = _GEN_1157 ? (_GEN_3460 ? ~_GEN_325 & _GEN_3458 : ~(_GEN_1161 & _GEN_325) & _GEN_3458) : _GEN_3458;
  wire        _GEN_3492 = _GEN_1157 ? (_GEN_3460 ? ~(&lcam_ldq_idx_0) & _GEN_3459 : ~(_GEN_1161 & (&lcam_ldq_idx_0)) & _GEN_3459) : _GEN_3459;
  wire        _GEN_3493 = _GEN_1165 | _GEN_1166;
  wire        _GEN_3494 = _GEN_1163 ? (_GEN_3493 ? (|lcam_ldq_idx_1) & _GEN_3461 : ~(_GEN_1161 & ~(|lcam_ldq_idx_1)) & _GEN_3461) : _GEN_3461;
  wire        _GEN_3495 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_336 & _GEN_3462 : ~(_GEN_1161 & _GEN_336) & _GEN_3462) : _GEN_3462;
  wire        _GEN_3496 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_337 & _GEN_3463 : ~(_GEN_1161 & _GEN_337) & _GEN_3463) : _GEN_3463;
  wire        _GEN_3497 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_338 & _GEN_3464 : ~(_GEN_1161 & _GEN_338) & _GEN_3464) : _GEN_3464;
  wire        _GEN_3498 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_339 & _GEN_3465 : ~(_GEN_1161 & _GEN_339) & _GEN_3465) : _GEN_3465;
  wire        _GEN_3499 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_340 & _GEN_3466 : ~(_GEN_1161 & _GEN_340) & _GEN_3466) : _GEN_3466;
  wire        _GEN_3500 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_341 & _GEN_3467 : ~(_GEN_1161 & _GEN_341) & _GEN_3467) : _GEN_3467;
  wire        _GEN_3501 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_342 & _GEN_3468 : ~(_GEN_1161 & _GEN_342) & _GEN_3468) : _GEN_3468;
  wire        _GEN_3502 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_343 & _GEN_3469 : ~(_GEN_1161 & _GEN_343) & _GEN_3469) : _GEN_3469;
  wire        _GEN_3503 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_344 & _GEN_3470 : ~(_GEN_1161 & _GEN_344) & _GEN_3470) : _GEN_3470;
  wire        _GEN_3504 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_345 & _GEN_3471 : ~(_GEN_1161 & _GEN_345) & _GEN_3471) : _GEN_3471;
  wire        _GEN_3505 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_346 & _GEN_3472 : ~(_GEN_1161 & _GEN_346) & _GEN_3472) : _GEN_3472;
  wire        _GEN_3506 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_347 & _GEN_3473 : ~(_GEN_1161 & _GEN_347) & _GEN_3473) : _GEN_3473;
  wire        _GEN_3507 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_348 & _GEN_3474 : ~(_GEN_1161 & _GEN_348) & _GEN_3474) : _GEN_3474;
  wire        _GEN_3508 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_349 & _GEN_3475 : ~(_GEN_1161 & _GEN_349) & _GEN_3475) : _GEN_3475;
  wire        _GEN_3509 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_350 & _GEN_3476 : ~(_GEN_1161 & _GEN_350) & _GEN_3476) : _GEN_3476;
  wire        _GEN_3510 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_351 & _GEN_3477 : ~(_GEN_1161 & _GEN_351) & _GEN_3477) : _GEN_3477;
  wire        _GEN_3511 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_352 & _GEN_3478 : ~(_GEN_1161 & _GEN_352) & _GEN_3478) : _GEN_3478;
  wire        _GEN_3512 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_353 & _GEN_3479 : ~(_GEN_1161 & _GEN_353) & _GEN_3479) : _GEN_3479;
  wire        _GEN_3513 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_354 & _GEN_3480 : ~(_GEN_1161 & _GEN_354) & _GEN_3480) : _GEN_3480;
  wire        _GEN_3514 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_355 & _GEN_3481 : ~(_GEN_1161 & _GEN_355) & _GEN_3481) : _GEN_3481;
  wire        _GEN_3515 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_356 & _GEN_3482 : ~(_GEN_1161 & _GEN_356) & _GEN_3482) : _GEN_3482;
  wire        _GEN_3516 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_357 & _GEN_3483 : ~(_GEN_1161 & _GEN_357) & _GEN_3483) : _GEN_3483;
  wire        _GEN_3517 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_358 & _GEN_3484 : ~(_GEN_1161 & _GEN_358) & _GEN_3484) : _GEN_3484;
  wire        _GEN_3518 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_359 & _GEN_3485 : ~(_GEN_1161 & _GEN_359) & _GEN_3485) : _GEN_3485;
  wire        _GEN_3519 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_360 & _GEN_3486 : ~(_GEN_1161 & _GEN_360) & _GEN_3486) : _GEN_3486;
  wire        _GEN_3520 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_361 & _GEN_3487 : ~(_GEN_1161 & _GEN_361) & _GEN_3487) : _GEN_3487;
  wire        _GEN_3521 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_362 & _GEN_3488 : ~(_GEN_1161 & _GEN_362) & _GEN_3488) : _GEN_3488;
  wire        _GEN_3522 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_363 & _GEN_3489 : ~(_GEN_1161 & _GEN_363) & _GEN_3489) : _GEN_3489;
  wire        _GEN_3523 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_364 & _GEN_3490 : ~(_GEN_1161 & _GEN_364) & _GEN_3490) : _GEN_3490;
  wire        _GEN_3524 = _GEN_1163 ? (_GEN_3493 ? ~_GEN_365 & _GEN_3491 : ~(_GEN_1161 & _GEN_365) & _GEN_3491) : _GEN_3491;
  wire        _GEN_3525 = _GEN_1163 ? (_GEN_3493 ? ~(&lcam_ldq_idx_1) & _GEN_3492 : ~(_GEN_1161 & (&lcam_ldq_idx_1)) & _GEN_3492) : _GEN_3492;
  wire        _GEN_3526 = _GEN_1170 | _GEN_1171;
  wire        _GEN_3527 = _GEN_1168 ? (_GEN_3526 ? (|lcam_ldq_idx_0) & _GEN_3494 : ~(_GEN_1172 & ~(|lcam_ldq_idx_0)) & _GEN_3494) : _GEN_3494;
  wire        _GEN_3528 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_296 & _GEN_3495 : ~(_GEN_1172 & _GEN_296) & _GEN_3495) : _GEN_3495;
  wire        _GEN_3529 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_297 & _GEN_3496 : ~(_GEN_1172 & _GEN_297) & _GEN_3496) : _GEN_3496;
  wire        _GEN_3530 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_298 & _GEN_3497 : ~(_GEN_1172 & _GEN_298) & _GEN_3497) : _GEN_3497;
  wire        _GEN_3531 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_299 & _GEN_3498 : ~(_GEN_1172 & _GEN_299) & _GEN_3498) : _GEN_3498;
  wire        _GEN_3532 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_300 & _GEN_3499 : ~(_GEN_1172 & _GEN_300) & _GEN_3499) : _GEN_3499;
  wire        _GEN_3533 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_301 & _GEN_3500 : ~(_GEN_1172 & _GEN_301) & _GEN_3500) : _GEN_3500;
  wire        _GEN_3534 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_302 & _GEN_3501 : ~(_GEN_1172 & _GEN_302) & _GEN_3501) : _GEN_3501;
  wire        _GEN_3535 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_303 & _GEN_3502 : ~(_GEN_1172 & _GEN_303) & _GEN_3502) : _GEN_3502;
  wire        _GEN_3536 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_304 & _GEN_3503 : ~(_GEN_1172 & _GEN_304) & _GEN_3503) : _GEN_3503;
  wire        _GEN_3537 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_305 & _GEN_3504 : ~(_GEN_1172 & _GEN_305) & _GEN_3504) : _GEN_3504;
  wire        _GEN_3538 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_306 & _GEN_3505 : ~(_GEN_1172 & _GEN_306) & _GEN_3505) : _GEN_3505;
  wire        _GEN_3539 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_307 & _GEN_3506 : ~(_GEN_1172 & _GEN_307) & _GEN_3506) : _GEN_3506;
  wire        _GEN_3540 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_308 & _GEN_3507 : ~(_GEN_1172 & _GEN_308) & _GEN_3507) : _GEN_3507;
  wire        _GEN_3541 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_309 & _GEN_3508 : ~(_GEN_1172 & _GEN_309) & _GEN_3508) : _GEN_3508;
  wire        _GEN_3542 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_310 & _GEN_3509 : ~(_GEN_1172 & _GEN_310) & _GEN_3509) : _GEN_3509;
  wire        _GEN_3543 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_311 & _GEN_3510 : ~(_GEN_1172 & _GEN_311) & _GEN_3510) : _GEN_3510;
  wire        _GEN_3544 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_312 & _GEN_3511 : ~(_GEN_1172 & _GEN_312) & _GEN_3511) : _GEN_3511;
  wire        _GEN_3545 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_313 & _GEN_3512 : ~(_GEN_1172 & _GEN_313) & _GEN_3512) : _GEN_3512;
  wire        _GEN_3546 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_314 & _GEN_3513 : ~(_GEN_1172 & _GEN_314) & _GEN_3513) : _GEN_3513;
  wire        _GEN_3547 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_315 & _GEN_3514 : ~(_GEN_1172 & _GEN_315) & _GEN_3514) : _GEN_3514;
  wire        _GEN_3548 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_316 & _GEN_3515 : ~(_GEN_1172 & _GEN_316) & _GEN_3515) : _GEN_3515;
  wire        _GEN_3549 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_317 & _GEN_3516 : ~(_GEN_1172 & _GEN_317) & _GEN_3516) : _GEN_3516;
  wire        _GEN_3550 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_318 & _GEN_3517 : ~(_GEN_1172 & _GEN_318) & _GEN_3517) : _GEN_3517;
  wire        _GEN_3551 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_319 & _GEN_3518 : ~(_GEN_1172 & _GEN_319) & _GEN_3518) : _GEN_3518;
  wire        _GEN_3552 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_320 & _GEN_3519 : ~(_GEN_1172 & _GEN_320) & _GEN_3519) : _GEN_3519;
  wire        _GEN_3553 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_321 & _GEN_3520 : ~(_GEN_1172 & _GEN_321) & _GEN_3520) : _GEN_3520;
  wire        _GEN_3554 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_322 & _GEN_3521 : ~(_GEN_1172 & _GEN_322) & _GEN_3521) : _GEN_3521;
  wire        _GEN_3555 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_323 & _GEN_3522 : ~(_GEN_1172 & _GEN_323) & _GEN_3522) : _GEN_3522;
  wire        _GEN_3556 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_324 & _GEN_3523 : ~(_GEN_1172 & _GEN_324) & _GEN_3523) : _GEN_3523;
  wire        _GEN_3557 = _GEN_1168 ? (_GEN_3526 ? ~_GEN_325 & _GEN_3524 : ~(_GEN_1172 & _GEN_325) & _GEN_3524) : _GEN_3524;
  wire        _GEN_3558 = _GEN_1168 ? (_GEN_3526 ? ~(&lcam_ldq_idx_0) & _GEN_3525 : ~(_GEN_1172 & (&lcam_ldq_idx_0)) & _GEN_3525) : _GEN_3525;
  wire        _GEN_3559 = _GEN_1176 | _GEN_1177;
  wire        _GEN_3560 = _GEN_1174 ? (_GEN_3559 ? (|lcam_ldq_idx_1) & _GEN_3527 : ~(_GEN_1172 & ~(|lcam_ldq_idx_1)) & _GEN_3527) : _GEN_3527;
  wire        _GEN_3561 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_336 & _GEN_3528 : ~(_GEN_1172 & _GEN_336) & _GEN_3528) : _GEN_3528;
  wire        _GEN_3562 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_337 & _GEN_3529 : ~(_GEN_1172 & _GEN_337) & _GEN_3529) : _GEN_3529;
  wire        _GEN_3563 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_338 & _GEN_3530 : ~(_GEN_1172 & _GEN_338) & _GEN_3530) : _GEN_3530;
  wire        _GEN_3564 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_339 & _GEN_3531 : ~(_GEN_1172 & _GEN_339) & _GEN_3531) : _GEN_3531;
  wire        _GEN_3565 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_340 & _GEN_3532 : ~(_GEN_1172 & _GEN_340) & _GEN_3532) : _GEN_3532;
  wire        _GEN_3566 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_341 & _GEN_3533 : ~(_GEN_1172 & _GEN_341) & _GEN_3533) : _GEN_3533;
  wire        _GEN_3567 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_342 & _GEN_3534 : ~(_GEN_1172 & _GEN_342) & _GEN_3534) : _GEN_3534;
  wire        _GEN_3568 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_343 & _GEN_3535 : ~(_GEN_1172 & _GEN_343) & _GEN_3535) : _GEN_3535;
  wire        _GEN_3569 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_344 & _GEN_3536 : ~(_GEN_1172 & _GEN_344) & _GEN_3536) : _GEN_3536;
  wire        _GEN_3570 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_345 & _GEN_3537 : ~(_GEN_1172 & _GEN_345) & _GEN_3537) : _GEN_3537;
  wire        _GEN_3571 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_346 & _GEN_3538 : ~(_GEN_1172 & _GEN_346) & _GEN_3538) : _GEN_3538;
  wire        _GEN_3572 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_347 & _GEN_3539 : ~(_GEN_1172 & _GEN_347) & _GEN_3539) : _GEN_3539;
  wire        _GEN_3573 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_348 & _GEN_3540 : ~(_GEN_1172 & _GEN_348) & _GEN_3540) : _GEN_3540;
  wire        _GEN_3574 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_349 & _GEN_3541 : ~(_GEN_1172 & _GEN_349) & _GEN_3541) : _GEN_3541;
  wire        _GEN_3575 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_350 & _GEN_3542 : ~(_GEN_1172 & _GEN_350) & _GEN_3542) : _GEN_3542;
  wire        _GEN_3576 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_351 & _GEN_3543 : ~(_GEN_1172 & _GEN_351) & _GEN_3543) : _GEN_3543;
  wire        _GEN_3577 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_352 & _GEN_3544 : ~(_GEN_1172 & _GEN_352) & _GEN_3544) : _GEN_3544;
  wire        _GEN_3578 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_353 & _GEN_3545 : ~(_GEN_1172 & _GEN_353) & _GEN_3545) : _GEN_3545;
  wire        _GEN_3579 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_354 & _GEN_3546 : ~(_GEN_1172 & _GEN_354) & _GEN_3546) : _GEN_3546;
  wire        _GEN_3580 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_355 & _GEN_3547 : ~(_GEN_1172 & _GEN_355) & _GEN_3547) : _GEN_3547;
  wire        _GEN_3581 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_356 & _GEN_3548 : ~(_GEN_1172 & _GEN_356) & _GEN_3548) : _GEN_3548;
  wire        _GEN_3582 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_357 & _GEN_3549 : ~(_GEN_1172 & _GEN_357) & _GEN_3549) : _GEN_3549;
  wire        _GEN_3583 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_358 & _GEN_3550 : ~(_GEN_1172 & _GEN_358) & _GEN_3550) : _GEN_3550;
  wire        _GEN_3584 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_359 & _GEN_3551 : ~(_GEN_1172 & _GEN_359) & _GEN_3551) : _GEN_3551;
  wire        _GEN_3585 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_360 & _GEN_3552 : ~(_GEN_1172 & _GEN_360) & _GEN_3552) : _GEN_3552;
  wire        _GEN_3586 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_361 & _GEN_3553 : ~(_GEN_1172 & _GEN_361) & _GEN_3553) : _GEN_3553;
  wire        _GEN_3587 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_362 & _GEN_3554 : ~(_GEN_1172 & _GEN_362) & _GEN_3554) : _GEN_3554;
  wire        _GEN_3588 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_363 & _GEN_3555 : ~(_GEN_1172 & _GEN_363) & _GEN_3555) : _GEN_3555;
  wire        _GEN_3589 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_364 & _GEN_3556 : ~(_GEN_1172 & _GEN_364) & _GEN_3556) : _GEN_3556;
  wire        _GEN_3590 = _GEN_1174 ? (_GEN_3559 ? ~_GEN_365 & _GEN_3557 : ~(_GEN_1172 & _GEN_365) & _GEN_3557) : _GEN_3557;
  wire        _GEN_3591 = _GEN_1174 ? (_GEN_3559 ? ~(&lcam_ldq_idx_1) & _GEN_3558 : ~(_GEN_1172 & (&lcam_ldq_idx_1)) & _GEN_3558) : _GEN_3558;
  wire        _GEN_3592 = _GEN_1181 | _GEN_1182;
  wire        _GEN_3593 = _GEN_1179 ? (_GEN_3592 ? (|lcam_ldq_idx_0) & _GEN_3560 : ~(_GEN_1183 & ~(|lcam_ldq_idx_0)) & _GEN_3560) : _GEN_3560;
  wire        _GEN_3594 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_296 & _GEN_3561 : ~(_GEN_1183 & _GEN_296) & _GEN_3561) : _GEN_3561;
  wire        _GEN_3595 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_297 & _GEN_3562 : ~(_GEN_1183 & _GEN_297) & _GEN_3562) : _GEN_3562;
  wire        _GEN_3596 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_298 & _GEN_3563 : ~(_GEN_1183 & _GEN_298) & _GEN_3563) : _GEN_3563;
  wire        _GEN_3597 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_299 & _GEN_3564 : ~(_GEN_1183 & _GEN_299) & _GEN_3564) : _GEN_3564;
  wire        _GEN_3598 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_300 & _GEN_3565 : ~(_GEN_1183 & _GEN_300) & _GEN_3565) : _GEN_3565;
  wire        _GEN_3599 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_301 & _GEN_3566 : ~(_GEN_1183 & _GEN_301) & _GEN_3566) : _GEN_3566;
  wire        _GEN_3600 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_302 & _GEN_3567 : ~(_GEN_1183 & _GEN_302) & _GEN_3567) : _GEN_3567;
  wire        _GEN_3601 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_303 & _GEN_3568 : ~(_GEN_1183 & _GEN_303) & _GEN_3568) : _GEN_3568;
  wire        _GEN_3602 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_304 & _GEN_3569 : ~(_GEN_1183 & _GEN_304) & _GEN_3569) : _GEN_3569;
  wire        _GEN_3603 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_305 & _GEN_3570 : ~(_GEN_1183 & _GEN_305) & _GEN_3570) : _GEN_3570;
  wire        _GEN_3604 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_306 & _GEN_3571 : ~(_GEN_1183 & _GEN_306) & _GEN_3571) : _GEN_3571;
  wire        _GEN_3605 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_307 & _GEN_3572 : ~(_GEN_1183 & _GEN_307) & _GEN_3572) : _GEN_3572;
  wire        _GEN_3606 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_308 & _GEN_3573 : ~(_GEN_1183 & _GEN_308) & _GEN_3573) : _GEN_3573;
  wire        _GEN_3607 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_309 & _GEN_3574 : ~(_GEN_1183 & _GEN_309) & _GEN_3574) : _GEN_3574;
  wire        _GEN_3608 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_310 & _GEN_3575 : ~(_GEN_1183 & _GEN_310) & _GEN_3575) : _GEN_3575;
  wire        _GEN_3609 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_311 & _GEN_3576 : ~(_GEN_1183 & _GEN_311) & _GEN_3576) : _GEN_3576;
  wire        _GEN_3610 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_312 & _GEN_3577 : ~(_GEN_1183 & _GEN_312) & _GEN_3577) : _GEN_3577;
  wire        _GEN_3611 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_313 & _GEN_3578 : ~(_GEN_1183 & _GEN_313) & _GEN_3578) : _GEN_3578;
  wire        _GEN_3612 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_314 & _GEN_3579 : ~(_GEN_1183 & _GEN_314) & _GEN_3579) : _GEN_3579;
  wire        _GEN_3613 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_315 & _GEN_3580 : ~(_GEN_1183 & _GEN_315) & _GEN_3580) : _GEN_3580;
  wire        _GEN_3614 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_316 & _GEN_3581 : ~(_GEN_1183 & _GEN_316) & _GEN_3581) : _GEN_3581;
  wire        _GEN_3615 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_317 & _GEN_3582 : ~(_GEN_1183 & _GEN_317) & _GEN_3582) : _GEN_3582;
  wire        _GEN_3616 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_318 & _GEN_3583 : ~(_GEN_1183 & _GEN_318) & _GEN_3583) : _GEN_3583;
  wire        _GEN_3617 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_319 & _GEN_3584 : ~(_GEN_1183 & _GEN_319) & _GEN_3584) : _GEN_3584;
  wire        _GEN_3618 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_320 & _GEN_3585 : ~(_GEN_1183 & _GEN_320) & _GEN_3585) : _GEN_3585;
  wire        _GEN_3619 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_321 & _GEN_3586 : ~(_GEN_1183 & _GEN_321) & _GEN_3586) : _GEN_3586;
  wire        _GEN_3620 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_322 & _GEN_3587 : ~(_GEN_1183 & _GEN_322) & _GEN_3587) : _GEN_3587;
  wire        _GEN_3621 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_323 & _GEN_3588 : ~(_GEN_1183 & _GEN_323) & _GEN_3588) : _GEN_3588;
  wire        _GEN_3622 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_324 & _GEN_3589 : ~(_GEN_1183 & _GEN_324) & _GEN_3589) : _GEN_3589;
  wire        _GEN_3623 = _GEN_1179 ? (_GEN_3592 ? ~_GEN_325 & _GEN_3590 : ~(_GEN_1183 & _GEN_325) & _GEN_3590) : _GEN_3590;
  wire        _GEN_3624 = _GEN_1179 ? (_GEN_3592 ? ~(&lcam_ldq_idx_0) & _GEN_3591 : ~(_GEN_1183 & (&lcam_ldq_idx_0)) & _GEN_3591) : _GEN_3591;
  wire        _GEN_3625 = _GEN_1187 | _GEN_1188;
  wire        _GEN_3626 = _GEN_1185 ? (_GEN_3625 ? (|lcam_ldq_idx_1) & _GEN_3593 : ~(_GEN_1183 & ~(|lcam_ldq_idx_1)) & _GEN_3593) : _GEN_3593;
  wire        _GEN_3627 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_336 & _GEN_3594 : ~(_GEN_1183 & _GEN_336) & _GEN_3594) : _GEN_3594;
  wire        _GEN_3628 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_337 & _GEN_3595 : ~(_GEN_1183 & _GEN_337) & _GEN_3595) : _GEN_3595;
  wire        _GEN_3629 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_338 & _GEN_3596 : ~(_GEN_1183 & _GEN_338) & _GEN_3596) : _GEN_3596;
  wire        _GEN_3630 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_339 & _GEN_3597 : ~(_GEN_1183 & _GEN_339) & _GEN_3597) : _GEN_3597;
  wire        _GEN_3631 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_340 & _GEN_3598 : ~(_GEN_1183 & _GEN_340) & _GEN_3598) : _GEN_3598;
  wire        _GEN_3632 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_341 & _GEN_3599 : ~(_GEN_1183 & _GEN_341) & _GEN_3599) : _GEN_3599;
  wire        _GEN_3633 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_342 & _GEN_3600 : ~(_GEN_1183 & _GEN_342) & _GEN_3600) : _GEN_3600;
  wire        _GEN_3634 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_343 & _GEN_3601 : ~(_GEN_1183 & _GEN_343) & _GEN_3601) : _GEN_3601;
  wire        _GEN_3635 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_344 & _GEN_3602 : ~(_GEN_1183 & _GEN_344) & _GEN_3602) : _GEN_3602;
  wire        _GEN_3636 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_345 & _GEN_3603 : ~(_GEN_1183 & _GEN_345) & _GEN_3603) : _GEN_3603;
  wire        _GEN_3637 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_346 & _GEN_3604 : ~(_GEN_1183 & _GEN_346) & _GEN_3604) : _GEN_3604;
  wire        _GEN_3638 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_347 & _GEN_3605 : ~(_GEN_1183 & _GEN_347) & _GEN_3605) : _GEN_3605;
  wire        _GEN_3639 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_348 & _GEN_3606 : ~(_GEN_1183 & _GEN_348) & _GEN_3606) : _GEN_3606;
  wire        _GEN_3640 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_349 & _GEN_3607 : ~(_GEN_1183 & _GEN_349) & _GEN_3607) : _GEN_3607;
  wire        _GEN_3641 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_350 & _GEN_3608 : ~(_GEN_1183 & _GEN_350) & _GEN_3608) : _GEN_3608;
  wire        _GEN_3642 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_351 & _GEN_3609 : ~(_GEN_1183 & _GEN_351) & _GEN_3609) : _GEN_3609;
  wire        _GEN_3643 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_352 & _GEN_3610 : ~(_GEN_1183 & _GEN_352) & _GEN_3610) : _GEN_3610;
  wire        _GEN_3644 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_353 & _GEN_3611 : ~(_GEN_1183 & _GEN_353) & _GEN_3611) : _GEN_3611;
  wire        _GEN_3645 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_354 & _GEN_3612 : ~(_GEN_1183 & _GEN_354) & _GEN_3612) : _GEN_3612;
  wire        _GEN_3646 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_355 & _GEN_3613 : ~(_GEN_1183 & _GEN_355) & _GEN_3613) : _GEN_3613;
  wire        _GEN_3647 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_356 & _GEN_3614 : ~(_GEN_1183 & _GEN_356) & _GEN_3614) : _GEN_3614;
  wire        _GEN_3648 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_357 & _GEN_3615 : ~(_GEN_1183 & _GEN_357) & _GEN_3615) : _GEN_3615;
  wire        _GEN_3649 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_358 & _GEN_3616 : ~(_GEN_1183 & _GEN_358) & _GEN_3616) : _GEN_3616;
  wire        _GEN_3650 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_359 & _GEN_3617 : ~(_GEN_1183 & _GEN_359) & _GEN_3617) : _GEN_3617;
  wire        _GEN_3651 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_360 & _GEN_3618 : ~(_GEN_1183 & _GEN_360) & _GEN_3618) : _GEN_3618;
  wire        _GEN_3652 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_361 & _GEN_3619 : ~(_GEN_1183 & _GEN_361) & _GEN_3619) : _GEN_3619;
  wire        _GEN_3653 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_362 & _GEN_3620 : ~(_GEN_1183 & _GEN_362) & _GEN_3620) : _GEN_3620;
  wire        _GEN_3654 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_363 & _GEN_3621 : ~(_GEN_1183 & _GEN_363) & _GEN_3621) : _GEN_3621;
  wire        _GEN_3655 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_364 & _GEN_3622 : ~(_GEN_1183 & _GEN_364) & _GEN_3622) : _GEN_3622;
  wire        _GEN_3656 = _GEN_1185 ? (_GEN_3625 ? ~_GEN_365 & _GEN_3623 : ~(_GEN_1183 & _GEN_365) & _GEN_3623) : _GEN_3623;
  wire        _GEN_3657 = _GEN_1185 ? (_GEN_3625 ? ~(&lcam_ldq_idx_1) & _GEN_3624 : ~(_GEN_1183 & (&lcam_ldq_idx_1)) & _GEN_3624) : _GEN_3624;
  wire        _GEN_3658 = _GEN_1192 | _GEN_1193;
  wire        _GEN_3659 = _GEN_1190 ? (_GEN_3658 ? (|lcam_ldq_idx_0) & _GEN_3626 : ~(_GEN_1194 & ~(|lcam_ldq_idx_0)) & _GEN_3626) : _GEN_3626;
  wire        _GEN_3660 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_296 & _GEN_3627 : ~(_GEN_1194 & _GEN_296) & _GEN_3627) : _GEN_3627;
  wire        _GEN_3661 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_297 & _GEN_3628 : ~(_GEN_1194 & _GEN_297) & _GEN_3628) : _GEN_3628;
  wire        _GEN_3662 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_298 & _GEN_3629 : ~(_GEN_1194 & _GEN_298) & _GEN_3629) : _GEN_3629;
  wire        _GEN_3663 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_299 & _GEN_3630 : ~(_GEN_1194 & _GEN_299) & _GEN_3630) : _GEN_3630;
  wire        _GEN_3664 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_300 & _GEN_3631 : ~(_GEN_1194 & _GEN_300) & _GEN_3631) : _GEN_3631;
  wire        _GEN_3665 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_301 & _GEN_3632 : ~(_GEN_1194 & _GEN_301) & _GEN_3632) : _GEN_3632;
  wire        _GEN_3666 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_302 & _GEN_3633 : ~(_GEN_1194 & _GEN_302) & _GEN_3633) : _GEN_3633;
  wire        _GEN_3667 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_303 & _GEN_3634 : ~(_GEN_1194 & _GEN_303) & _GEN_3634) : _GEN_3634;
  wire        _GEN_3668 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_304 & _GEN_3635 : ~(_GEN_1194 & _GEN_304) & _GEN_3635) : _GEN_3635;
  wire        _GEN_3669 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_305 & _GEN_3636 : ~(_GEN_1194 & _GEN_305) & _GEN_3636) : _GEN_3636;
  wire        _GEN_3670 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_306 & _GEN_3637 : ~(_GEN_1194 & _GEN_306) & _GEN_3637) : _GEN_3637;
  wire        _GEN_3671 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_307 & _GEN_3638 : ~(_GEN_1194 & _GEN_307) & _GEN_3638) : _GEN_3638;
  wire        _GEN_3672 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_308 & _GEN_3639 : ~(_GEN_1194 & _GEN_308) & _GEN_3639) : _GEN_3639;
  wire        _GEN_3673 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_309 & _GEN_3640 : ~(_GEN_1194 & _GEN_309) & _GEN_3640) : _GEN_3640;
  wire        _GEN_3674 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_310 & _GEN_3641 : ~(_GEN_1194 & _GEN_310) & _GEN_3641) : _GEN_3641;
  wire        _GEN_3675 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_311 & _GEN_3642 : ~(_GEN_1194 & _GEN_311) & _GEN_3642) : _GEN_3642;
  wire        _GEN_3676 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_312 & _GEN_3643 : ~(_GEN_1194 & _GEN_312) & _GEN_3643) : _GEN_3643;
  wire        _GEN_3677 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_313 & _GEN_3644 : ~(_GEN_1194 & _GEN_313) & _GEN_3644) : _GEN_3644;
  wire        _GEN_3678 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_314 & _GEN_3645 : ~(_GEN_1194 & _GEN_314) & _GEN_3645) : _GEN_3645;
  wire        _GEN_3679 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_315 & _GEN_3646 : ~(_GEN_1194 & _GEN_315) & _GEN_3646) : _GEN_3646;
  wire        _GEN_3680 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_316 & _GEN_3647 : ~(_GEN_1194 & _GEN_316) & _GEN_3647) : _GEN_3647;
  wire        _GEN_3681 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_317 & _GEN_3648 : ~(_GEN_1194 & _GEN_317) & _GEN_3648) : _GEN_3648;
  wire        _GEN_3682 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_318 & _GEN_3649 : ~(_GEN_1194 & _GEN_318) & _GEN_3649) : _GEN_3649;
  wire        _GEN_3683 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_319 & _GEN_3650 : ~(_GEN_1194 & _GEN_319) & _GEN_3650) : _GEN_3650;
  wire        _GEN_3684 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_320 & _GEN_3651 : ~(_GEN_1194 & _GEN_320) & _GEN_3651) : _GEN_3651;
  wire        _GEN_3685 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_321 & _GEN_3652 : ~(_GEN_1194 & _GEN_321) & _GEN_3652) : _GEN_3652;
  wire        _GEN_3686 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_322 & _GEN_3653 : ~(_GEN_1194 & _GEN_322) & _GEN_3653) : _GEN_3653;
  wire        _GEN_3687 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_323 & _GEN_3654 : ~(_GEN_1194 & _GEN_323) & _GEN_3654) : _GEN_3654;
  wire        _GEN_3688 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_324 & _GEN_3655 : ~(_GEN_1194 & _GEN_324) & _GEN_3655) : _GEN_3655;
  wire        _GEN_3689 = _GEN_1190 ? (_GEN_3658 ? ~_GEN_325 & _GEN_3656 : ~(_GEN_1194 & _GEN_325) & _GEN_3656) : _GEN_3656;
  wire        _GEN_3690 = _GEN_1190 ? (_GEN_3658 ? ~(&lcam_ldq_idx_0) & _GEN_3657 : ~(_GEN_1194 & (&lcam_ldq_idx_0)) & _GEN_3657) : _GEN_3657;
  wire        _GEN_3691 = _GEN_1198 | _GEN_1199;
  wire        _GEN_3692 = _GEN_1196 ? (_GEN_3691 ? (|lcam_ldq_idx_1) & _GEN_3659 : ~(_GEN_1194 & ~(|lcam_ldq_idx_1)) & _GEN_3659) : _GEN_3659;
  wire        _GEN_3693 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_336 & _GEN_3660 : ~(_GEN_1194 & _GEN_336) & _GEN_3660) : _GEN_3660;
  wire        _GEN_3694 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_337 & _GEN_3661 : ~(_GEN_1194 & _GEN_337) & _GEN_3661) : _GEN_3661;
  wire        _GEN_3695 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_338 & _GEN_3662 : ~(_GEN_1194 & _GEN_338) & _GEN_3662) : _GEN_3662;
  wire        _GEN_3696 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_339 & _GEN_3663 : ~(_GEN_1194 & _GEN_339) & _GEN_3663) : _GEN_3663;
  wire        _GEN_3697 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_340 & _GEN_3664 : ~(_GEN_1194 & _GEN_340) & _GEN_3664) : _GEN_3664;
  wire        _GEN_3698 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_341 & _GEN_3665 : ~(_GEN_1194 & _GEN_341) & _GEN_3665) : _GEN_3665;
  wire        _GEN_3699 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_342 & _GEN_3666 : ~(_GEN_1194 & _GEN_342) & _GEN_3666) : _GEN_3666;
  wire        _GEN_3700 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_343 & _GEN_3667 : ~(_GEN_1194 & _GEN_343) & _GEN_3667) : _GEN_3667;
  wire        _GEN_3701 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_344 & _GEN_3668 : ~(_GEN_1194 & _GEN_344) & _GEN_3668) : _GEN_3668;
  wire        _GEN_3702 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_345 & _GEN_3669 : ~(_GEN_1194 & _GEN_345) & _GEN_3669) : _GEN_3669;
  wire        _GEN_3703 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_346 & _GEN_3670 : ~(_GEN_1194 & _GEN_346) & _GEN_3670) : _GEN_3670;
  wire        _GEN_3704 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_347 & _GEN_3671 : ~(_GEN_1194 & _GEN_347) & _GEN_3671) : _GEN_3671;
  wire        _GEN_3705 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_348 & _GEN_3672 : ~(_GEN_1194 & _GEN_348) & _GEN_3672) : _GEN_3672;
  wire        _GEN_3706 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_349 & _GEN_3673 : ~(_GEN_1194 & _GEN_349) & _GEN_3673) : _GEN_3673;
  wire        _GEN_3707 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_350 & _GEN_3674 : ~(_GEN_1194 & _GEN_350) & _GEN_3674) : _GEN_3674;
  wire        _GEN_3708 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_351 & _GEN_3675 : ~(_GEN_1194 & _GEN_351) & _GEN_3675) : _GEN_3675;
  wire        _GEN_3709 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_352 & _GEN_3676 : ~(_GEN_1194 & _GEN_352) & _GEN_3676) : _GEN_3676;
  wire        _GEN_3710 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_353 & _GEN_3677 : ~(_GEN_1194 & _GEN_353) & _GEN_3677) : _GEN_3677;
  wire        _GEN_3711 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_354 & _GEN_3678 : ~(_GEN_1194 & _GEN_354) & _GEN_3678) : _GEN_3678;
  wire        _GEN_3712 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_355 & _GEN_3679 : ~(_GEN_1194 & _GEN_355) & _GEN_3679) : _GEN_3679;
  wire        _GEN_3713 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_356 & _GEN_3680 : ~(_GEN_1194 & _GEN_356) & _GEN_3680) : _GEN_3680;
  wire        _GEN_3714 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_357 & _GEN_3681 : ~(_GEN_1194 & _GEN_357) & _GEN_3681) : _GEN_3681;
  wire        _GEN_3715 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_358 & _GEN_3682 : ~(_GEN_1194 & _GEN_358) & _GEN_3682) : _GEN_3682;
  wire        _GEN_3716 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_359 & _GEN_3683 : ~(_GEN_1194 & _GEN_359) & _GEN_3683) : _GEN_3683;
  wire        _GEN_3717 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_360 & _GEN_3684 : ~(_GEN_1194 & _GEN_360) & _GEN_3684) : _GEN_3684;
  wire        _GEN_3718 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_361 & _GEN_3685 : ~(_GEN_1194 & _GEN_361) & _GEN_3685) : _GEN_3685;
  wire        _GEN_3719 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_362 & _GEN_3686 : ~(_GEN_1194 & _GEN_362) & _GEN_3686) : _GEN_3686;
  wire        _GEN_3720 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_363 & _GEN_3687 : ~(_GEN_1194 & _GEN_363) & _GEN_3687) : _GEN_3687;
  wire        _GEN_3721 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_364 & _GEN_3688 : ~(_GEN_1194 & _GEN_364) & _GEN_3688) : _GEN_3688;
  wire        _GEN_3722 = _GEN_1196 ? (_GEN_3691 ? ~_GEN_365 & _GEN_3689 : ~(_GEN_1194 & _GEN_365) & _GEN_3689) : _GEN_3689;
  wire        _GEN_3723 = _GEN_1196 ? (_GEN_3691 ? ~(&lcam_ldq_idx_1) & _GEN_3690 : ~(_GEN_1194 & (&lcam_ldq_idx_1)) & _GEN_3690) : _GEN_3690;
  wire        _GEN_3724 = _GEN_1203 | _GEN_1204;
  wire        _GEN_3725 = _GEN_1201 ? (_GEN_3724 ? (|lcam_ldq_idx_0) & _GEN_3692 : ~(_GEN_1205 & ~(|lcam_ldq_idx_0)) & _GEN_3692) : _GEN_3692;
  wire        _GEN_3726 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_296 & _GEN_3693 : ~(_GEN_1205 & _GEN_296) & _GEN_3693) : _GEN_3693;
  wire        _GEN_3727 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_297 & _GEN_3694 : ~(_GEN_1205 & _GEN_297) & _GEN_3694) : _GEN_3694;
  wire        _GEN_3728 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_298 & _GEN_3695 : ~(_GEN_1205 & _GEN_298) & _GEN_3695) : _GEN_3695;
  wire        _GEN_3729 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_299 & _GEN_3696 : ~(_GEN_1205 & _GEN_299) & _GEN_3696) : _GEN_3696;
  wire        _GEN_3730 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_300 & _GEN_3697 : ~(_GEN_1205 & _GEN_300) & _GEN_3697) : _GEN_3697;
  wire        _GEN_3731 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_301 & _GEN_3698 : ~(_GEN_1205 & _GEN_301) & _GEN_3698) : _GEN_3698;
  wire        _GEN_3732 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_302 & _GEN_3699 : ~(_GEN_1205 & _GEN_302) & _GEN_3699) : _GEN_3699;
  wire        _GEN_3733 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_303 & _GEN_3700 : ~(_GEN_1205 & _GEN_303) & _GEN_3700) : _GEN_3700;
  wire        _GEN_3734 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_304 & _GEN_3701 : ~(_GEN_1205 & _GEN_304) & _GEN_3701) : _GEN_3701;
  wire        _GEN_3735 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_305 & _GEN_3702 : ~(_GEN_1205 & _GEN_305) & _GEN_3702) : _GEN_3702;
  wire        _GEN_3736 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_306 & _GEN_3703 : ~(_GEN_1205 & _GEN_306) & _GEN_3703) : _GEN_3703;
  wire        _GEN_3737 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_307 & _GEN_3704 : ~(_GEN_1205 & _GEN_307) & _GEN_3704) : _GEN_3704;
  wire        _GEN_3738 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_308 & _GEN_3705 : ~(_GEN_1205 & _GEN_308) & _GEN_3705) : _GEN_3705;
  wire        _GEN_3739 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_309 & _GEN_3706 : ~(_GEN_1205 & _GEN_309) & _GEN_3706) : _GEN_3706;
  wire        _GEN_3740 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_310 & _GEN_3707 : ~(_GEN_1205 & _GEN_310) & _GEN_3707) : _GEN_3707;
  wire        _GEN_3741 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_311 & _GEN_3708 : ~(_GEN_1205 & _GEN_311) & _GEN_3708) : _GEN_3708;
  wire        _GEN_3742 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_312 & _GEN_3709 : ~(_GEN_1205 & _GEN_312) & _GEN_3709) : _GEN_3709;
  wire        _GEN_3743 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_313 & _GEN_3710 : ~(_GEN_1205 & _GEN_313) & _GEN_3710) : _GEN_3710;
  wire        _GEN_3744 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_314 & _GEN_3711 : ~(_GEN_1205 & _GEN_314) & _GEN_3711) : _GEN_3711;
  wire        _GEN_3745 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_315 & _GEN_3712 : ~(_GEN_1205 & _GEN_315) & _GEN_3712) : _GEN_3712;
  wire        _GEN_3746 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_316 & _GEN_3713 : ~(_GEN_1205 & _GEN_316) & _GEN_3713) : _GEN_3713;
  wire        _GEN_3747 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_317 & _GEN_3714 : ~(_GEN_1205 & _GEN_317) & _GEN_3714) : _GEN_3714;
  wire        _GEN_3748 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_318 & _GEN_3715 : ~(_GEN_1205 & _GEN_318) & _GEN_3715) : _GEN_3715;
  wire        _GEN_3749 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_319 & _GEN_3716 : ~(_GEN_1205 & _GEN_319) & _GEN_3716) : _GEN_3716;
  wire        _GEN_3750 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_320 & _GEN_3717 : ~(_GEN_1205 & _GEN_320) & _GEN_3717) : _GEN_3717;
  wire        _GEN_3751 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_321 & _GEN_3718 : ~(_GEN_1205 & _GEN_321) & _GEN_3718) : _GEN_3718;
  wire        _GEN_3752 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_322 & _GEN_3719 : ~(_GEN_1205 & _GEN_322) & _GEN_3719) : _GEN_3719;
  wire        _GEN_3753 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_323 & _GEN_3720 : ~(_GEN_1205 & _GEN_323) & _GEN_3720) : _GEN_3720;
  wire        _GEN_3754 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_324 & _GEN_3721 : ~(_GEN_1205 & _GEN_324) & _GEN_3721) : _GEN_3721;
  wire        _GEN_3755 = _GEN_1201 ? (_GEN_3724 ? ~_GEN_325 & _GEN_3722 : ~(_GEN_1205 & _GEN_325) & _GEN_3722) : _GEN_3722;
  wire        _GEN_3756 = _GEN_1201 ? (_GEN_3724 ? ~(&lcam_ldq_idx_0) & _GEN_3723 : ~(_GEN_1205 & (&lcam_ldq_idx_0)) & _GEN_3723) : _GEN_3723;
  wire        _GEN_3757 = _GEN_1209 | _GEN_1210;
  wire        _GEN_3758 = _GEN_1207 ? (_GEN_3757 ? (|lcam_ldq_idx_1) & _GEN_3725 : ~(_GEN_1205 & ~(|lcam_ldq_idx_1)) & _GEN_3725) : _GEN_3725;
  wire        _GEN_3759 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_336 & _GEN_3726 : ~(_GEN_1205 & _GEN_336) & _GEN_3726) : _GEN_3726;
  wire        _GEN_3760 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_337 & _GEN_3727 : ~(_GEN_1205 & _GEN_337) & _GEN_3727) : _GEN_3727;
  wire        _GEN_3761 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_338 & _GEN_3728 : ~(_GEN_1205 & _GEN_338) & _GEN_3728) : _GEN_3728;
  wire        _GEN_3762 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_339 & _GEN_3729 : ~(_GEN_1205 & _GEN_339) & _GEN_3729) : _GEN_3729;
  wire        _GEN_3763 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_340 & _GEN_3730 : ~(_GEN_1205 & _GEN_340) & _GEN_3730) : _GEN_3730;
  wire        _GEN_3764 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_341 & _GEN_3731 : ~(_GEN_1205 & _GEN_341) & _GEN_3731) : _GEN_3731;
  wire        _GEN_3765 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_342 & _GEN_3732 : ~(_GEN_1205 & _GEN_342) & _GEN_3732) : _GEN_3732;
  wire        _GEN_3766 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_343 & _GEN_3733 : ~(_GEN_1205 & _GEN_343) & _GEN_3733) : _GEN_3733;
  wire        _GEN_3767 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_344 & _GEN_3734 : ~(_GEN_1205 & _GEN_344) & _GEN_3734) : _GEN_3734;
  wire        _GEN_3768 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_345 & _GEN_3735 : ~(_GEN_1205 & _GEN_345) & _GEN_3735) : _GEN_3735;
  wire        _GEN_3769 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_346 & _GEN_3736 : ~(_GEN_1205 & _GEN_346) & _GEN_3736) : _GEN_3736;
  wire        _GEN_3770 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_347 & _GEN_3737 : ~(_GEN_1205 & _GEN_347) & _GEN_3737) : _GEN_3737;
  wire        _GEN_3771 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_348 & _GEN_3738 : ~(_GEN_1205 & _GEN_348) & _GEN_3738) : _GEN_3738;
  wire        _GEN_3772 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_349 & _GEN_3739 : ~(_GEN_1205 & _GEN_349) & _GEN_3739) : _GEN_3739;
  wire        _GEN_3773 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_350 & _GEN_3740 : ~(_GEN_1205 & _GEN_350) & _GEN_3740) : _GEN_3740;
  wire        _GEN_3774 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_351 & _GEN_3741 : ~(_GEN_1205 & _GEN_351) & _GEN_3741) : _GEN_3741;
  wire        _GEN_3775 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_352 & _GEN_3742 : ~(_GEN_1205 & _GEN_352) & _GEN_3742) : _GEN_3742;
  wire        _GEN_3776 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_353 & _GEN_3743 : ~(_GEN_1205 & _GEN_353) & _GEN_3743) : _GEN_3743;
  wire        _GEN_3777 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_354 & _GEN_3744 : ~(_GEN_1205 & _GEN_354) & _GEN_3744) : _GEN_3744;
  wire        _GEN_3778 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_355 & _GEN_3745 : ~(_GEN_1205 & _GEN_355) & _GEN_3745) : _GEN_3745;
  wire        _GEN_3779 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_356 & _GEN_3746 : ~(_GEN_1205 & _GEN_356) & _GEN_3746) : _GEN_3746;
  wire        _GEN_3780 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_357 & _GEN_3747 : ~(_GEN_1205 & _GEN_357) & _GEN_3747) : _GEN_3747;
  wire        _GEN_3781 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_358 & _GEN_3748 : ~(_GEN_1205 & _GEN_358) & _GEN_3748) : _GEN_3748;
  wire        _GEN_3782 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_359 & _GEN_3749 : ~(_GEN_1205 & _GEN_359) & _GEN_3749) : _GEN_3749;
  wire        _GEN_3783 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_360 & _GEN_3750 : ~(_GEN_1205 & _GEN_360) & _GEN_3750) : _GEN_3750;
  wire        _GEN_3784 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_361 & _GEN_3751 : ~(_GEN_1205 & _GEN_361) & _GEN_3751) : _GEN_3751;
  wire        _GEN_3785 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_362 & _GEN_3752 : ~(_GEN_1205 & _GEN_362) & _GEN_3752) : _GEN_3752;
  wire        _GEN_3786 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_363 & _GEN_3753 : ~(_GEN_1205 & _GEN_363) & _GEN_3753) : _GEN_3753;
  wire        _GEN_3787 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_364 & _GEN_3754 : ~(_GEN_1205 & _GEN_364) & _GEN_3754) : _GEN_3754;
  wire        _GEN_3788 = _GEN_1207 ? (_GEN_3757 ? ~_GEN_365 & _GEN_3755 : ~(_GEN_1205 & _GEN_365) & _GEN_3755) : _GEN_3755;
  wire        _GEN_3789 = _GEN_1207 ? (_GEN_3757 ? ~(&lcam_ldq_idx_1) & _GEN_3756 : ~(_GEN_1205 & (&lcam_ldq_idx_1)) & _GEN_3756) : _GEN_3756;
  wire        _GEN_3790 = _GEN_1214 | _GEN_1215;
  wire        _GEN_3791 = _GEN_1212 ? (_GEN_3790 ? (|lcam_ldq_idx_0) & _GEN_3758 : ~(_GEN_1216 & ~(|lcam_ldq_idx_0)) & _GEN_3758) : _GEN_3758;
  wire        _GEN_3792 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_296 & _GEN_3759 : ~(_GEN_1216 & _GEN_296) & _GEN_3759) : _GEN_3759;
  wire        _GEN_3793 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_297 & _GEN_3760 : ~(_GEN_1216 & _GEN_297) & _GEN_3760) : _GEN_3760;
  wire        _GEN_3794 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_298 & _GEN_3761 : ~(_GEN_1216 & _GEN_298) & _GEN_3761) : _GEN_3761;
  wire        _GEN_3795 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_299 & _GEN_3762 : ~(_GEN_1216 & _GEN_299) & _GEN_3762) : _GEN_3762;
  wire        _GEN_3796 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_300 & _GEN_3763 : ~(_GEN_1216 & _GEN_300) & _GEN_3763) : _GEN_3763;
  wire        _GEN_3797 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_301 & _GEN_3764 : ~(_GEN_1216 & _GEN_301) & _GEN_3764) : _GEN_3764;
  wire        _GEN_3798 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_302 & _GEN_3765 : ~(_GEN_1216 & _GEN_302) & _GEN_3765) : _GEN_3765;
  wire        _GEN_3799 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_303 & _GEN_3766 : ~(_GEN_1216 & _GEN_303) & _GEN_3766) : _GEN_3766;
  wire        _GEN_3800 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_304 & _GEN_3767 : ~(_GEN_1216 & _GEN_304) & _GEN_3767) : _GEN_3767;
  wire        _GEN_3801 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_305 & _GEN_3768 : ~(_GEN_1216 & _GEN_305) & _GEN_3768) : _GEN_3768;
  wire        _GEN_3802 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_306 & _GEN_3769 : ~(_GEN_1216 & _GEN_306) & _GEN_3769) : _GEN_3769;
  wire        _GEN_3803 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_307 & _GEN_3770 : ~(_GEN_1216 & _GEN_307) & _GEN_3770) : _GEN_3770;
  wire        _GEN_3804 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_308 & _GEN_3771 : ~(_GEN_1216 & _GEN_308) & _GEN_3771) : _GEN_3771;
  wire        _GEN_3805 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_309 & _GEN_3772 : ~(_GEN_1216 & _GEN_309) & _GEN_3772) : _GEN_3772;
  wire        _GEN_3806 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_310 & _GEN_3773 : ~(_GEN_1216 & _GEN_310) & _GEN_3773) : _GEN_3773;
  wire        _GEN_3807 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_311 & _GEN_3774 : ~(_GEN_1216 & _GEN_311) & _GEN_3774) : _GEN_3774;
  wire        _GEN_3808 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_312 & _GEN_3775 : ~(_GEN_1216 & _GEN_312) & _GEN_3775) : _GEN_3775;
  wire        _GEN_3809 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_313 & _GEN_3776 : ~(_GEN_1216 & _GEN_313) & _GEN_3776) : _GEN_3776;
  wire        _GEN_3810 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_314 & _GEN_3777 : ~(_GEN_1216 & _GEN_314) & _GEN_3777) : _GEN_3777;
  wire        _GEN_3811 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_315 & _GEN_3778 : ~(_GEN_1216 & _GEN_315) & _GEN_3778) : _GEN_3778;
  wire        _GEN_3812 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_316 & _GEN_3779 : ~(_GEN_1216 & _GEN_316) & _GEN_3779) : _GEN_3779;
  wire        _GEN_3813 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_317 & _GEN_3780 : ~(_GEN_1216 & _GEN_317) & _GEN_3780) : _GEN_3780;
  wire        _GEN_3814 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_318 & _GEN_3781 : ~(_GEN_1216 & _GEN_318) & _GEN_3781) : _GEN_3781;
  wire        _GEN_3815 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_319 & _GEN_3782 : ~(_GEN_1216 & _GEN_319) & _GEN_3782) : _GEN_3782;
  wire        _GEN_3816 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_320 & _GEN_3783 : ~(_GEN_1216 & _GEN_320) & _GEN_3783) : _GEN_3783;
  wire        _GEN_3817 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_321 & _GEN_3784 : ~(_GEN_1216 & _GEN_321) & _GEN_3784) : _GEN_3784;
  wire        _GEN_3818 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_322 & _GEN_3785 : ~(_GEN_1216 & _GEN_322) & _GEN_3785) : _GEN_3785;
  wire        _GEN_3819 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_323 & _GEN_3786 : ~(_GEN_1216 & _GEN_323) & _GEN_3786) : _GEN_3786;
  wire        _GEN_3820 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_324 & _GEN_3787 : ~(_GEN_1216 & _GEN_324) & _GEN_3787) : _GEN_3787;
  wire        _GEN_3821 = _GEN_1212 ? (_GEN_3790 ? ~_GEN_325 & _GEN_3788 : ~(_GEN_1216 & _GEN_325) & _GEN_3788) : _GEN_3788;
  wire        _GEN_3822 = _GEN_1212 ? (_GEN_3790 ? ~(&lcam_ldq_idx_0) & _GEN_3789 : ~(_GEN_1216 & (&lcam_ldq_idx_0)) & _GEN_3789) : _GEN_3789;
  wire        _GEN_3823 = _GEN_1220 | _GEN_1221;
  wire        _GEN_3824 = _GEN_1218 ? (_GEN_3823 ? (|lcam_ldq_idx_1) & _GEN_3791 : ~(_GEN_1216 & ~(|lcam_ldq_idx_1)) & _GEN_3791) : _GEN_3791;
  wire        _GEN_3825 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_336 & _GEN_3792 : ~(_GEN_1216 & _GEN_336) & _GEN_3792) : _GEN_3792;
  wire        _GEN_3826 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_337 & _GEN_3793 : ~(_GEN_1216 & _GEN_337) & _GEN_3793) : _GEN_3793;
  wire        _GEN_3827 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_338 & _GEN_3794 : ~(_GEN_1216 & _GEN_338) & _GEN_3794) : _GEN_3794;
  wire        _GEN_3828 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_339 & _GEN_3795 : ~(_GEN_1216 & _GEN_339) & _GEN_3795) : _GEN_3795;
  wire        _GEN_3829 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_340 & _GEN_3796 : ~(_GEN_1216 & _GEN_340) & _GEN_3796) : _GEN_3796;
  wire        _GEN_3830 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_341 & _GEN_3797 : ~(_GEN_1216 & _GEN_341) & _GEN_3797) : _GEN_3797;
  wire        _GEN_3831 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_342 & _GEN_3798 : ~(_GEN_1216 & _GEN_342) & _GEN_3798) : _GEN_3798;
  wire        _GEN_3832 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_343 & _GEN_3799 : ~(_GEN_1216 & _GEN_343) & _GEN_3799) : _GEN_3799;
  wire        _GEN_3833 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_344 & _GEN_3800 : ~(_GEN_1216 & _GEN_344) & _GEN_3800) : _GEN_3800;
  wire        _GEN_3834 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_345 & _GEN_3801 : ~(_GEN_1216 & _GEN_345) & _GEN_3801) : _GEN_3801;
  wire        _GEN_3835 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_346 & _GEN_3802 : ~(_GEN_1216 & _GEN_346) & _GEN_3802) : _GEN_3802;
  wire        _GEN_3836 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_347 & _GEN_3803 : ~(_GEN_1216 & _GEN_347) & _GEN_3803) : _GEN_3803;
  wire        _GEN_3837 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_348 & _GEN_3804 : ~(_GEN_1216 & _GEN_348) & _GEN_3804) : _GEN_3804;
  wire        _GEN_3838 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_349 & _GEN_3805 : ~(_GEN_1216 & _GEN_349) & _GEN_3805) : _GEN_3805;
  wire        _GEN_3839 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_350 & _GEN_3806 : ~(_GEN_1216 & _GEN_350) & _GEN_3806) : _GEN_3806;
  wire        _GEN_3840 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_351 & _GEN_3807 : ~(_GEN_1216 & _GEN_351) & _GEN_3807) : _GEN_3807;
  wire        _GEN_3841 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_352 & _GEN_3808 : ~(_GEN_1216 & _GEN_352) & _GEN_3808) : _GEN_3808;
  wire        _GEN_3842 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_353 & _GEN_3809 : ~(_GEN_1216 & _GEN_353) & _GEN_3809) : _GEN_3809;
  wire        _GEN_3843 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_354 & _GEN_3810 : ~(_GEN_1216 & _GEN_354) & _GEN_3810) : _GEN_3810;
  wire        _GEN_3844 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_355 & _GEN_3811 : ~(_GEN_1216 & _GEN_355) & _GEN_3811) : _GEN_3811;
  wire        _GEN_3845 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_356 & _GEN_3812 : ~(_GEN_1216 & _GEN_356) & _GEN_3812) : _GEN_3812;
  wire        _GEN_3846 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_357 & _GEN_3813 : ~(_GEN_1216 & _GEN_357) & _GEN_3813) : _GEN_3813;
  wire        _GEN_3847 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_358 & _GEN_3814 : ~(_GEN_1216 & _GEN_358) & _GEN_3814) : _GEN_3814;
  wire        _GEN_3848 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_359 & _GEN_3815 : ~(_GEN_1216 & _GEN_359) & _GEN_3815) : _GEN_3815;
  wire        _GEN_3849 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_360 & _GEN_3816 : ~(_GEN_1216 & _GEN_360) & _GEN_3816) : _GEN_3816;
  wire        _GEN_3850 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_361 & _GEN_3817 : ~(_GEN_1216 & _GEN_361) & _GEN_3817) : _GEN_3817;
  wire        _GEN_3851 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_362 & _GEN_3818 : ~(_GEN_1216 & _GEN_362) & _GEN_3818) : _GEN_3818;
  wire        _GEN_3852 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_363 & _GEN_3819 : ~(_GEN_1216 & _GEN_363) & _GEN_3819) : _GEN_3819;
  wire        _GEN_3853 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_364 & _GEN_3820 : ~(_GEN_1216 & _GEN_364) & _GEN_3820) : _GEN_3820;
  wire        _GEN_3854 = _GEN_1218 ? (_GEN_3823 ? ~_GEN_365 & _GEN_3821 : ~(_GEN_1216 & _GEN_365) & _GEN_3821) : _GEN_3821;
  wire        _GEN_3855 = _GEN_1218 ? (_GEN_3823 ? ~(&lcam_ldq_idx_1) & _GEN_3822 : ~(_GEN_1216 & (&lcam_ldq_idx_1)) & _GEN_3822) : _GEN_3822;
  wire        _GEN_3856 = _GEN_1225 | _GEN_1226;
  wire        _GEN_3857 = _GEN_1223 ? (_GEN_3856 ? (|lcam_ldq_idx_0) & _GEN_3824 : ~(_GEN_1227 & ~(|lcam_ldq_idx_0)) & _GEN_3824) : _GEN_3824;
  wire        _GEN_3858 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_296 & _GEN_3825 : ~(_GEN_1227 & _GEN_296) & _GEN_3825) : _GEN_3825;
  wire        _GEN_3859 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_297 & _GEN_3826 : ~(_GEN_1227 & _GEN_297) & _GEN_3826) : _GEN_3826;
  wire        _GEN_3860 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_298 & _GEN_3827 : ~(_GEN_1227 & _GEN_298) & _GEN_3827) : _GEN_3827;
  wire        _GEN_3861 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_299 & _GEN_3828 : ~(_GEN_1227 & _GEN_299) & _GEN_3828) : _GEN_3828;
  wire        _GEN_3862 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_300 & _GEN_3829 : ~(_GEN_1227 & _GEN_300) & _GEN_3829) : _GEN_3829;
  wire        _GEN_3863 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_301 & _GEN_3830 : ~(_GEN_1227 & _GEN_301) & _GEN_3830) : _GEN_3830;
  wire        _GEN_3864 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_302 & _GEN_3831 : ~(_GEN_1227 & _GEN_302) & _GEN_3831) : _GEN_3831;
  wire        _GEN_3865 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_303 & _GEN_3832 : ~(_GEN_1227 & _GEN_303) & _GEN_3832) : _GEN_3832;
  wire        _GEN_3866 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_304 & _GEN_3833 : ~(_GEN_1227 & _GEN_304) & _GEN_3833) : _GEN_3833;
  wire        _GEN_3867 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_305 & _GEN_3834 : ~(_GEN_1227 & _GEN_305) & _GEN_3834) : _GEN_3834;
  wire        _GEN_3868 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_306 & _GEN_3835 : ~(_GEN_1227 & _GEN_306) & _GEN_3835) : _GEN_3835;
  wire        _GEN_3869 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_307 & _GEN_3836 : ~(_GEN_1227 & _GEN_307) & _GEN_3836) : _GEN_3836;
  wire        _GEN_3870 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_308 & _GEN_3837 : ~(_GEN_1227 & _GEN_308) & _GEN_3837) : _GEN_3837;
  wire        _GEN_3871 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_309 & _GEN_3838 : ~(_GEN_1227 & _GEN_309) & _GEN_3838) : _GEN_3838;
  wire        _GEN_3872 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_310 & _GEN_3839 : ~(_GEN_1227 & _GEN_310) & _GEN_3839) : _GEN_3839;
  wire        _GEN_3873 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_311 & _GEN_3840 : ~(_GEN_1227 & _GEN_311) & _GEN_3840) : _GEN_3840;
  wire        _GEN_3874 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_312 & _GEN_3841 : ~(_GEN_1227 & _GEN_312) & _GEN_3841) : _GEN_3841;
  wire        _GEN_3875 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_313 & _GEN_3842 : ~(_GEN_1227 & _GEN_313) & _GEN_3842) : _GEN_3842;
  wire        _GEN_3876 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_314 & _GEN_3843 : ~(_GEN_1227 & _GEN_314) & _GEN_3843) : _GEN_3843;
  wire        _GEN_3877 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_315 & _GEN_3844 : ~(_GEN_1227 & _GEN_315) & _GEN_3844) : _GEN_3844;
  wire        _GEN_3878 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_316 & _GEN_3845 : ~(_GEN_1227 & _GEN_316) & _GEN_3845) : _GEN_3845;
  wire        _GEN_3879 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_317 & _GEN_3846 : ~(_GEN_1227 & _GEN_317) & _GEN_3846) : _GEN_3846;
  wire        _GEN_3880 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_318 & _GEN_3847 : ~(_GEN_1227 & _GEN_318) & _GEN_3847) : _GEN_3847;
  wire        _GEN_3881 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_319 & _GEN_3848 : ~(_GEN_1227 & _GEN_319) & _GEN_3848) : _GEN_3848;
  wire        _GEN_3882 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_320 & _GEN_3849 : ~(_GEN_1227 & _GEN_320) & _GEN_3849) : _GEN_3849;
  wire        _GEN_3883 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_321 & _GEN_3850 : ~(_GEN_1227 & _GEN_321) & _GEN_3850) : _GEN_3850;
  wire        _GEN_3884 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_322 & _GEN_3851 : ~(_GEN_1227 & _GEN_322) & _GEN_3851) : _GEN_3851;
  wire        _GEN_3885 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_323 & _GEN_3852 : ~(_GEN_1227 & _GEN_323) & _GEN_3852) : _GEN_3852;
  wire        _GEN_3886 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_324 & _GEN_3853 : ~(_GEN_1227 & _GEN_324) & _GEN_3853) : _GEN_3853;
  wire        _GEN_3887 = _GEN_1223 ? (_GEN_3856 ? ~_GEN_325 & _GEN_3854 : ~(_GEN_1227 & _GEN_325) & _GEN_3854) : _GEN_3854;
  wire        _GEN_3888 = _GEN_1223 ? (_GEN_3856 ? ~(&lcam_ldq_idx_0) & _GEN_3855 : ~(_GEN_1227 & (&lcam_ldq_idx_0)) & _GEN_3855) : _GEN_3855;
  wire        _GEN_3889 = _GEN_1231 | _GEN_1232;
  wire        _GEN_3890 = _GEN_1229 ? (_GEN_3889 ? (|lcam_ldq_idx_1) & _GEN_3857 : ~(_GEN_1227 & ~(|lcam_ldq_idx_1)) & _GEN_3857) : _GEN_3857;
  wire        _GEN_3891 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_336 & _GEN_3858 : ~(_GEN_1227 & _GEN_336) & _GEN_3858) : _GEN_3858;
  wire        _GEN_3892 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_337 & _GEN_3859 : ~(_GEN_1227 & _GEN_337) & _GEN_3859) : _GEN_3859;
  wire        _GEN_3893 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_338 & _GEN_3860 : ~(_GEN_1227 & _GEN_338) & _GEN_3860) : _GEN_3860;
  wire        _GEN_3894 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_339 & _GEN_3861 : ~(_GEN_1227 & _GEN_339) & _GEN_3861) : _GEN_3861;
  wire        _GEN_3895 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_340 & _GEN_3862 : ~(_GEN_1227 & _GEN_340) & _GEN_3862) : _GEN_3862;
  wire        _GEN_3896 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_341 & _GEN_3863 : ~(_GEN_1227 & _GEN_341) & _GEN_3863) : _GEN_3863;
  wire        _GEN_3897 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_342 & _GEN_3864 : ~(_GEN_1227 & _GEN_342) & _GEN_3864) : _GEN_3864;
  wire        _GEN_3898 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_343 & _GEN_3865 : ~(_GEN_1227 & _GEN_343) & _GEN_3865) : _GEN_3865;
  wire        _GEN_3899 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_344 & _GEN_3866 : ~(_GEN_1227 & _GEN_344) & _GEN_3866) : _GEN_3866;
  wire        _GEN_3900 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_345 & _GEN_3867 : ~(_GEN_1227 & _GEN_345) & _GEN_3867) : _GEN_3867;
  wire        _GEN_3901 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_346 & _GEN_3868 : ~(_GEN_1227 & _GEN_346) & _GEN_3868) : _GEN_3868;
  wire        _GEN_3902 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_347 & _GEN_3869 : ~(_GEN_1227 & _GEN_347) & _GEN_3869) : _GEN_3869;
  wire        _GEN_3903 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_348 & _GEN_3870 : ~(_GEN_1227 & _GEN_348) & _GEN_3870) : _GEN_3870;
  wire        _GEN_3904 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_349 & _GEN_3871 : ~(_GEN_1227 & _GEN_349) & _GEN_3871) : _GEN_3871;
  wire        _GEN_3905 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_350 & _GEN_3872 : ~(_GEN_1227 & _GEN_350) & _GEN_3872) : _GEN_3872;
  wire        _GEN_3906 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_351 & _GEN_3873 : ~(_GEN_1227 & _GEN_351) & _GEN_3873) : _GEN_3873;
  wire        _GEN_3907 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_352 & _GEN_3874 : ~(_GEN_1227 & _GEN_352) & _GEN_3874) : _GEN_3874;
  wire        _GEN_3908 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_353 & _GEN_3875 : ~(_GEN_1227 & _GEN_353) & _GEN_3875) : _GEN_3875;
  wire        _GEN_3909 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_354 & _GEN_3876 : ~(_GEN_1227 & _GEN_354) & _GEN_3876) : _GEN_3876;
  wire        _GEN_3910 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_355 & _GEN_3877 : ~(_GEN_1227 & _GEN_355) & _GEN_3877) : _GEN_3877;
  wire        _GEN_3911 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_356 & _GEN_3878 : ~(_GEN_1227 & _GEN_356) & _GEN_3878) : _GEN_3878;
  wire        _GEN_3912 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_357 & _GEN_3879 : ~(_GEN_1227 & _GEN_357) & _GEN_3879) : _GEN_3879;
  wire        _GEN_3913 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_358 & _GEN_3880 : ~(_GEN_1227 & _GEN_358) & _GEN_3880) : _GEN_3880;
  wire        _GEN_3914 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_359 & _GEN_3881 : ~(_GEN_1227 & _GEN_359) & _GEN_3881) : _GEN_3881;
  wire        _GEN_3915 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_360 & _GEN_3882 : ~(_GEN_1227 & _GEN_360) & _GEN_3882) : _GEN_3882;
  wire        _GEN_3916 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_361 & _GEN_3883 : ~(_GEN_1227 & _GEN_361) & _GEN_3883) : _GEN_3883;
  wire        _GEN_3917 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_362 & _GEN_3884 : ~(_GEN_1227 & _GEN_362) & _GEN_3884) : _GEN_3884;
  wire        _GEN_3918 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_363 & _GEN_3885 : ~(_GEN_1227 & _GEN_363) & _GEN_3885) : _GEN_3885;
  wire        _GEN_3919 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_364 & _GEN_3886 : ~(_GEN_1227 & _GEN_364) & _GEN_3886) : _GEN_3886;
  wire        _GEN_3920 = _GEN_1229 ? (_GEN_3889 ? ~_GEN_365 & _GEN_3887 : ~(_GEN_1227 & _GEN_365) & _GEN_3887) : _GEN_3887;
  wire        _GEN_3921 = _GEN_1229 ? (_GEN_3889 ? ~(&lcam_ldq_idx_1) & _GEN_3888 : ~(_GEN_1227 & (&lcam_ldq_idx_1)) & _GEN_3888) : _GEN_3888;
  wire        _GEN_3922 = _GEN_1236 | _GEN_1237;
  wire        _GEN_3923 = _GEN_1234 ? (_GEN_3922 ? (|lcam_ldq_idx_0) & _GEN_3890 : ~(_GEN_1238 & ~(|lcam_ldq_idx_0)) & _GEN_3890) : _GEN_3890;
  wire        _GEN_3924 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_296 & _GEN_3891 : ~(_GEN_1238 & _GEN_296) & _GEN_3891) : _GEN_3891;
  wire        _GEN_3925 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_297 & _GEN_3892 : ~(_GEN_1238 & _GEN_297) & _GEN_3892) : _GEN_3892;
  wire        _GEN_3926 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_298 & _GEN_3893 : ~(_GEN_1238 & _GEN_298) & _GEN_3893) : _GEN_3893;
  wire        _GEN_3927 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_299 & _GEN_3894 : ~(_GEN_1238 & _GEN_299) & _GEN_3894) : _GEN_3894;
  wire        _GEN_3928 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_300 & _GEN_3895 : ~(_GEN_1238 & _GEN_300) & _GEN_3895) : _GEN_3895;
  wire        _GEN_3929 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_301 & _GEN_3896 : ~(_GEN_1238 & _GEN_301) & _GEN_3896) : _GEN_3896;
  wire        _GEN_3930 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_302 & _GEN_3897 : ~(_GEN_1238 & _GEN_302) & _GEN_3897) : _GEN_3897;
  wire        _GEN_3931 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_303 & _GEN_3898 : ~(_GEN_1238 & _GEN_303) & _GEN_3898) : _GEN_3898;
  wire        _GEN_3932 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_304 & _GEN_3899 : ~(_GEN_1238 & _GEN_304) & _GEN_3899) : _GEN_3899;
  wire        _GEN_3933 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_305 & _GEN_3900 : ~(_GEN_1238 & _GEN_305) & _GEN_3900) : _GEN_3900;
  wire        _GEN_3934 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_306 & _GEN_3901 : ~(_GEN_1238 & _GEN_306) & _GEN_3901) : _GEN_3901;
  wire        _GEN_3935 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_307 & _GEN_3902 : ~(_GEN_1238 & _GEN_307) & _GEN_3902) : _GEN_3902;
  wire        _GEN_3936 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_308 & _GEN_3903 : ~(_GEN_1238 & _GEN_308) & _GEN_3903) : _GEN_3903;
  wire        _GEN_3937 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_309 & _GEN_3904 : ~(_GEN_1238 & _GEN_309) & _GEN_3904) : _GEN_3904;
  wire        _GEN_3938 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_310 & _GEN_3905 : ~(_GEN_1238 & _GEN_310) & _GEN_3905) : _GEN_3905;
  wire        _GEN_3939 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_311 & _GEN_3906 : ~(_GEN_1238 & _GEN_311) & _GEN_3906) : _GEN_3906;
  wire        _GEN_3940 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_312 & _GEN_3907 : ~(_GEN_1238 & _GEN_312) & _GEN_3907) : _GEN_3907;
  wire        _GEN_3941 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_313 & _GEN_3908 : ~(_GEN_1238 & _GEN_313) & _GEN_3908) : _GEN_3908;
  wire        _GEN_3942 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_314 & _GEN_3909 : ~(_GEN_1238 & _GEN_314) & _GEN_3909) : _GEN_3909;
  wire        _GEN_3943 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_315 & _GEN_3910 : ~(_GEN_1238 & _GEN_315) & _GEN_3910) : _GEN_3910;
  wire        _GEN_3944 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_316 & _GEN_3911 : ~(_GEN_1238 & _GEN_316) & _GEN_3911) : _GEN_3911;
  wire        _GEN_3945 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_317 & _GEN_3912 : ~(_GEN_1238 & _GEN_317) & _GEN_3912) : _GEN_3912;
  wire        _GEN_3946 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_318 & _GEN_3913 : ~(_GEN_1238 & _GEN_318) & _GEN_3913) : _GEN_3913;
  wire        _GEN_3947 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_319 & _GEN_3914 : ~(_GEN_1238 & _GEN_319) & _GEN_3914) : _GEN_3914;
  wire        _GEN_3948 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_320 & _GEN_3915 : ~(_GEN_1238 & _GEN_320) & _GEN_3915) : _GEN_3915;
  wire        _GEN_3949 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_321 & _GEN_3916 : ~(_GEN_1238 & _GEN_321) & _GEN_3916) : _GEN_3916;
  wire        _GEN_3950 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_322 & _GEN_3917 : ~(_GEN_1238 & _GEN_322) & _GEN_3917) : _GEN_3917;
  wire        _GEN_3951 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_323 & _GEN_3918 : ~(_GEN_1238 & _GEN_323) & _GEN_3918) : _GEN_3918;
  wire        _GEN_3952 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_324 & _GEN_3919 : ~(_GEN_1238 & _GEN_324) & _GEN_3919) : _GEN_3919;
  wire        _GEN_3953 = _GEN_1234 ? (_GEN_3922 ? ~_GEN_325 & _GEN_3920 : ~(_GEN_1238 & _GEN_325) & _GEN_3920) : _GEN_3920;
  wire        _GEN_3954 = _GEN_1234 ? (_GEN_3922 ? ~(&lcam_ldq_idx_0) & _GEN_3921 : ~(_GEN_1238 & (&lcam_ldq_idx_0)) & _GEN_3921) : _GEN_3921;
  wire        _GEN_3955 = _GEN_1242 | _GEN_1243;
  wire        _GEN_3956 = _GEN_1240 ? (_GEN_3955 ? (|lcam_ldq_idx_1) & _GEN_3923 : ~(_GEN_1238 & ~(|lcam_ldq_idx_1)) & _GEN_3923) : _GEN_3923;
  wire        _GEN_3957 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_336 & _GEN_3924 : ~(_GEN_1238 & _GEN_336) & _GEN_3924) : _GEN_3924;
  wire        _GEN_3958 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_337 & _GEN_3925 : ~(_GEN_1238 & _GEN_337) & _GEN_3925) : _GEN_3925;
  wire        _GEN_3959 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_338 & _GEN_3926 : ~(_GEN_1238 & _GEN_338) & _GEN_3926) : _GEN_3926;
  wire        _GEN_3960 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_339 & _GEN_3927 : ~(_GEN_1238 & _GEN_339) & _GEN_3927) : _GEN_3927;
  wire        _GEN_3961 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_340 & _GEN_3928 : ~(_GEN_1238 & _GEN_340) & _GEN_3928) : _GEN_3928;
  wire        _GEN_3962 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_341 & _GEN_3929 : ~(_GEN_1238 & _GEN_341) & _GEN_3929) : _GEN_3929;
  wire        _GEN_3963 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_342 & _GEN_3930 : ~(_GEN_1238 & _GEN_342) & _GEN_3930) : _GEN_3930;
  wire        _GEN_3964 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_343 & _GEN_3931 : ~(_GEN_1238 & _GEN_343) & _GEN_3931) : _GEN_3931;
  wire        _GEN_3965 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_344 & _GEN_3932 : ~(_GEN_1238 & _GEN_344) & _GEN_3932) : _GEN_3932;
  wire        _GEN_3966 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_345 & _GEN_3933 : ~(_GEN_1238 & _GEN_345) & _GEN_3933) : _GEN_3933;
  wire        _GEN_3967 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_346 & _GEN_3934 : ~(_GEN_1238 & _GEN_346) & _GEN_3934) : _GEN_3934;
  wire        _GEN_3968 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_347 & _GEN_3935 : ~(_GEN_1238 & _GEN_347) & _GEN_3935) : _GEN_3935;
  wire        _GEN_3969 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_348 & _GEN_3936 : ~(_GEN_1238 & _GEN_348) & _GEN_3936) : _GEN_3936;
  wire        _GEN_3970 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_349 & _GEN_3937 : ~(_GEN_1238 & _GEN_349) & _GEN_3937) : _GEN_3937;
  wire        _GEN_3971 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_350 & _GEN_3938 : ~(_GEN_1238 & _GEN_350) & _GEN_3938) : _GEN_3938;
  wire        _GEN_3972 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_351 & _GEN_3939 : ~(_GEN_1238 & _GEN_351) & _GEN_3939) : _GEN_3939;
  wire        _GEN_3973 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_352 & _GEN_3940 : ~(_GEN_1238 & _GEN_352) & _GEN_3940) : _GEN_3940;
  wire        _GEN_3974 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_353 & _GEN_3941 : ~(_GEN_1238 & _GEN_353) & _GEN_3941) : _GEN_3941;
  wire        _GEN_3975 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_354 & _GEN_3942 : ~(_GEN_1238 & _GEN_354) & _GEN_3942) : _GEN_3942;
  wire        _GEN_3976 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_355 & _GEN_3943 : ~(_GEN_1238 & _GEN_355) & _GEN_3943) : _GEN_3943;
  wire        _GEN_3977 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_356 & _GEN_3944 : ~(_GEN_1238 & _GEN_356) & _GEN_3944) : _GEN_3944;
  wire        _GEN_3978 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_357 & _GEN_3945 : ~(_GEN_1238 & _GEN_357) & _GEN_3945) : _GEN_3945;
  wire        _GEN_3979 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_358 & _GEN_3946 : ~(_GEN_1238 & _GEN_358) & _GEN_3946) : _GEN_3946;
  wire        _GEN_3980 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_359 & _GEN_3947 : ~(_GEN_1238 & _GEN_359) & _GEN_3947) : _GEN_3947;
  wire        _GEN_3981 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_360 & _GEN_3948 : ~(_GEN_1238 & _GEN_360) & _GEN_3948) : _GEN_3948;
  wire        _GEN_3982 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_361 & _GEN_3949 : ~(_GEN_1238 & _GEN_361) & _GEN_3949) : _GEN_3949;
  wire        _GEN_3983 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_362 & _GEN_3950 : ~(_GEN_1238 & _GEN_362) & _GEN_3950) : _GEN_3950;
  wire        _GEN_3984 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_363 & _GEN_3951 : ~(_GEN_1238 & _GEN_363) & _GEN_3951) : _GEN_3951;
  wire        _GEN_3985 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_364 & _GEN_3952 : ~(_GEN_1238 & _GEN_364) & _GEN_3952) : _GEN_3952;
  wire        _GEN_3986 = _GEN_1240 ? (_GEN_3955 ? ~_GEN_365 & _GEN_3953 : ~(_GEN_1238 & _GEN_365) & _GEN_3953) : _GEN_3953;
  wire        _GEN_3987 = _GEN_1240 ? (_GEN_3955 ? ~(&lcam_ldq_idx_1) & _GEN_3954 : ~(_GEN_1238 & (&lcam_ldq_idx_1)) & _GEN_3954) : _GEN_3954;
  wire        _GEN_3988 = _GEN_1247 | _GEN_1248;
  wire        _GEN_3989 = _GEN_1245 ? (_GEN_3988 ? (|lcam_ldq_idx_0) & _GEN_3956 : ~(_GEN_1249 & ~(|lcam_ldq_idx_0)) & _GEN_3956) : _GEN_3956;
  wire        _GEN_3990 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_296 & _GEN_3957 : ~(_GEN_1249 & _GEN_296) & _GEN_3957) : _GEN_3957;
  wire        _GEN_3991 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_297 & _GEN_3958 : ~(_GEN_1249 & _GEN_297) & _GEN_3958) : _GEN_3958;
  wire        _GEN_3992 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_298 & _GEN_3959 : ~(_GEN_1249 & _GEN_298) & _GEN_3959) : _GEN_3959;
  wire        _GEN_3993 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_299 & _GEN_3960 : ~(_GEN_1249 & _GEN_299) & _GEN_3960) : _GEN_3960;
  wire        _GEN_3994 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_300 & _GEN_3961 : ~(_GEN_1249 & _GEN_300) & _GEN_3961) : _GEN_3961;
  wire        _GEN_3995 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_301 & _GEN_3962 : ~(_GEN_1249 & _GEN_301) & _GEN_3962) : _GEN_3962;
  wire        _GEN_3996 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_302 & _GEN_3963 : ~(_GEN_1249 & _GEN_302) & _GEN_3963) : _GEN_3963;
  wire        _GEN_3997 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_303 & _GEN_3964 : ~(_GEN_1249 & _GEN_303) & _GEN_3964) : _GEN_3964;
  wire        _GEN_3998 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_304 & _GEN_3965 : ~(_GEN_1249 & _GEN_304) & _GEN_3965) : _GEN_3965;
  wire        _GEN_3999 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_305 & _GEN_3966 : ~(_GEN_1249 & _GEN_305) & _GEN_3966) : _GEN_3966;
  wire        _GEN_4000 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_306 & _GEN_3967 : ~(_GEN_1249 & _GEN_306) & _GEN_3967) : _GEN_3967;
  wire        _GEN_4001 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_307 & _GEN_3968 : ~(_GEN_1249 & _GEN_307) & _GEN_3968) : _GEN_3968;
  wire        _GEN_4002 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_308 & _GEN_3969 : ~(_GEN_1249 & _GEN_308) & _GEN_3969) : _GEN_3969;
  wire        _GEN_4003 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_309 & _GEN_3970 : ~(_GEN_1249 & _GEN_309) & _GEN_3970) : _GEN_3970;
  wire        _GEN_4004 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_310 & _GEN_3971 : ~(_GEN_1249 & _GEN_310) & _GEN_3971) : _GEN_3971;
  wire        _GEN_4005 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_311 & _GEN_3972 : ~(_GEN_1249 & _GEN_311) & _GEN_3972) : _GEN_3972;
  wire        _GEN_4006 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_312 & _GEN_3973 : ~(_GEN_1249 & _GEN_312) & _GEN_3973) : _GEN_3973;
  wire        _GEN_4007 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_313 & _GEN_3974 : ~(_GEN_1249 & _GEN_313) & _GEN_3974) : _GEN_3974;
  wire        _GEN_4008 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_314 & _GEN_3975 : ~(_GEN_1249 & _GEN_314) & _GEN_3975) : _GEN_3975;
  wire        _GEN_4009 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_315 & _GEN_3976 : ~(_GEN_1249 & _GEN_315) & _GEN_3976) : _GEN_3976;
  wire        _GEN_4010 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_316 & _GEN_3977 : ~(_GEN_1249 & _GEN_316) & _GEN_3977) : _GEN_3977;
  wire        _GEN_4011 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_317 & _GEN_3978 : ~(_GEN_1249 & _GEN_317) & _GEN_3978) : _GEN_3978;
  wire        _GEN_4012 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_318 & _GEN_3979 : ~(_GEN_1249 & _GEN_318) & _GEN_3979) : _GEN_3979;
  wire        _GEN_4013 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_319 & _GEN_3980 : ~(_GEN_1249 & _GEN_319) & _GEN_3980) : _GEN_3980;
  wire        _GEN_4014 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_320 & _GEN_3981 : ~(_GEN_1249 & _GEN_320) & _GEN_3981) : _GEN_3981;
  wire        _GEN_4015 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_321 & _GEN_3982 : ~(_GEN_1249 & _GEN_321) & _GEN_3982) : _GEN_3982;
  wire        _GEN_4016 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_322 & _GEN_3983 : ~(_GEN_1249 & _GEN_322) & _GEN_3983) : _GEN_3983;
  wire        _GEN_4017 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_323 & _GEN_3984 : ~(_GEN_1249 & _GEN_323) & _GEN_3984) : _GEN_3984;
  wire        _GEN_4018 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_324 & _GEN_3985 : ~(_GEN_1249 & _GEN_324) & _GEN_3985) : _GEN_3985;
  wire        _GEN_4019 = _GEN_1245 ? (_GEN_3988 ? ~_GEN_325 & _GEN_3986 : ~(_GEN_1249 & _GEN_325) & _GEN_3986) : _GEN_3986;
  wire        _GEN_4020 = _GEN_1245 ? (_GEN_3988 ? ~(&lcam_ldq_idx_0) & _GEN_3987 : ~(_GEN_1249 & (&lcam_ldq_idx_0)) & _GEN_3987) : _GEN_3987;
  wire        _GEN_4021 = _GEN_1253 | _GEN_1254;
  wire        _GEN_4022 = _GEN_1251 ? (_GEN_4021 ? (|lcam_ldq_idx_1) & _GEN_3989 : ~(_GEN_1249 & ~(|lcam_ldq_idx_1)) & _GEN_3989) : _GEN_3989;
  wire        _GEN_4023 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_336 & _GEN_3990 : ~(_GEN_1249 & _GEN_336) & _GEN_3990) : _GEN_3990;
  wire        _GEN_4024 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_337 & _GEN_3991 : ~(_GEN_1249 & _GEN_337) & _GEN_3991) : _GEN_3991;
  wire        _GEN_4025 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_338 & _GEN_3992 : ~(_GEN_1249 & _GEN_338) & _GEN_3992) : _GEN_3992;
  wire        _GEN_4026 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_339 & _GEN_3993 : ~(_GEN_1249 & _GEN_339) & _GEN_3993) : _GEN_3993;
  wire        _GEN_4027 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_340 & _GEN_3994 : ~(_GEN_1249 & _GEN_340) & _GEN_3994) : _GEN_3994;
  wire        _GEN_4028 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_341 & _GEN_3995 : ~(_GEN_1249 & _GEN_341) & _GEN_3995) : _GEN_3995;
  wire        _GEN_4029 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_342 & _GEN_3996 : ~(_GEN_1249 & _GEN_342) & _GEN_3996) : _GEN_3996;
  wire        _GEN_4030 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_343 & _GEN_3997 : ~(_GEN_1249 & _GEN_343) & _GEN_3997) : _GEN_3997;
  wire        _GEN_4031 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_344 & _GEN_3998 : ~(_GEN_1249 & _GEN_344) & _GEN_3998) : _GEN_3998;
  wire        _GEN_4032 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_345 & _GEN_3999 : ~(_GEN_1249 & _GEN_345) & _GEN_3999) : _GEN_3999;
  wire        _GEN_4033 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_346 & _GEN_4000 : ~(_GEN_1249 & _GEN_346) & _GEN_4000) : _GEN_4000;
  wire        _GEN_4034 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_347 & _GEN_4001 : ~(_GEN_1249 & _GEN_347) & _GEN_4001) : _GEN_4001;
  wire        _GEN_4035 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_348 & _GEN_4002 : ~(_GEN_1249 & _GEN_348) & _GEN_4002) : _GEN_4002;
  wire        _GEN_4036 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_349 & _GEN_4003 : ~(_GEN_1249 & _GEN_349) & _GEN_4003) : _GEN_4003;
  wire        _GEN_4037 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_350 & _GEN_4004 : ~(_GEN_1249 & _GEN_350) & _GEN_4004) : _GEN_4004;
  wire        _GEN_4038 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_351 & _GEN_4005 : ~(_GEN_1249 & _GEN_351) & _GEN_4005) : _GEN_4005;
  wire        _GEN_4039 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_352 & _GEN_4006 : ~(_GEN_1249 & _GEN_352) & _GEN_4006) : _GEN_4006;
  wire        _GEN_4040 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_353 & _GEN_4007 : ~(_GEN_1249 & _GEN_353) & _GEN_4007) : _GEN_4007;
  wire        _GEN_4041 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_354 & _GEN_4008 : ~(_GEN_1249 & _GEN_354) & _GEN_4008) : _GEN_4008;
  wire        _GEN_4042 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_355 & _GEN_4009 : ~(_GEN_1249 & _GEN_355) & _GEN_4009) : _GEN_4009;
  wire        _GEN_4043 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_356 & _GEN_4010 : ~(_GEN_1249 & _GEN_356) & _GEN_4010) : _GEN_4010;
  wire        _GEN_4044 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_357 & _GEN_4011 : ~(_GEN_1249 & _GEN_357) & _GEN_4011) : _GEN_4011;
  wire        _GEN_4045 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_358 & _GEN_4012 : ~(_GEN_1249 & _GEN_358) & _GEN_4012) : _GEN_4012;
  wire        _GEN_4046 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_359 & _GEN_4013 : ~(_GEN_1249 & _GEN_359) & _GEN_4013) : _GEN_4013;
  wire        _GEN_4047 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_360 & _GEN_4014 : ~(_GEN_1249 & _GEN_360) & _GEN_4014) : _GEN_4014;
  wire        _GEN_4048 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_361 & _GEN_4015 : ~(_GEN_1249 & _GEN_361) & _GEN_4015) : _GEN_4015;
  wire        _GEN_4049 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_362 & _GEN_4016 : ~(_GEN_1249 & _GEN_362) & _GEN_4016) : _GEN_4016;
  wire        _GEN_4050 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_363 & _GEN_4017 : ~(_GEN_1249 & _GEN_363) & _GEN_4017) : _GEN_4017;
  wire        _GEN_4051 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_364 & _GEN_4018 : ~(_GEN_1249 & _GEN_364) & _GEN_4018) : _GEN_4018;
  wire        _GEN_4052 = _GEN_1251 ? (_GEN_4021 ? ~_GEN_365 & _GEN_4019 : ~(_GEN_1249 & _GEN_365) & _GEN_4019) : _GEN_4019;
  wire        _GEN_4053 = _GEN_1251 ? (_GEN_4021 ? ~(&lcam_ldq_idx_1) & _GEN_4020 : ~(_GEN_1249 & (&lcam_ldq_idx_1)) & _GEN_4020) : _GEN_4020;
  wire        _GEN_4054 = _GEN_1258 | _GEN_1259;
  wire        _GEN_4055 = _GEN_1256 ? (_GEN_4054 ? (|lcam_ldq_idx_0) & _GEN_4022 : ~(_GEN_1260 & ~(|lcam_ldq_idx_0)) & _GEN_4022) : _GEN_4022;
  wire        _GEN_4056 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_296 & _GEN_4023 : ~(_GEN_1260 & _GEN_296) & _GEN_4023) : _GEN_4023;
  wire        _GEN_4057 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_297 & _GEN_4024 : ~(_GEN_1260 & _GEN_297) & _GEN_4024) : _GEN_4024;
  wire        _GEN_4058 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_298 & _GEN_4025 : ~(_GEN_1260 & _GEN_298) & _GEN_4025) : _GEN_4025;
  wire        _GEN_4059 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_299 & _GEN_4026 : ~(_GEN_1260 & _GEN_299) & _GEN_4026) : _GEN_4026;
  wire        _GEN_4060 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_300 & _GEN_4027 : ~(_GEN_1260 & _GEN_300) & _GEN_4027) : _GEN_4027;
  wire        _GEN_4061 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_301 & _GEN_4028 : ~(_GEN_1260 & _GEN_301) & _GEN_4028) : _GEN_4028;
  wire        _GEN_4062 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_302 & _GEN_4029 : ~(_GEN_1260 & _GEN_302) & _GEN_4029) : _GEN_4029;
  wire        _GEN_4063 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_303 & _GEN_4030 : ~(_GEN_1260 & _GEN_303) & _GEN_4030) : _GEN_4030;
  wire        _GEN_4064 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_304 & _GEN_4031 : ~(_GEN_1260 & _GEN_304) & _GEN_4031) : _GEN_4031;
  wire        _GEN_4065 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_305 & _GEN_4032 : ~(_GEN_1260 & _GEN_305) & _GEN_4032) : _GEN_4032;
  wire        _GEN_4066 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_306 & _GEN_4033 : ~(_GEN_1260 & _GEN_306) & _GEN_4033) : _GEN_4033;
  wire        _GEN_4067 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_307 & _GEN_4034 : ~(_GEN_1260 & _GEN_307) & _GEN_4034) : _GEN_4034;
  wire        _GEN_4068 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_308 & _GEN_4035 : ~(_GEN_1260 & _GEN_308) & _GEN_4035) : _GEN_4035;
  wire        _GEN_4069 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_309 & _GEN_4036 : ~(_GEN_1260 & _GEN_309) & _GEN_4036) : _GEN_4036;
  wire        _GEN_4070 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_310 & _GEN_4037 : ~(_GEN_1260 & _GEN_310) & _GEN_4037) : _GEN_4037;
  wire        _GEN_4071 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_311 & _GEN_4038 : ~(_GEN_1260 & _GEN_311) & _GEN_4038) : _GEN_4038;
  wire        _GEN_4072 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_312 & _GEN_4039 : ~(_GEN_1260 & _GEN_312) & _GEN_4039) : _GEN_4039;
  wire        _GEN_4073 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_313 & _GEN_4040 : ~(_GEN_1260 & _GEN_313) & _GEN_4040) : _GEN_4040;
  wire        _GEN_4074 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_314 & _GEN_4041 : ~(_GEN_1260 & _GEN_314) & _GEN_4041) : _GEN_4041;
  wire        _GEN_4075 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_315 & _GEN_4042 : ~(_GEN_1260 & _GEN_315) & _GEN_4042) : _GEN_4042;
  wire        _GEN_4076 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_316 & _GEN_4043 : ~(_GEN_1260 & _GEN_316) & _GEN_4043) : _GEN_4043;
  wire        _GEN_4077 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_317 & _GEN_4044 : ~(_GEN_1260 & _GEN_317) & _GEN_4044) : _GEN_4044;
  wire        _GEN_4078 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_318 & _GEN_4045 : ~(_GEN_1260 & _GEN_318) & _GEN_4045) : _GEN_4045;
  wire        _GEN_4079 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_319 & _GEN_4046 : ~(_GEN_1260 & _GEN_319) & _GEN_4046) : _GEN_4046;
  wire        _GEN_4080 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_320 & _GEN_4047 : ~(_GEN_1260 & _GEN_320) & _GEN_4047) : _GEN_4047;
  wire        _GEN_4081 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_321 & _GEN_4048 : ~(_GEN_1260 & _GEN_321) & _GEN_4048) : _GEN_4048;
  wire        _GEN_4082 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_322 & _GEN_4049 : ~(_GEN_1260 & _GEN_322) & _GEN_4049) : _GEN_4049;
  wire        _GEN_4083 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_323 & _GEN_4050 : ~(_GEN_1260 & _GEN_323) & _GEN_4050) : _GEN_4050;
  wire        _GEN_4084 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_324 & _GEN_4051 : ~(_GEN_1260 & _GEN_324) & _GEN_4051) : _GEN_4051;
  wire        _GEN_4085 = _GEN_1256 ? (_GEN_4054 ? ~_GEN_325 & _GEN_4052 : ~(_GEN_1260 & _GEN_325) & _GEN_4052) : _GEN_4052;
  wire        _GEN_4086 = _GEN_1256 ? (_GEN_4054 ? ~(&lcam_ldq_idx_0) & _GEN_4053 : ~(_GEN_1260 & (&lcam_ldq_idx_0)) & _GEN_4053) : _GEN_4053;
  wire        _GEN_4087 = _GEN_1264 | _GEN_1265;
  wire        _GEN_4088 = _GEN_1262 ? (_GEN_4087 ? (|lcam_ldq_idx_1) & _GEN_4055 : ~(_GEN_1260 & ~(|lcam_ldq_idx_1)) & _GEN_4055) : _GEN_4055;
  wire        _GEN_4089 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_336 & _GEN_4056 : ~(_GEN_1260 & _GEN_336) & _GEN_4056) : _GEN_4056;
  wire        _GEN_4090 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_337 & _GEN_4057 : ~(_GEN_1260 & _GEN_337) & _GEN_4057) : _GEN_4057;
  wire        _GEN_4091 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_338 & _GEN_4058 : ~(_GEN_1260 & _GEN_338) & _GEN_4058) : _GEN_4058;
  wire        _GEN_4092 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_339 & _GEN_4059 : ~(_GEN_1260 & _GEN_339) & _GEN_4059) : _GEN_4059;
  wire        _GEN_4093 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_340 & _GEN_4060 : ~(_GEN_1260 & _GEN_340) & _GEN_4060) : _GEN_4060;
  wire        _GEN_4094 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_341 & _GEN_4061 : ~(_GEN_1260 & _GEN_341) & _GEN_4061) : _GEN_4061;
  wire        _GEN_4095 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_342 & _GEN_4062 : ~(_GEN_1260 & _GEN_342) & _GEN_4062) : _GEN_4062;
  wire        _GEN_4096 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_343 & _GEN_4063 : ~(_GEN_1260 & _GEN_343) & _GEN_4063) : _GEN_4063;
  wire        _GEN_4097 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_344 & _GEN_4064 : ~(_GEN_1260 & _GEN_344) & _GEN_4064) : _GEN_4064;
  wire        _GEN_4098 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_345 & _GEN_4065 : ~(_GEN_1260 & _GEN_345) & _GEN_4065) : _GEN_4065;
  wire        _GEN_4099 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_346 & _GEN_4066 : ~(_GEN_1260 & _GEN_346) & _GEN_4066) : _GEN_4066;
  wire        _GEN_4100 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_347 & _GEN_4067 : ~(_GEN_1260 & _GEN_347) & _GEN_4067) : _GEN_4067;
  wire        _GEN_4101 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_348 & _GEN_4068 : ~(_GEN_1260 & _GEN_348) & _GEN_4068) : _GEN_4068;
  wire        _GEN_4102 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_349 & _GEN_4069 : ~(_GEN_1260 & _GEN_349) & _GEN_4069) : _GEN_4069;
  wire        _GEN_4103 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_350 & _GEN_4070 : ~(_GEN_1260 & _GEN_350) & _GEN_4070) : _GEN_4070;
  wire        _GEN_4104 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_351 & _GEN_4071 : ~(_GEN_1260 & _GEN_351) & _GEN_4071) : _GEN_4071;
  wire        _GEN_4105 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_352 & _GEN_4072 : ~(_GEN_1260 & _GEN_352) & _GEN_4072) : _GEN_4072;
  wire        _GEN_4106 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_353 & _GEN_4073 : ~(_GEN_1260 & _GEN_353) & _GEN_4073) : _GEN_4073;
  wire        _GEN_4107 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_354 & _GEN_4074 : ~(_GEN_1260 & _GEN_354) & _GEN_4074) : _GEN_4074;
  wire        _GEN_4108 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_355 & _GEN_4075 : ~(_GEN_1260 & _GEN_355) & _GEN_4075) : _GEN_4075;
  wire        _GEN_4109 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_356 & _GEN_4076 : ~(_GEN_1260 & _GEN_356) & _GEN_4076) : _GEN_4076;
  wire        _GEN_4110 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_357 & _GEN_4077 : ~(_GEN_1260 & _GEN_357) & _GEN_4077) : _GEN_4077;
  wire        _GEN_4111 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_358 & _GEN_4078 : ~(_GEN_1260 & _GEN_358) & _GEN_4078) : _GEN_4078;
  wire        _GEN_4112 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_359 & _GEN_4079 : ~(_GEN_1260 & _GEN_359) & _GEN_4079) : _GEN_4079;
  wire        _GEN_4113 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_360 & _GEN_4080 : ~(_GEN_1260 & _GEN_360) & _GEN_4080) : _GEN_4080;
  wire        _GEN_4114 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_361 & _GEN_4081 : ~(_GEN_1260 & _GEN_361) & _GEN_4081) : _GEN_4081;
  wire        _GEN_4115 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_362 & _GEN_4082 : ~(_GEN_1260 & _GEN_362) & _GEN_4082) : _GEN_4082;
  wire        _GEN_4116 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_363 & _GEN_4083 : ~(_GEN_1260 & _GEN_363) & _GEN_4083) : _GEN_4083;
  wire        _GEN_4117 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_364 & _GEN_4084 : ~(_GEN_1260 & _GEN_364) & _GEN_4084) : _GEN_4084;
  wire        _GEN_4118 = _GEN_1262 ? (_GEN_4087 ? ~_GEN_365 & _GEN_4085 : ~(_GEN_1260 & _GEN_365) & _GEN_4085) : _GEN_4085;
  wire        _GEN_4119 = _GEN_1262 ? (_GEN_4087 ? ~(&lcam_ldq_idx_1) & _GEN_4086 : ~(_GEN_1260 & (&lcam_ldq_idx_1)) & _GEN_4086) : _GEN_4086;
  wire        _GEN_4120 = _GEN_1269 | _GEN_1270;
  wire        _GEN_4121 = _GEN_1267 ? (_GEN_4120 ? (|lcam_ldq_idx_0) & _GEN_4088 : ~(_GEN_1271 & ~(|lcam_ldq_idx_0)) & _GEN_4088) : _GEN_4088;
  wire        _GEN_4122 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_296 & _GEN_4089 : ~(_GEN_1271 & _GEN_296) & _GEN_4089) : _GEN_4089;
  wire        _GEN_4123 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_297 & _GEN_4090 : ~(_GEN_1271 & _GEN_297) & _GEN_4090) : _GEN_4090;
  wire        _GEN_4124 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_298 & _GEN_4091 : ~(_GEN_1271 & _GEN_298) & _GEN_4091) : _GEN_4091;
  wire        _GEN_4125 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_299 & _GEN_4092 : ~(_GEN_1271 & _GEN_299) & _GEN_4092) : _GEN_4092;
  wire        _GEN_4126 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_300 & _GEN_4093 : ~(_GEN_1271 & _GEN_300) & _GEN_4093) : _GEN_4093;
  wire        _GEN_4127 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_301 & _GEN_4094 : ~(_GEN_1271 & _GEN_301) & _GEN_4094) : _GEN_4094;
  wire        _GEN_4128 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_302 & _GEN_4095 : ~(_GEN_1271 & _GEN_302) & _GEN_4095) : _GEN_4095;
  wire        _GEN_4129 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_303 & _GEN_4096 : ~(_GEN_1271 & _GEN_303) & _GEN_4096) : _GEN_4096;
  wire        _GEN_4130 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_304 & _GEN_4097 : ~(_GEN_1271 & _GEN_304) & _GEN_4097) : _GEN_4097;
  wire        _GEN_4131 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_305 & _GEN_4098 : ~(_GEN_1271 & _GEN_305) & _GEN_4098) : _GEN_4098;
  wire        _GEN_4132 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_306 & _GEN_4099 : ~(_GEN_1271 & _GEN_306) & _GEN_4099) : _GEN_4099;
  wire        _GEN_4133 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_307 & _GEN_4100 : ~(_GEN_1271 & _GEN_307) & _GEN_4100) : _GEN_4100;
  wire        _GEN_4134 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_308 & _GEN_4101 : ~(_GEN_1271 & _GEN_308) & _GEN_4101) : _GEN_4101;
  wire        _GEN_4135 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_309 & _GEN_4102 : ~(_GEN_1271 & _GEN_309) & _GEN_4102) : _GEN_4102;
  wire        _GEN_4136 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_310 & _GEN_4103 : ~(_GEN_1271 & _GEN_310) & _GEN_4103) : _GEN_4103;
  wire        _GEN_4137 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_311 & _GEN_4104 : ~(_GEN_1271 & _GEN_311) & _GEN_4104) : _GEN_4104;
  wire        _GEN_4138 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_312 & _GEN_4105 : ~(_GEN_1271 & _GEN_312) & _GEN_4105) : _GEN_4105;
  wire        _GEN_4139 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_313 & _GEN_4106 : ~(_GEN_1271 & _GEN_313) & _GEN_4106) : _GEN_4106;
  wire        _GEN_4140 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_314 & _GEN_4107 : ~(_GEN_1271 & _GEN_314) & _GEN_4107) : _GEN_4107;
  wire        _GEN_4141 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_315 & _GEN_4108 : ~(_GEN_1271 & _GEN_315) & _GEN_4108) : _GEN_4108;
  wire        _GEN_4142 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_316 & _GEN_4109 : ~(_GEN_1271 & _GEN_316) & _GEN_4109) : _GEN_4109;
  wire        _GEN_4143 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_317 & _GEN_4110 : ~(_GEN_1271 & _GEN_317) & _GEN_4110) : _GEN_4110;
  wire        _GEN_4144 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_318 & _GEN_4111 : ~(_GEN_1271 & _GEN_318) & _GEN_4111) : _GEN_4111;
  wire        _GEN_4145 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_319 & _GEN_4112 : ~(_GEN_1271 & _GEN_319) & _GEN_4112) : _GEN_4112;
  wire        _GEN_4146 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_320 & _GEN_4113 : ~(_GEN_1271 & _GEN_320) & _GEN_4113) : _GEN_4113;
  wire        _GEN_4147 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_321 & _GEN_4114 : ~(_GEN_1271 & _GEN_321) & _GEN_4114) : _GEN_4114;
  wire        _GEN_4148 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_322 & _GEN_4115 : ~(_GEN_1271 & _GEN_322) & _GEN_4115) : _GEN_4115;
  wire        _GEN_4149 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_323 & _GEN_4116 : ~(_GEN_1271 & _GEN_323) & _GEN_4116) : _GEN_4116;
  wire        _GEN_4150 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_324 & _GEN_4117 : ~(_GEN_1271 & _GEN_324) & _GEN_4117) : _GEN_4117;
  wire        _GEN_4151 = _GEN_1267 ? (_GEN_4120 ? ~_GEN_325 & _GEN_4118 : ~(_GEN_1271 & _GEN_325) & _GEN_4118) : _GEN_4118;
  wire        _GEN_4152 = _GEN_1267 ? (_GEN_4120 ? ~(&lcam_ldq_idx_0) & _GEN_4119 : ~(_GEN_1271 & (&lcam_ldq_idx_0)) & _GEN_4119) : _GEN_4119;
  wire        _GEN_4153 = _GEN_1275 | _GEN_1276;
  wire        _GEN_4154 = _GEN_1273 ? (_GEN_4153 ? (|lcam_ldq_idx_1) & _GEN_4121 : ~(_GEN_1271 & ~(|lcam_ldq_idx_1)) & _GEN_4121) : _GEN_4121;
  wire        _GEN_4155 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_336 & _GEN_4122 : ~(_GEN_1271 & _GEN_336) & _GEN_4122) : _GEN_4122;
  wire        _GEN_4156 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_337 & _GEN_4123 : ~(_GEN_1271 & _GEN_337) & _GEN_4123) : _GEN_4123;
  wire        _GEN_4157 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_338 & _GEN_4124 : ~(_GEN_1271 & _GEN_338) & _GEN_4124) : _GEN_4124;
  wire        _GEN_4158 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_339 & _GEN_4125 : ~(_GEN_1271 & _GEN_339) & _GEN_4125) : _GEN_4125;
  wire        _GEN_4159 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_340 & _GEN_4126 : ~(_GEN_1271 & _GEN_340) & _GEN_4126) : _GEN_4126;
  wire        _GEN_4160 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_341 & _GEN_4127 : ~(_GEN_1271 & _GEN_341) & _GEN_4127) : _GEN_4127;
  wire        _GEN_4161 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_342 & _GEN_4128 : ~(_GEN_1271 & _GEN_342) & _GEN_4128) : _GEN_4128;
  wire        _GEN_4162 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_343 & _GEN_4129 : ~(_GEN_1271 & _GEN_343) & _GEN_4129) : _GEN_4129;
  wire        _GEN_4163 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_344 & _GEN_4130 : ~(_GEN_1271 & _GEN_344) & _GEN_4130) : _GEN_4130;
  wire        _GEN_4164 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_345 & _GEN_4131 : ~(_GEN_1271 & _GEN_345) & _GEN_4131) : _GEN_4131;
  wire        _GEN_4165 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_346 & _GEN_4132 : ~(_GEN_1271 & _GEN_346) & _GEN_4132) : _GEN_4132;
  wire        _GEN_4166 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_347 & _GEN_4133 : ~(_GEN_1271 & _GEN_347) & _GEN_4133) : _GEN_4133;
  wire        _GEN_4167 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_348 & _GEN_4134 : ~(_GEN_1271 & _GEN_348) & _GEN_4134) : _GEN_4134;
  wire        _GEN_4168 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_349 & _GEN_4135 : ~(_GEN_1271 & _GEN_349) & _GEN_4135) : _GEN_4135;
  wire        _GEN_4169 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_350 & _GEN_4136 : ~(_GEN_1271 & _GEN_350) & _GEN_4136) : _GEN_4136;
  wire        _GEN_4170 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_351 & _GEN_4137 : ~(_GEN_1271 & _GEN_351) & _GEN_4137) : _GEN_4137;
  wire        _GEN_4171 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_352 & _GEN_4138 : ~(_GEN_1271 & _GEN_352) & _GEN_4138) : _GEN_4138;
  wire        _GEN_4172 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_353 & _GEN_4139 : ~(_GEN_1271 & _GEN_353) & _GEN_4139) : _GEN_4139;
  wire        _GEN_4173 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_354 & _GEN_4140 : ~(_GEN_1271 & _GEN_354) & _GEN_4140) : _GEN_4140;
  wire        _GEN_4174 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_355 & _GEN_4141 : ~(_GEN_1271 & _GEN_355) & _GEN_4141) : _GEN_4141;
  wire        _GEN_4175 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_356 & _GEN_4142 : ~(_GEN_1271 & _GEN_356) & _GEN_4142) : _GEN_4142;
  wire        _GEN_4176 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_357 & _GEN_4143 : ~(_GEN_1271 & _GEN_357) & _GEN_4143) : _GEN_4143;
  wire        _GEN_4177 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_358 & _GEN_4144 : ~(_GEN_1271 & _GEN_358) & _GEN_4144) : _GEN_4144;
  wire        _GEN_4178 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_359 & _GEN_4145 : ~(_GEN_1271 & _GEN_359) & _GEN_4145) : _GEN_4145;
  wire        _GEN_4179 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_360 & _GEN_4146 : ~(_GEN_1271 & _GEN_360) & _GEN_4146) : _GEN_4146;
  wire        _GEN_4180 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_361 & _GEN_4147 : ~(_GEN_1271 & _GEN_361) & _GEN_4147) : _GEN_4147;
  wire        _GEN_4181 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_362 & _GEN_4148 : ~(_GEN_1271 & _GEN_362) & _GEN_4148) : _GEN_4148;
  wire        _GEN_4182 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_363 & _GEN_4149 : ~(_GEN_1271 & _GEN_363) & _GEN_4149) : _GEN_4149;
  wire        _GEN_4183 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_364 & _GEN_4150 : ~(_GEN_1271 & _GEN_364) & _GEN_4150) : _GEN_4150;
  wire        _GEN_4184 = _GEN_1273 ? (_GEN_4153 ? ~_GEN_365 & _GEN_4151 : ~(_GEN_1271 & _GEN_365) & _GEN_4151) : _GEN_4151;
  wire        _GEN_4185 = _GEN_1273 ? (_GEN_4153 ? ~(&lcam_ldq_idx_1) & _GEN_4152 : ~(_GEN_1271 & (&lcam_ldq_idx_1)) & _GEN_4152) : _GEN_4152;
  wire        _GEN_4186 = _GEN_1280 | _GEN_1281;
  wire        _GEN_4187 = _GEN_1278 ? (_GEN_4186 ? (|lcam_ldq_idx_0) & _GEN_4154 : ~(_GEN_1282 & ~(|lcam_ldq_idx_0)) & _GEN_4154) : _GEN_4154;
  wire        _GEN_4188 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_296 & _GEN_4155 : ~(_GEN_1282 & _GEN_296) & _GEN_4155) : _GEN_4155;
  wire        _GEN_4189 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_297 & _GEN_4156 : ~(_GEN_1282 & _GEN_297) & _GEN_4156) : _GEN_4156;
  wire        _GEN_4190 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_298 & _GEN_4157 : ~(_GEN_1282 & _GEN_298) & _GEN_4157) : _GEN_4157;
  wire        _GEN_4191 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_299 & _GEN_4158 : ~(_GEN_1282 & _GEN_299) & _GEN_4158) : _GEN_4158;
  wire        _GEN_4192 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_300 & _GEN_4159 : ~(_GEN_1282 & _GEN_300) & _GEN_4159) : _GEN_4159;
  wire        _GEN_4193 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_301 & _GEN_4160 : ~(_GEN_1282 & _GEN_301) & _GEN_4160) : _GEN_4160;
  wire        _GEN_4194 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_302 & _GEN_4161 : ~(_GEN_1282 & _GEN_302) & _GEN_4161) : _GEN_4161;
  wire        _GEN_4195 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_303 & _GEN_4162 : ~(_GEN_1282 & _GEN_303) & _GEN_4162) : _GEN_4162;
  wire        _GEN_4196 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_304 & _GEN_4163 : ~(_GEN_1282 & _GEN_304) & _GEN_4163) : _GEN_4163;
  wire        _GEN_4197 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_305 & _GEN_4164 : ~(_GEN_1282 & _GEN_305) & _GEN_4164) : _GEN_4164;
  wire        _GEN_4198 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_306 & _GEN_4165 : ~(_GEN_1282 & _GEN_306) & _GEN_4165) : _GEN_4165;
  wire        _GEN_4199 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_307 & _GEN_4166 : ~(_GEN_1282 & _GEN_307) & _GEN_4166) : _GEN_4166;
  wire        _GEN_4200 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_308 & _GEN_4167 : ~(_GEN_1282 & _GEN_308) & _GEN_4167) : _GEN_4167;
  wire        _GEN_4201 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_309 & _GEN_4168 : ~(_GEN_1282 & _GEN_309) & _GEN_4168) : _GEN_4168;
  wire        _GEN_4202 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_310 & _GEN_4169 : ~(_GEN_1282 & _GEN_310) & _GEN_4169) : _GEN_4169;
  wire        _GEN_4203 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_311 & _GEN_4170 : ~(_GEN_1282 & _GEN_311) & _GEN_4170) : _GEN_4170;
  wire        _GEN_4204 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_312 & _GEN_4171 : ~(_GEN_1282 & _GEN_312) & _GEN_4171) : _GEN_4171;
  wire        _GEN_4205 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_313 & _GEN_4172 : ~(_GEN_1282 & _GEN_313) & _GEN_4172) : _GEN_4172;
  wire        _GEN_4206 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_314 & _GEN_4173 : ~(_GEN_1282 & _GEN_314) & _GEN_4173) : _GEN_4173;
  wire        _GEN_4207 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_315 & _GEN_4174 : ~(_GEN_1282 & _GEN_315) & _GEN_4174) : _GEN_4174;
  wire        _GEN_4208 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_316 & _GEN_4175 : ~(_GEN_1282 & _GEN_316) & _GEN_4175) : _GEN_4175;
  wire        _GEN_4209 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_317 & _GEN_4176 : ~(_GEN_1282 & _GEN_317) & _GEN_4176) : _GEN_4176;
  wire        _GEN_4210 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_318 & _GEN_4177 : ~(_GEN_1282 & _GEN_318) & _GEN_4177) : _GEN_4177;
  wire        _GEN_4211 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_319 & _GEN_4178 : ~(_GEN_1282 & _GEN_319) & _GEN_4178) : _GEN_4178;
  wire        _GEN_4212 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_320 & _GEN_4179 : ~(_GEN_1282 & _GEN_320) & _GEN_4179) : _GEN_4179;
  wire        _GEN_4213 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_321 & _GEN_4180 : ~(_GEN_1282 & _GEN_321) & _GEN_4180) : _GEN_4180;
  wire        _GEN_4214 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_322 & _GEN_4181 : ~(_GEN_1282 & _GEN_322) & _GEN_4181) : _GEN_4181;
  wire        _GEN_4215 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_323 & _GEN_4182 : ~(_GEN_1282 & _GEN_323) & _GEN_4182) : _GEN_4182;
  wire        _GEN_4216 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_324 & _GEN_4183 : ~(_GEN_1282 & _GEN_324) & _GEN_4183) : _GEN_4183;
  wire        _GEN_4217 = _GEN_1278 ? (_GEN_4186 ? ~_GEN_325 & _GEN_4184 : ~(_GEN_1282 & _GEN_325) & _GEN_4184) : _GEN_4184;
  wire        _GEN_4218 = _GEN_1278 ? (_GEN_4186 ? ~(&lcam_ldq_idx_0) & _GEN_4185 : ~(_GEN_1282 & (&lcam_ldq_idx_0)) & _GEN_4185) : _GEN_4185;
  wire        _GEN_4219 = _GEN_1286 | _GEN_1287;
  wire        _GEN_4220 = _GEN_1284 ? (_GEN_4219 ? (|lcam_ldq_idx_1) & _GEN_4187 : ~(_GEN_1282 & ~(|lcam_ldq_idx_1)) & _GEN_4187) : _GEN_4187;
  wire        _GEN_4221 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_336 & _GEN_4188 : ~(_GEN_1282 & _GEN_336) & _GEN_4188) : _GEN_4188;
  wire        _GEN_4222 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_337 & _GEN_4189 : ~(_GEN_1282 & _GEN_337) & _GEN_4189) : _GEN_4189;
  wire        _GEN_4223 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_338 & _GEN_4190 : ~(_GEN_1282 & _GEN_338) & _GEN_4190) : _GEN_4190;
  wire        _GEN_4224 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_339 & _GEN_4191 : ~(_GEN_1282 & _GEN_339) & _GEN_4191) : _GEN_4191;
  wire        _GEN_4225 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_340 & _GEN_4192 : ~(_GEN_1282 & _GEN_340) & _GEN_4192) : _GEN_4192;
  wire        _GEN_4226 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_341 & _GEN_4193 : ~(_GEN_1282 & _GEN_341) & _GEN_4193) : _GEN_4193;
  wire        _GEN_4227 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_342 & _GEN_4194 : ~(_GEN_1282 & _GEN_342) & _GEN_4194) : _GEN_4194;
  wire        _GEN_4228 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_343 & _GEN_4195 : ~(_GEN_1282 & _GEN_343) & _GEN_4195) : _GEN_4195;
  wire        _GEN_4229 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_344 & _GEN_4196 : ~(_GEN_1282 & _GEN_344) & _GEN_4196) : _GEN_4196;
  wire        _GEN_4230 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_345 & _GEN_4197 : ~(_GEN_1282 & _GEN_345) & _GEN_4197) : _GEN_4197;
  wire        _GEN_4231 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_346 & _GEN_4198 : ~(_GEN_1282 & _GEN_346) & _GEN_4198) : _GEN_4198;
  wire        _GEN_4232 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_347 & _GEN_4199 : ~(_GEN_1282 & _GEN_347) & _GEN_4199) : _GEN_4199;
  wire        _GEN_4233 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_348 & _GEN_4200 : ~(_GEN_1282 & _GEN_348) & _GEN_4200) : _GEN_4200;
  wire        _GEN_4234 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_349 & _GEN_4201 : ~(_GEN_1282 & _GEN_349) & _GEN_4201) : _GEN_4201;
  wire        _GEN_4235 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_350 & _GEN_4202 : ~(_GEN_1282 & _GEN_350) & _GEN_4202) : _GEN_4202;
  wire        _GEN_4236 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_351 & _GEN_4203 : ~(_GEN_1282 & _GEN_351) & _GEN_4203) : _GEN_4203;
  wire        _GEN_4237 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_352 & _GEN_4204 : ~(_GEN_1282 & _GEN_352) & _GEN_4204) : _GEN_4204;
  wire        _GEN_4238 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_353 & _GEN_4205 : ~(_GEN_1282 & _GEN_353) & _GEN_4205) : _GEN_4205;
  wire        _GEN_4239 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_354 & _GEN_4206 : ~(_GEN_1282 & _GEN_354) & _GEN_4206) : _GEN_4206;
  wire        _GEN_4240 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_355 & _GEN_4207 : ~(_GEN_1282 & _GEN_355) & _GEN_4207) : _GEN_4207;
  wire        _GEN_4241 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_356 & _GEN_4208 : ~(_GEN_1282 & _GEN_356) & _GEN_4208) : _GEN_4208;
  wire        _GEN_4242 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_357 & _GEN_4209 : ~(_GEN_1282 & _GEN_357) & _GEN_4209) : _GEN_4209;
  wire        _GEN_4243 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_358 & _GEN_4210 : ~(_GEN_1282 & _GEN_358) & _GEN_4210) : _GEN_4210;
  wire        _GEN_4244 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_359 & _GEN_4211 : ~(_GEN_1282 & _GEN_359) & _GEN_4211) : _GEN_4211;
  wire        _GEN_4245 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_360 & _GEN_4212 : ~(_GEN_1282 & _GEN_360) & _GEN_4212) : _GEN_4212;
  wire        _GEN_4246 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_361 & _GEN_4213 : ~(_GEN_1282 & _GEN_361) & _GEN_4213) : _GEN_4213;
  wire        _GEN_4247 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_362 & _GEN_4214 : ~(_GEN_1282 & _GEN_362) & _GEN_4214) : _GEN_4214;
  wire        _GEN_4248 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_363 & _GEN_4215 : ~(_GEN_1282 & _GEN_363) & _GEN_4215) : _GEN_4215;
  wire        _GEN_4249 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_364 & _GEN_4216 : ~(_GEN_1282 & _GEN_364) & _GEN_4216) : _GEN_4216;
  wire        _GEN_4250 = _GEN_1284 ? (_GEN_4219 ? ~_GEN_365 & _GEN_4217 : ~(_GEN_1282 & _GEN_365) & _GEN_4217) : _GEN_4217;
  wire        _GEN_4251 = _GEN_1284 ? (_GEN_4219 ? ~(&lcam_ldq_idx_1) & _GEN_4218 : ~(_GEN_1282 & (&lcam_ldq_idx_1)) & _GEN_4218) : _GEN_4218;
  wire        _GEN_4252 = _GEN_1291 | _GEN_1292;
  wire        _GEN_4253 = _GEN_1289 ? (_GEN_4252 ? (|lcam_ldq_idx_0) & _GEN_4220 : ~(_GEN_1293 & ~(|lcam_ldq_idx_0)) & _GEN_4220) : _GEN_4220;
  wire        _GEN_4254 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_296 & _GEN_4221 : ~(_GEN_1293 & _GEN_296) & _GEN_4221) : _GEN_4221;
  wire        _GEN_4255 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_297 & _GEN_4222 : ~(_GEN_1293 & _GEN_297) & _GEN_4222) : _GEN_4222;
  wire        _GEN_4256 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_298 & _GEN_4223 : ~(_GEN_1293 & _GEN_298) & _GEN_4223) : _GEN_4223;
  wire        _GEN_4257 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_299 & _GEN_4224 : ~(_GEN_1293 & _GEN_299) & _GEN_4224) : _GEN_4224;
  wire        _GEN_4258 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_300 & _GEN_4225 : ~(_GEN_1293 & _GEN_300) & _GEN_4225) : _GEN_4225;
  wire        _GEN_4259 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_301 & _GEN_4226 : ~(_GEN_1293 & _GEN_301) & _GEN_4226) : _GEN_4226;
  wire        _GEN_4260 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_302 & _GEN_4227 : ~(_GEN_1293 & _GEN_302) & _GEN_4227) : _GEN_4227;
  wire        _GEN_4261 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_303 & _GEN_4228 : ~(_GEN_1293 & _GEN_303) & _GEN_4228) : _GEN_4228;
  wire        _GEN_4262 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_304 & _GEN_4229 : ~(_GEN_1293 & _GEN_304) & _GEN_4229) : _GEN_4229;
  wire        _GEN_4263 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_305 & _GEN_4230 : ~(_GEN_1293 & _GEN_305) & _GEN_4230) : _GEN_4230;
  wire        _GEN_4264 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_306 & _GEN_4231 : ~(_GEN_1293 & _GEN_306) & _GEN_4231) : _GEN_4231;
  wire        _GEN_4265 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_307 & _GEN_4232 : ~(_GEN_1293 & _GEN_307) & _GEN_4232) : _GEN_4232;
  wire        _GEN_4266 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_308 & _GEN_4233 : ~(_GEN_1293 & _GEN_308) & _GEN_4233) : _GEN_4233;
  wire        _GEN_4267 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_309 & _GEN_4234 : ~(_GEN_1293 & _GEN_309) & _GEN_4234) : _GEN_4234;
  wire        _GEN_4268 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_310 & _GEN_4235 : ~(_GEN_1293 & _GEN_310) & _GEN_4235) : _GEN_4235;
  wire        _GEN_4269 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_311 & _GEN_4236 : ~(_GEN_1293 & _GEN_311) & _GEN_4236) : _GEN_4236;
  wire        _GEN_4270 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_312 & _GEN_4237 : ~(_GEN_1293 & _GEN_312) & _GEN_4237) : _GEN_4237;
  wire        _GEN_4271 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_313 & _GEN_4238 : ~(_GEN_1293 & _GEN_313) & _GEN_4238) : _GEN_4238;
  wire        _GEN_4272 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_314 & _GEN_4239 : ~(_GEN_1293 & _GEN_314) & _GEN_4239) : _GEN_4239;
  wire        _GEN_4273 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_315 & _GEN_4240 : ~(_GEN_1293 & _GEN_315) & _GEN_4240) : _GEN_4240;
  wire        _GEN_4274 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_316 & _GEN_4241 : ~(_GEN_1293 & _GEN_316) & _GEN_4241) : _GEN_4241;
  wire        _GEN_4275 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_317 & _GEN_4242 : ~(_GEN_1293 & _GEN_317) & _GEN_4242) : _GEN_4242;
  wire        _GEN_4276 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_318 & _GEN_4243 : ~(_GEN_1293 & _GEN_318) & _GEN_4243) : _GEN_4243;
  wire        _GEN_4277 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_319 & _GEN_4244 : ~(_GEN_1293 & _GEN_319) & _GEN_4244) : _GEN_4244;
  wire        _GEN_4278 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_320 & _GEN_4245 : ~(_GEN_1293 & _GEN_320) & _GEN_4245) : _GEN_4245;
  wire        _GEN_4279 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_321 & _GEN_4246 : ~(_GEN_1293 & _GEN_321) & _GEN_4246) : _GEN_4246;
  wire        _GEN_4280 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_322 & _GEN_4247 : ~(_GEN_1293 & _GEN_322) & _GEN_4247) : _GEN_4247;
  wire        _GEN_4281 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_323 & _GEN_4248 : ~(_GEN_1293 & _GEN_323) & _GEN_4248) : _GEN_4248;
  wire        _GEN_4282 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_324 & _GEN_4249 : ~(_GEN_1293 & _GEN_324) & _GEN_4249) : _GEN_4249;
  wire        _GEN_4283 = _GEN_1289 ? (_GEN_4252 ? ~_GEN_325 & _GEN_4250 : ~(_GEN_1293 & _GEN_325) & _GEN_4250) : _GEN_4250;
  wire        _GEN_4284 = _GEN_1289 ? (_GEN_4252 ? ~(&lcam_ldq_idx_0) & _GEN_4251 : ~(_GEN_1293 & (&lcam_ldq_idx_0)) & _GEN_4251) : _GEN_4251;
  wire        _GEN_4285 = _GEN_1297 | _GEN_1298;
  wire        _GEN_4286 = _GEN_1295 ? (_GEN_4285 ? (|lcam_ldq_idx_1) & _GEN_4253 : ~(_GEN_1293 & ~(|lcam_ldq_idx_1)) & _GEN_4253) : _GEN_4253;
  wire        _GEN_4287 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_336 & _GEN_4254 : ~(_GEN_1293 & _GEN_336) & _GEN_4254) : _GEN_4254;
  wire        _GEN_4288 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_337 & _GEN_4255 : ~(_GEN_1293 & _GEN_337) & _GEN_4255) : _GEN_4255;
  wire        _GEN_4289 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_338 & _GEN_4256 : ~(_GEN_1293 & _GEN_338) & _GEN_4256) : _GEN_4256;
  wire        _GEN_4290 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_339 & _GEN_4257 : ~(_GEN_1293 & _GEN_339) & _GEN_4257) : _GEN_4257;
  wire        _GEN_4291 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_340 & _GEN_4258 : ~(_GEN_1293 & _GEN_340) & _GEN_4258) : _GEN_4258;
  wire        _GEN_4292 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_341 & _GEN_4259 : ~(_GEN_1293 & _GEN_341) & _GEN_4259) : _GEN_4259;
  wire        _GEN_4293 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_342 & _GEN_4260 : ~(_GEN_1293 & _GEN_342) & _GEN_4260) : _GEN_4260;
  wire        _GEN_4294 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_343 & _GEN_4261 : ~(_GEN_1293 & _GEN_343) & _GEN_4261) : _GEN_4261;
  wire        _GEN_4295 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_344 & _GEN_4262 : ~(_GEN_1293 & _GEN_344) & _GEN_4262) : _GEN_4262;
  wire        _GEN_4296 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_345 & _GEN_4263 : ~(_GEN_1293 & _GEN_345) & _GEN_4263) : _GEN_4263;
  wire        _GEN_4297 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_346 & _GEN_4264 : ~(_GEN_1293 & _GEN_346) & _GEN_4264) : _GEN_4264;
  wire        _GEN_4298 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_347 & _GEN_4265 : ~(_GEN_1293 & _GEN_347) & _GEN_4265) : _GEN_4265;
  wire        _GEN_4299 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_348 & _GEN_4266 : ~(_GEN_1293 & _GEN_348) & _GEN_4266) : _GEN_4266;
  wire        _GEN_4300 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_349 & _GEN_4267 : ~(_GEN_1293 & _GEN_349) & _GEN_4267) : _GEN_4267;
  wire        _GEN_4301 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_350 & _GEN_4268 : ~(_GEN_1293 & _GEN_350) & _GEN_4268) : _GEN_4268;
  wire        _GEN_4302 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_351 & _GEN_4269 : ~(_GEN_1293 & _GEN_351) & _GEN_4269) : _GEN_4269;
  wire        _GEN_4303 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_352 & _GEN_4270 : ~(_GEN_1293 & _GEN_352) & _GEN_4270) : _GEN_4270;
  wire        _GEN_4304 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_353 & _GEN_4271 : ~(_GEN_1293 & _GEN_353) & _GEN_4271) : _GEN_4271;
  wire        _GEN_4305 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_354 & _GEN_4272 : ~(_GEN_1293 & _GEN_354) & _GEN_4272) : _GEN_4272;
  wire        _GEN_4306 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_355 & _GEN_4273 : ~(_GEN_1293 & _GEN_355) & _GEN_4273) : _GEN_4273;
  wire        _GEN_4307 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_356 & _GEN_4274 : ~(_GEN_1293 & _GEN_356) & _GEN_4274) : _GEN_4274;
  wire        _GEN_4308 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_357 & _GEN_4275 : ~(_GEN_1293 & _GEN_357) & _GEN_4275) : _GEN_4275;
  wire        _GEN_4309 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_358 & _GEN_4276 : ~(_GEN_1293 & _GEN_358) & _GEN_4276) : _GEN_4276;
  wire        _GEN_4310 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_359 & _GEN_4277 : ~(_GEN_1293 & _GEN_359) & _GEN_4277) : _GEN_4277;
  wire        _GEN_4311 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_360 & _GEN_4278 : ~(_GEN_1293 & _GEN_360) & _GEN_4278) : _GEN_4278;
  wire        _GEN_4312 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_361 & _GEN_4279 : ~(_GEN_1293 & _GEN_361) & _GEN_4279) : _GEN_4279;
  wire        _GEN_4313 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_362 & _GEN_4280 : ~(_GEN_1293 & _GEN_362) & _GEN_4280) : _GEN_4280;
  wire        _GEN_4314 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_363 & _GEN_4281 : ~(_GEN_1293 & _GEN_363) & _GEN_4281) : _GEN_4281;
  wire        _GEN_4315 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_364 & _GEN_4282 : ~(_GEN_1293 & _GEN_364) & _GEN_4282) : _GEN_4282;
  wire        _GEN_4316 = _GEN_1295 ? (_GEN_4285 ? ~_GEN_365 & _GEN_4283 : ~(_GEN_1293 & _GEN_365) & _GEN_4283) : _GEN_4283;
  wire        _GEN_4317 = _GEN_1295 ? (_GEN_4285 ? ~(&lcam_ldq_idx_1) & _GEN_4284 : ~(_GEN_1293 & (&lcam_ldq_idx_1)) & _GEN_4284) : _GEN_4284;
  wire        _GEN_4318 = _GEN_1302 | _GEN_1303;
  wire        _GEN_4319 = _GEN_1300 ? (_GEN_4318 ? (|lcam_ldq_idx_0) & _GEN_4286 : ~(_GEN_1304 & ~(|lcam_ldq_idx_0)) & _GEN_4286) : _GEN_4286;
  wire        _GEN_4320 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_296 & _GEN_4287 : ~(_GEN_1304 & _GEN_296) & _GEN_4287) : _GEN_4287;
  wire        _GEN_4321 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_297 & _GEN_4288 : ~(_GEN_1304 & _GEN_297) & _GEN_4288) : _GEN_4288;
  wire        _GEN_4322 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_298 & _GEN_4289 : ~(_GEN_1304 & _GEN_298) & _GEN_4289) : _GEN_4289;
  wire        _GEN_4323 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_299 & _GEN_4290 : ~(_GEN_1304 & _GEN_299) & _GEN_4290) : _GEN_4290;
  wire        _GEN_4324 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_300 & _GEN_4291 : ~(_GEN_1304 & _GEN_300) & _GEN_4291) : _GEN_4291;
  wire        _GEN_4325 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_301 & _GEN_4292 : ~(_GEN_1304 & _GEN_301) & _GEN_4292) : _GEN_4292;
  wire        _GEN_4326 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_302 & _GEN_4293 : ~(_GEN_1304 & _GEN_302) & _GEN_4293) : _GEN_4293;
  wire        _GEN_4327 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_303 & _GEN_4294 : ~(_GEN_1304 & _GEN_303) & _GEN_4294) : _GEN_4294;
  wire        _GEN_4328 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_304 & _GEN_4295 : ~(_GEN_1304 & _GEN_304) & _GEN_4295) : _GEN_4295;
  wire        _GEN_4329 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_305 & _GEN_4296 : ~(_GEN_1304 & _GEN_305) & _GEN_4296) : _GEN_4296;
  wire        _GEN_4330 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_306 & _GEN_4297 : ~(_GEN_1304 & _GEN_306) & _GEN_4297) : _GEN_4297;
  wire        _GEN_4331 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_307 & _GEN_4298 : ~(_GEN_1304 & _GEN_307) & _GEN_4298) : _GEN_4298;
  wire        _GEN_4332 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_308 & _GEN_4299 : ~(_GEN_1304 & _GEN_308) & _GEN_4299) : _GEN_4299;
  wire        _GEN_4333 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_309 & _GEN_4300 : ~(_GEN_1304 & _GEN_309) & _GEN_4300) : _GEN_4300;
  wire        _GEN_4334 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_310 & _GEN_4301 : ~(_GEN_1304 & _GEN_310) & _GEN_4301) : _GEN_4301;
  wire        _GEN_4335 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_311 & _GEN_4302 : ~(_GEN_1304 & _GEN_311) & _GEN_4302) : _GEN_4302;
  wire        _GEN_4336 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_312 & _GEN_4303 : ~(_GEN_1304 & _GEN_312) & _GEN_4303) : _GEN_4303;
  wire        _GEN_4337 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_313 & _GEN_4304 : ~(_GEN_1304 & _GEN_313) & _GEN_4304) : _GEN_4304;
  wire        _GEN_4338 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_314 & _GEN_4305 : ~(_GEN_1304 & _GEN_314) & _GEN_4305) : _GEN_4305;
  wire        _GEN_4339 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_315 & _GEN_4306 : ~(_GEN_1304 & _GEN_315) & _GEN_4306) : _GEN_4306;
  wire        _GEN_4340 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_316 & _GEN_4307 : ~(_GEN_1304 & _GEN_316) & _GEN_4307) : _GEN_4307;
  wire        _GEN_4341 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_317 & _GEN_4308 : ~(_GEN_1304 & _GEN_317) & _GEN_4308) : _GEN_4308;
  wire        _GEN_4342 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_318 & _GEN_4309 : ~(_GEN_1304 & _GEN_318) & _GEN_4309) : _GEN_4309;
  wire        _GEN_4343 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_319 & _GEN_4310 : ~(_GEN_1304 & _GEN_319) & _GEN_4310) : _GEN_4310;
  wire        _GEN_4344 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_320 & _GEN_4311 : ~(_GEN_1304 & _GEN_320) & _GEN_4311) : _GEN_4311;
  wire        _GEN_4345 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_321 & _GEN_4312 : ~(_GEN_1304 & _GEN_321) & _GEN_4312) : _GEN_4312;
  wire        _GEN_4346 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_322 & _GEN_4313 : ~(_GEN_1304 & _GEN_322) & _GEN_4313) : _GEN_4313;
  wire        _GEN_4347 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_323 & _GEN_4314 : ~(_GEN_1304 & _GEN_323) & _GEN_4314) : _GEN_4314;
  wire        _GEN_4348 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_324 & _GEN_4315 : ~(_GEN_1304 & _GEN_324) & _GEN_4315) : _GEN_4315;
  wire        _GEN_4349 = _GEN_1300 ? (_GEN_4318 ? ~_GEN_325 & _GEN_4316 : ~(_GEN_1304 & _GEN_325) & _GEN_4316) : _GEN_4316;
  wire        _GEN_4350 = _GEN_1300 ? (_GEN_4318 ? ~(&lcam_ldq_idx_0) & _GEN_4317 : ~(_GEN_1304 & (&lcam_ldq_idx_0)) & _GEN_4317) : _GEN_4317;
  wire        _GEN_4351 = _GEN_1308 | _GEN_1309;
  wire        _GEN_4352 = _GEN_1306 ? (_GEN_4351 ? (|lcam_ldq_idx_1) & _GEN_4319 : ~(_GEN_1304 & ~(|lcam_ldq_idx_1)) & _GEN_4319) : _GEN_4319;
  wire        _GEN_4353 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_336 & _GEN_4320 : ~(_GEN_1304 & _GEN_336) & _GEN_4320) : _GEN_4320;
  wire        _GEN_4354 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_337 & _GEN_4321 : ~(_GEN_1304 & _GEN_337) & _GEN_4321) : _GEN_4321;
  wire        _GEN_4355 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_338 & _GEN_4322 : ~(_GEN_1304 & _GEN_338) & _GEN_4322) : _GEN_4322;
  wire        _GEN_4356 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_339 & _GEN_4323 : ~(_GEN_1304 & _GEN_339) & _GEN_4323) : _GEN_4323;
  wire        _GEN_4357 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_340 & _GEN_4324 : ~(_GEN_1304 & _GEN_340) & _GEN_4324) : _GEN_4324;
  wire        _GEN_4358 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_341 & _GEN_4325 : ~(_GEN_1304 & _GEN_341) & _GEN_4325) : _GEN_4325;
  wire        _GEN_4359 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_342 & _GEN_4326 : ~(_GEN_1304 & _GEN_342) & _GEN_4326) : _GEN_4326;
  wire        _GEN_4360 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_343 & _GEN_4327 : ~(_GEN_1304 & _GEN_343) & _GEN_4327) : _GEN_4327;
  wire        _GEN_4361 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_344 & _GEN_4328 : ~(_GEN_1304 & _GEN_344) & _GEN_4328) : _GEN_4328;
  wire        _GEN_4362 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_345 & _GEN_4329 : ~(_GEN_1304 & _GEN_345) & _GEN_4329) : _GEN_4329;
  wire        _GEN_4363 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_346 & _GEN_4330 : ~(_GEN_1304 & _GEN_346) & _GEN_4330) : _GEN_4330;
  wire        _GEN_4364 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_347 & _GEN_4331 : ~(_GEN_1304 & _GEN_347) & _GEN_4331) : _GEN_4331;
  wire        _GEN_4365 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_348 & _GEN_4332 : ~(_GEN_1304 & _GEN_348) & _GEN_4332) : _GEN_4332;
  wire        _GEN_4366 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_349 & _GEN_4333 : ~(_GEN_1304 & _GEN_349) & _GEN_4333) : _GEN_4333;
  wire        _GEN_4367 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_350 & _GEN_4334 : ~(_GEN_1304 & _GEN_350) & _GEN_4334) : _GEN_4334;
  wire        _GEN_4368 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_351 & _GEN_4335 : ~(_GEN_1304 & _GEN_351) & _GEN_4335) : _GEN_4335;
  wire        _GEN_4369 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_352 & _GEN_4336 : ~(_GEN_1304 & _GEN_352) & _GEN_4336) : _GEN_4336;
  wire        _GEN_4370 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_353 & _GEN_4337 : ~(_GEN_1304 & _GEN_353) & _GEN_4337) : _GEN_4337;
  wire        _GEN_4371 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_354 & _GEN_4338 : ~(_GEN_1304 & _GEN_354) & _GEN_4338) : _GEN_4338;
  wire        _GEN_4372 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_355 & _GEN_4339 : ~(_GEN_1304 & _GEN_355) & _GEN_4339) : _GEN_4339;
  wire        _GEN_4373 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_356 & _GEN_4340 : ~(_GEN_1304 & _GEN_356) & _GEN_4340) : _GEN_4340;
  wire        _GEN_4374 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_357 & _GEN_4341 : ~(_GEN_1304 & _GEN_357) & _GEN_4341) : _GEN_4341;
  wire        _GEN_4375 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_358 & _GEN_4342 : ~(_GEN_1304 & _GEN_358) & _GEN_4342) : _GEN_4342;
  wire        _GEN_4376 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_359 & _GEN_4343 : ~(_GEN_1304 & _GEN_359) & _GEN_4343) : _GEN_4343;
  wire        _GEN_4377 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_360 & _GEN_4344 : ~(_GEN_1304 & _GEN_360) & _GEN_4344) : _GEN_4344;
  wire        _GEN_4378 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_361 & _GEN_4345 : ~(_GEN_1304 & _GEN_361) & _GEN_4345) : _GEN_4345;
  wire        _GEN_4379 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_362 & _GEN_4346 : ~(_GEN_1304 & _GEN_362) & _GEN_4346) : _GEN_4346;
  wire        _GEN_4380 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_363 & _GEN_4347 : ~(_GEN_1304 & _GEN_363) & _GEN_4347) : _GEN_4347;
  wire        _GEN_4381 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_364 & _GEN_4348 : ~(_GEN_1304 & _GEN_364) & _GEN_4348) : _GEN_4348;
  wire        _GEN_4382 = _GEN_1306 ? (_GEN_4351 ? ~_GEN_365 & _GEN_4349 : ~(_GEN_1304 & _GEN_365) & _GEN_4349) : _GEN_4349;
  wire        _GEN_4383 = _GEN_1306 ? (_GEN_4351 ? ~(&lcam_ldq_idx_1) & _GEN_4350 : ~(_GEN_1304 & (&lcam_ldq_idx_1)) & _GEN_4350) : _GEN_4350;
  wire        _GEN_4384 = _GEN_1313 | _GEN_1314;
  wire        _GEN_4385 = _GEN_1311 ? (_GEN_4384 ? (|lcam_ldq_idx_0) & _GEN_4352 : ~(_GEN_1315 & ~(|lcam_ldq_idx_0)) & _GEN_4352) : _GEN_4352;
  wire        _GEN_4386 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_296 & _GEN_4353 : ~(_GEN_1315 & _GEN_296) & _GEN_4353) : _GEN_4353;
  wire        _GEN_4387 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_297 & _GEN_4354 : ~(_GEN_1315 & _GEN_297) & _GEN_4354) : _GEN_4354;
  wire        _GEN_4388 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_298 & _GEN_4355 : ~(_GEN_1315 & _GEN_298) & _GEN_4355) : _GEN_4355;
  wire        _GEN_4389 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_299 & _GEN_4356 : ~(_GEN_1315 & _GEN_299) & _GEN_4356) : _GEN_4356;
  wire        _GEN_4390 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_300 & _GEN_4357 : ~(_GEN_1315 & _GEN_300) & _GEN_4357) : _GEN_4357;
  wire        _GEN_4391 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_301 & _GEN_4358 : ~(_GEN_1315 & _GEN_301) & _GEN_4358) : _GEN_4358;
  wire        _GEN_4392 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_302 & _GEN_4359 : ~(_GEN_1315 & _GEN_302) & _GEN_4359) : _GEN_4359;
  wire        _GEN_4393 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_303 & _GEN_4360 : ~(_GEN_1315 & _GEN_303) & _GEN_4360) : _GEN_4360;
  wire        _GEN_4394 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_304 & _GEN_4361 : ~(_GEN_1315 & _GEN_304) & _GEN_4361) : _GEN_4361;
  wire        _GEN_4395 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_305 & _GEN_4362 : ~(_GEN_1315 & _GEN_305) & _GEN_4362) : _GEN_4362;
  wire        _GEN_4396 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_306 & _GEN_4363 : ~(_GEN_1315 & _GEN_306) & _GEN_4363) : _GEN_4363;
  wire        _GEN_4397 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_307 & _GEN_4364 : ~(_GEN_1315 & _GEN_307) & _GEN_4364) : _GEN_4364;
  wire        _GEN_4398 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_308 & _GEN_4365 : ~(_GEN_1315 & _GEN_308) & _GEN_4365) : _GEN_4365;
  wire        _GEN_4399 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_309 & _GEN_4366 : ~(_GEN_1315 & _GEN_309) & _GEN_4366) : _GEN_4366;
  wire        _GEN_4400 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_310 & _GEN_4367 : ~(_GEN_1315 & _GEN_310) & _GEN_4367) : _GEN_4367;
  wire        _GEN_4401 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_311 & _GEN_4368 : ~(_GEN_1315 & _GEN_311) & _GEN_4368) : _GEN_4368;
  wire        _GEN_4402 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_312 & _GEN_4369 : ~(_GEN_1315 & _GEN_312) & _GEN_4369) : _GEN_4369;
  wire        _GEN_4403 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_313 & _GEN_4370 : ~(_GEN_1315 & _GEN_313) & _GEN_4370) : _GEN_4370;
  wire        _GEN_4404 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_314 & _GEN_4371 : ~(_GEN_1315 & _GEN_314) & _GEN_4371) : _GEN_4371;
  wire        _GEN_4405 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_315 & _GEN_4372 : ~(_GEN_1315 & _GEN_315) & _GEN_4372) : _GEN_4372;
  wire        _GEN_4406 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_316 & _GEN_4373 : ~(_GEN_1315 & _GEN_316) & _GEN_4373) : _GEN_4373;
  wire        _GEN_4407 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_317 & _GEN_4374 : ~(_GEN_1315 & _GEN_317) & _GEN_4374) : _GEN_4374;
  wire        _GEN_4408 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_318 & _GEN_4375 : ~(_GEN_1315 & _GEN_318) & _GEN_4375) : _GEN_4375;
  wire        _GEN_4409 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_319 & _GEN_4376 : ~(_GEN_1315 & _GEN_319) & _GEN_4376) : _GEN_4376;
  wire        _GEN_4410 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_320 & _GEN_4377 : ~(_GEN_1315 & _GEN_320) & _GEN_4377) : _GEN_4377;
  wire        _GEN_4411 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_321 & _GEN_4378 : ~(_GEN_1315 & _GEN_321) & _GEN_4378) : _GEN_4378;
  wire        _GEN_4412 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_322 & _GEN_4379 : ~(_GEN_1315 & _GEN_322) & _GEN_4379) : _GEN_4379;
  wire        _GEN_4413 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_323 & _GEN_4380 : ~(_GEN_1315 & _GEN_323) & _GEN_4380) : _GEN_4380;
  wire        _GEN_4414 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_324 & _GEN_4381 : ~(_GEN_1315 & _GEN_324) & _GEN_4381) : _GEN_4381;
  wire        _GEN_4415 = _GEN_1311 ? (_GEN_4384 ? ~_GEN_325 & _GEN_4382 : ~(_GEN_1315 & _GEN_325) & _GEN_4382) : _GEN_4382;
  wire        _GEN_4416 = _GEN_1311 ? (_GEN_4384 ? ~(&lcam_ldq_idx_0) & _GEN_4383 : ~(_GEN_1315 & (&lcam_ldq_idx_0)) & _GEN_4383) : _GEN_4383;
  wire        _GEN_4417 = _GEN_1319 | _GEN_1320;
  wire        _GEN_4418 = _GEN_1317 ? (_GEN_4417 ? (|lcam_ldq_idx_1) & _GEN_4385 : ~(_GEN_1315 & ~(|lcam_ldq_idx_1)) & _GEN_4385) : _GEN_4385;
  wire        _GEN_4419 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_336 & _GEN_4386 : ~(_GEN_1315 & _GEN_336) & _GEN_4386) : _GEN_4386;
  wire        _GEN_4420 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_337 & _GEN_4387 : ~(_GEN_1315 & _GEN_337) & _GEN_4387) : _GEN_4387;
  wire        _GEN_4421 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_338 & _GEN_4388 : ~(_GEN_1315 & _GEN_338) & _GEN_4388) : _GEN_4388;
  wire        _GEN_4422 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_339 & _GEN_4389 : ~(_GEN_1315 & _GEN_339) & _GEN_4389) : _GEN_4389;
  wire        _GEN_4423 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_340 & _GEN_4390 : ~(_GEN_1315 & _GEN_340) & _GEN_4390) : _GEN_4390;
  wire        _GEN_4424 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_341 & _GEN_4391 : ~(_GEN_1315 & _GEN_341) & _GEN_4391) : _GEN_4391;
  wire        _GEN_4425 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_342 & _GEN_4392 : ~(_GEN_1315 & _GEN_342) & _GEN_4392) : _GEN_4392;
  wire        _GEN_4426 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_343 & _GEN_4393 : ~(_GEN_1315 & _GEN_343) & _GEN_4393) : _GEN_4393;
  wire        _GEN_4427 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_344 & _GEN_4394 : ~(_GEN_1315 & _GEN_344) & _GEN_4394) : _GEN_4394;
  wire        _GEN_4428 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_345 & _GEN_4395 : ~(_GEN_1315 & _GEN_345) & _GEN_4395) : _GEN_4395;
  wire        _GEN_4429 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_346 & _GEN_4396 : ~(_GEN_1315 & _GEN_346) & _GEN_4396) : _GEN_4396;
  wire        _GEN_4430 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_347 & _GEN_4397 : ~(_GEN_1315 & _GEN_347) & _GEN_4397) : _GEN_4397;
  wire        _GEN_4431 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_348 & _GEN_4398 : ~(_GEN_1315 & _GEN_348) & _GEN_4398) : _GEN_4398;
  wire        _GEN_4432 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_349 & _GEN_4399 : ~(_GEN_1315 & _GEN_349) & _GEN_4399) : _GEN_4399;
  wire        _GEN_4433 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_350 & _GEN_4400 : ~(_GEN_1315 & _GEN_350) & _GEN_4400) : _GEN_4400;
  wire        _GEN_4434 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_351 & _GEN_4401 : ~(_GEN_1315 & _GEN_351) & _GEN_4401) : _GEN_4401;
  wire        _GEN_4435 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_352 & _GEN_4402 : ~(_GEN_1315 & _GEN_352) & _GEN_4402) : _GEN_4402;
  wire        _GEN_4436 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_353 & _GEN_4403 : ~(_GEN_1315 & _GEN_353) & _GEN_4403) : _GEN_4403;
  wire        _GEN_4437 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_354 & _GEN_4404 : ~(_GEN_1315 & _GEN_354) & _GEN_4404) : _GEN_4404;
  wire        _GEN_4438 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_355 & _GEN_4405 : ~(_GEN_1315 & _GEN_355) & _GEN_4405) : _GEN_4405;
  wire        _GEN_4439 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_356 & _GEN_4406 : ~(_GEN_1315 & _GEN_356) & _GEN_4406) : _GEN_4406;
  wire        _GEN_4440 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_357 & _GEN_4407 : ~(_GEN_1315 & _GEN_357) & _GEN_4407) : _GEN_4407;
  wire        _GEN_4441 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_358 & _GEN_4408 : ~(_GEN_1315 & _GEN_358) & _GEN_4408) : _GEN_4408;
  wire        _GEN_4442 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_359 & _GEN_4409 : ~(_GEN_1315 & _GEN_359) & _GEN_4409) : _GEN_4409;
  wire        _GEN_4443 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_360 & _GEN_4410 : ~(_GEN_1315 & _GEN_360) & _GEN_4410) : _GEN_4410;
  wire        _GEN_4444 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_361 & _GEN_4411 : ~(_GEN_1315 & _GEN_361) & _GEN_4411) : _GEN_4411;
  wire        _GEN_4445 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_362 & _GEN_4412 : ~(_GEN_1315 & _GEN_362) & _GEN_4412) : _GEN_4412;
  wire        _GEN_4446 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_363 & _GEN_4413 : ~(_GEN_1315 & _GEN_363) & _GEN_4413) : _GEN_4413;
  wire        _GEN_4447 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_364 & _GEN_4414 : ~(_GEN_1315 & _GEN_364) & _GEN_4414) : _GEN_4414;
  wire        _GEN_4448 = _GEN_1317 ? (_GEN_4417 ? ~_GEN_365 & _GEN_4415 : ~(_GEN_1315 & _GEN_365) & _GEN_4415) : _GEN_4415;
  wire        _GEN_4449 = _GEN_1317 ? (_GEN_4417 ? ~(&lcam_ldq_idx_1) & _GEN_4416 : ~(_GEN_1315 & (&lcam_ldq_idx_1)) & _GEN_4416) : _GEN_4416;
  wire        _GEN_4450 = _GEN_1324 | _GEN_1325;
  wire        _GEN_4451 = _GEN_1322 ? (_GEN_4450 ? (|lcam_ldq_idx_0) & _GEN_4418 : ~(_GEN_1326 & ~(|lcam_ldq_idx_0)) & _GEN_4418) : _GEN_4418;
  wire        _GEN_4452 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_296 & _GEN_4419 : ~(_GEN_1326 & _GEN_296) & _GEN_4419) : _GEN_4419;
  wire        _GEN_4453 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_297 & _GEN_4420 : ~(_GEN_1326 & _GEN_297) & _GEN_4420) : _GEN_4420;
  wire        _GEN_4454 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_298 & _GEN_4421 : ~(_GEN_1326 & _GEN_298) & _GEN_4421) : _GEN_4421;
  wire        _GEN_4455 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_299 & _GEN_4422 : ~(_GEN_1326 & _GEN_299) & _GEN_4422) : _GEN_4422;
  wire        _GEN_4456 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_300 & _GEN_4423 : ~(_GEN_1326 & _GEN_300) & _GEN_4423) : _GEN_4423;
  wire        _GEN_4457 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_301 & _GEN_4424 : ~(_GEN_1326 & _GEN_301) & _GEN_4424) : _GEN_4424;
  wire        _GEN_4458 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_302 & _GEN_4425 : ~(_GEN_1326 & _GEN_302) & _GEN_4425) : _GEN_4425;
  wire        _GEN_4459 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_303 & _GEN_4426 : ~(_GEN_1326 & _GEN_303) & _GEN_4426) : _GEN_4426;
  wire        _GEN_4460 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_304 & _GEN_4427 : ~(_GEN_1326 & _GEN_304) & _GEN_4427) : _GEN_4427;
  wire        _GEN_4461 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_305 & _GEN_4428 : ~(_GEN_1326 & _GEN_305) & _GEN_4428) : _GEN_4428;
  wire        _GEN_4462 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_306 & _GEN_4429 : ~(_GEN_1326 & _GEN_306) & _GEN_4429) : _GEN_4429;
  wire        _GEN_4463 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_307 & _GEN_4430 : ~(_GEN_1326 & _GEN_307) & _GEN_4430) : _GEN_4430;
  wire        _GEN_4464 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_308 & _GEN_4431 : ~(_GEN_1326 & _GEN_308) & _GEN_4431) : _GEN_4431;
  wire        _GEN_4465 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_309 & _GEN_4432 : ~(_GEN_1326 & _GEN_309) & _GEN_4432) : _GEN_4432;
  wire        _GEN_4466 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_310 & _GEN_4433 : ~(_GEN_1326 & _GEN_310) & _GEN_4433) : _GEN_4433;
  wire        _GEN_4467 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_311 & _GEN_4434 : ~(_GEN_1326 & _GEN_311) & _GEN_4434) : _GEN_4434;
  wire        _GEN_4468 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_312 & _GEN_4435 : ~(_GEN_1326 & _GEN_312) & _GEN_4435) : _GEN_4435;
  wire        _GEN_4469 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_313 & _GEN_4436 : ~(_GEN_1326 & _GEN_313) & _GEN_4436) : _GEN_4436;
  wire        _GEN_4470 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_314 & _GEN_4437 : ~(_GEN_1326 & _GEN_314) & _GEN_4437) : _GEN_4437;
  wire        _GEN_4471 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_315 & _GEN_4438 : ~(_GEN_1326 & _GEN_315) & _GEN_4438) : _GEN_4438;
  wire        _GEN_4472 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_316 & _GEN_4439 : ~(_GEN_1326 & _GEN_316) & _GEN_4439) : _GEN_4439;
  wire        _GEN_4473 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_317 & _GEN_4440 : ~(_GEN_1326 & _GEN_317) & _GEN_4440) : _GEN_4440;
  wire        _GEN_4474 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_318 & _GEN_4441 : ~(_GEN_1326 & _GEN_318) & _GEN_4441) : _GEN_4441;
  wire        _GEN_4475 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_319 & _GEN_4442 : ~(_GEN_1326 & _GEN_319) & _GEN_4442) : _GEN_4442;
  wire        _GEN_4476 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_320 & _GEN_4443 : ~(_GEN_1326 & _GEN_320) & _GEN_4443) : _GEN_4443;
  wire        _GEN_4477 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_321 & _GEN_4444 : ~(_GEN_1326 & _GEN_321) & _GEN_4444) : _GEN_4444;
  wire        _GEN_4478 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_322 & _GEN_4445 : ~(_GEN_1326 & _GEN_322) & _GEN_4445) : _GEN_4445;
  wire        _GEN_4479 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_323 & _GEN_4446 : ~(_GEN_1326 & _GEN_323) & _GEN_4446) : _GEN_4446;
  wire        _GEN_4480 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_324 & _GEN_4447 : ~(_GEN_1326 & _GEN_324) & _GEN_4447) : _GEN_4447;
  wire        _GEN_4481 = _GEN_1322 ? (_GEN_4450 ? ~_GEN_325 & _GEN_4448 : ~(_GEN_1326 & _GEN_325) & _GEN_4448) : _GEN_4448;
  wire        _GEN_4482 = _GEN_1322 ? (_GEN_4450 ? ~(&lcam_ldq_idx_0) & _GEN_4449 : ~(_GEN_1326 & (&lcam_ldq_idx_0)) & _GEN_4449) : _GEN_4449;
  wire        _GEN_4483 = _GEN_1330 | _GEN_1331;
  wire        _GEN_4484 = _GEN_1328 ? (_GEN_4483 ? (|lcam_ldq_idx_1) & _GEN_4451 : ~(_GEN_1326 & ~(|lcam_ldq_idx_1)) & _GEN_4451) : _GEN_4451;
  wire        _GEN_4485 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_336 & _GEN_4452 : ~(_GEN_1326 & _GEN_336) & _GEN_4452) : _GEN_4452;
  wire        _GEN_4486 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_337 & _GEN_4453 : ~(_GEN_1326 & _GEN_337) & _GEN_4453) : _GEN_4453;
  wire        _GEN_4487 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_338 & _GEN_4454 : ~(_GEN_1326 & _GEN_338) & _GEN_4454) : _GEN_4454;
  wire        _GEN_4488 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_339 & _GEN_4455 : ~(_GEN_1326 & _GEN_339) & _GEN_4455) : _GEN_4455;
  wire        _GEN_4489 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_340 & _GEN_4456 : ~(_GEN_1326 & _GEN_340) & _GEN_4456) : _GEN_4456;
  wire        _GEN_4490 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_341 & _GEN_4457 : ~(_GEN_1326 & _GEN_341) & _GEN_4457) : _GEN_4457;
  wire        _GEN_4491 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_342 & _GEN_4458 : ~(_GEN_1326 & _GEN_342) & _GEN_4458) : _GEN_4458;
  wire        _GEN_4492 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_343 & _GEN_4459 : ~(_GEN_1326 & _GEN_343) & _GEN_4459) : _GEN_4459;
  wire        _GEN_4493 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_344 & _GEN_4460 : ~(_GEN_1326 & _GEN_344) & _GEN_4460) : _GEN_4460;
  wire        _GEN_4494 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_345 & _GEN_4461 : ~(_GEN_1326 & _GEN_345) & _GEN_4461) : _GEN_4461;
  wire        _GEN_4495 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_346 & _GEN_4462 : ~(_GEN_1326 & _GEN_346) & _GEN_4462) : _GEN_4462;
  wire        _GEN_4496 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_347 & _GEN_4463 : ~(_GEN_1326 & _GEN_347) & _GEN_4463) : _GEN_4463;
  wire        _GEN_4497 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_348 & _GEN_4464 : ~(_GEN_1326 & _GEN_348) & _GEN_4464) : _GEN_4464;
  wire        _GEN_4498 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_349 & _GEN_4465 : ~(_GEN_1326 & _GEN_349) & _GEN_4465) : _GEN_4465;
  wire        _GEN_4499 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_350 & _GEN_4466 : ~(_GEN_1326 & _GEN_350) & _GEN_4466) : _GEN_4466;
  wire        _GEN_4500 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_351 & _GEN_4467 : ~(_GEN_1326 & _GEN_351) & _GEN_4467) : _GEN_4467;
  wire        _GEN_4501 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_352 & _GEN_4468 : ~(_GEN_1326 & _GEN_352) & _GEN_4468) : _GEN_4468;
  wire        _GEN_4502 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_353 & _GEN_4469 : ~(_GEN_1326 & _GEN_353) & _GEN_4469) : _GEN_4469;
  wire        _GEN_4503 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_354 & _GEN_4470 : ~(_GEN_1326 & _GEN_354) & _GEN_4470) : _GEN_4470;
  wire        _GEN_4504 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_355 & _GEN_4471 : ~(_GEN_1326 & _GEN_355) & _GEN_4471) : _GEN_4471;
  wire        _GEN_4505 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_356 & _GEN_4472 : ~(_GEN_1326 & _GEN_356) & _GEN_4472) : _GEN_4472;
  wire        _GEN_4506 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_357 & _GEN_4473 : ~(_GEN_1326 & _GEN_357) & _GEN_4473) : _GEN_4473;
  wire        _GEN_4507 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_358 & _GEN_4474 : ~(_GEN_1326 & _GEN_358) & _GEN_4474) : _GEN_4474;
  wire        _GEN_4508 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_359 & _GEN_4475 : ~(_GEN_1326 & _GEN_359) & _GEN_4475) : _GEN_4475;
  wire        _GEN_4509 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_360 & _GEN_4476 : ~(_GEN_1326 & _GEN_360) & _GEN_4476) : _GEN_4476;
  wire        _GEN_4510 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_361 & _GEN_4477 : ~(_GEN_1326 & _GEN_361) & _GEN_4477) : _GEN_4477;
  wire        _GEN_4511 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_362 & _GEN_4478 : ~(_GEN_1326 & _GEN_362) & _GEN_4478) : _GEN_4478;
  wire        _GEN_4512 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_363 & _GEN_4479 : ~(_GEN_1326 & _GEN_363) & _GEN_4479) : _GEN_4479;
  wire        _GEN_4513 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_364 & _GEN_4480 : ~(_GEN_1326 & _GEN_364) & _GEN_4480) : _GEN_4480;
  wire        _GEN_4514 = _GEN_1328 ? (_GEN_4483 ? ~_GEN_365 & _GEN_4481 : ~(_GEN_1326 & _GEN_365) & _GEN_4481) : _GEN_4481;
  wire        _GEN_4515 = _GEN_1328 ? (_GEN_4483 ? ~(&lcam_ldq_idx_1) & _GEN_4482 : ~(_GEN_1326 & (&lcam_ldq_idx_1)) & _GEN_4482) : _GEN_4482;
  wire        _GEN_4516 = _GEN_1335 | _GEN_1336;
  wire        _GEN_4517 = _GEN_1333 ? (_GEN_4516 ? (|lcam_ldq_idx_0) & _GEN_4484 : ~(_GEN_1337 & ~(|lcam_ldq_idx_0)) & _GEN_4484) : _GEN_4484;
  wire        _GEN_4518 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_296 & _GEN_4485 : ~(_GEN_1337 & _GEN_296) & _GEN_4485) : _GEN_4485;
  wire        _GEN_4519 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_297 & _GEN_4486 : ~(_GEN_1337 & _GEN_297) & _GEN_4486) : _GEN_4486;
  wire        _GEN_4520 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_298 & _GEN_4487 : ~(_GEN_1337 & _GEN_298) & _GEN_4487) : _GEN_4487;
  wire        _GEN_4521 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_299 & _GEN_4488 : ~(_GEN_1337 & _GEN_299) & _GEN_4488) : _GEN_4488;
  wire        _GEN_4522 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_300 & _GEN_4489 : ~(_GEN_1337 & _GEN_300) & _GEN_4489) : _GEN_4489;
  wire        _GEN_4523 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_301 & _GEN_4490 : ~(_GEN_1337 & _GEN_301) & _GEN_4490) : _GEN_4490;
  wire        _GEN_4524 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_302 & _GEN_4491 : ~(_GEN_1337 & _GEN_302) & _GEN_4491) : _GEN_4491;
  wire        _GEN_4525 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_303 & _GEN_4492 : ~(_GEN_1337 & _GEN_303) & _GEN_4492) : _GEN_4492;
  wire        _GEN_4526 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_304 & _GEN_4493 : ~(_GEN_1337 & _GEN_304) & _GEN_4493) : _GEN_4493;
  wire        _GEN_4527 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_305 & _GEN_4494 : ~(_GEN_1337 & _GEN_305) & _GEN_4494) : _GEN_4494;
  wire        _GEN_4528 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_306 & _GEN_4495 : ~(_GEN_1337 & _GEN_306) & _GEN_4495) : _GEN_4495;
  wire        _GEN_4529 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_307 & _GEN_4496 : ~(_GEN_1337 & _GEN_307) & _GEN_4496) : _GEN_4496;
  wire        _GEN_4530 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_308 & _GEN_4497 : ~(_GEN_1337 & _GEN_308) & _GEN_4497) : _GEN_4497;
  wire        _GEN_4531 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_309 & _GEN_4498 : ~(_GEN_1337 & _GEN_309) & _GEN_4498) : _GEN_4498;
  wire        _GEN_4532 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_310 & _GEN_4499 : ~(_GEN_1337 & _GEN_310) & _GEN_4499) : _GEN_4499;
  wire        _GEN_4533 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_311 & _GEN_4500 : ~(_GEN_1337 & _GEN_311) & _GEN_4500) : _GEN_4500;
  wire        _GEN_4534 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_312 & _GEN_4501 : ~(_GEN_1337 & _GEN_312) & _GEN_4501) : _GEN_4501;
  wire        _GEN_4535 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_313 & _GEN_4502 : ~(_GEN_1337 & _GEN_313) & _GEN_4502) : _GEN_4502;
  wire        _GEN_4536 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_314 & _GEN_4503 : ~(_GEN_1337 & _GEN_314) & _GEN_4503) : _GEN_4503;
  wire        _GEN_4537 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_315 & _GEN_4504 : ~(_GEN_1337 & _GEN_315) & _GEN_4504) : _GEN_4504;
  wire        _GEN_4538 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_316 & _GEN_4505 : ~(_GEN_1337 & _GEN_316) & _GEN_4505) : _GEN_4505;
  wire        _GEN_4539 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_317 & _GEN_4506 : ~(_GEN_1337 & _GEN_317) & _GEN_4506) : _GEN_4506;
  wire        _GEN_4540 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_318 & _GEN_4507 : ~(_GEN_1337 & _GEN_318) & _GEN_4507) : _GEN_4507;
  wire        _GEN_4541 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_319 & _GEN_4508 : ~(_GEN_1337 & _GEN_319) & _GEN_4508) : _GEN_4508;
  wire        _GEN_4542 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_320 & _GEN_4509 : ~(_GEN_1337 & _GEN_320) & _GEN_4509) : _GEN_4509;
  wire        _GEN_4543 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_321 & _GEN_4510 : ~(_GEN_1337 & _GEN_321) & _GEN_4510) : _GEN_4510;
  wire        _GEN_4544 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_322 & _GEN_4511 : ~(_GEN_1337 & _GEN_322) & _GEN_4511) : _GEN_4511;
  wire        _GEN_4545 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_323 & _GEN_4512 : ~(_GEN_1337 & _GEN_323) & _GEN_4512) : _GEN_4512;
  wire        _GEN_4546 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_324 & _GEN_4513 : ~(_GEN_1337 & _GEN_324) & _GEN_4513) : _GEN_4513;
  wire        _GEN_4547 = _GEN_1333 ? (_GEN_4516 ? ~_GEN_325 & _GEN_4514 : ~(_GEN_1337 & _GEN_325) & _GEN_4514) : _GEN_4514;
  wire        _GEN_4548 = _GEN_1333 ? (_GEN_4516 ? ~(&lcam_ldq_idx_0) & _GEN_4515 : ~(_GEN_1337 & (&lcam_ldq_idx_0)) & _GEN_4515) : _GEN_4515;
  wire        _GEN_4549 = _GEN_1341 | _GEN_1342;
  wire        _GEN_4550 = _GEN_1339 ? (_GEN_4549 ? (|lcam_ldq_idx_1) & _GEN_4517 : ~(_GEN_1337 & ~(|lcam_ldq_idx_1)) & _GEN_4517) : _GEN_4517;
  wire        _GEN_4551 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_336 & _GEN_4518 : ~(_GEN_1337 & _GEN_336) & _GEN_4518) : _GEN_4518;
  wire        _GEN_4552 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_337 & _GEN_4519 : ~(_GEN_1337 & _GEN_337) & _GEN_4519) : _GEN_4519;
  wire        _GEN_4553 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_338 & _GEN_4520 : ~(_GEN_1337 & _GEN_338) & _GEN_4520) : _GEN_4520;
  wire        _GEN_4554 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_339 & _GEN_4521 : ~(_GEN_1337 & _GEN_339) & _GEN_4521) : _GEN_4521;
  wire        _GEN_4555 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_340 & _GEN_4522 : ~(_GEN_1337 & _GEN_340) & _GEN_4522) : _GEN_4522;
  wire        _GEN_4556 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_341 & _GEN_4523 : ~(_GEN_1337 & _GEN_341) & _GEN_4523) : _GEN_4523;
  wire        _GEN_4557 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_342 & _GEN_4524 : ~(_GEN_1337 & _GEN_342) & _GEN_4524) : _GEN_4524;
  wire        _GEN_4558 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_343 & _GEN_4525 : ~(_GEN_1337 & _GEN_343) & _GEN_4525) : _GEN_4525;
  wire        _GEN_4559 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_344 & _GEN_4526 : ~(_GEN_1337 & _GEN_344) & _GEN_4526) : _GEN_4526;
  wire        _GEN_4560 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_345 & _GEN_4527 : ~(_GEN_1337 & _GEN_345) & _GEN_4527) : _GEN_4527;
  wire        _GEN_4561 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_346 & _GEN_4528 : ~(_GEN_1337 & _GEN_346) & _GEN_4528) : _GEN_4528;
  wire        _GEN_4562 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_347 & _GEN_4529 : ~(_GEN_1337 & _GEN_347) & _GEN_4529) : _GEN_4529;
  wire        _GEN_4563 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_348 & _GEN_4530 : ~(_GEN_1337 & _GEN_348) & _GEN_4530) : _GEN_4530;
  wire        _GEN_4564 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_349 & _GEN_4531 : ~(_GEN_1337 & _GEN_349) & _GEN_4531) : _GEN_4531;
  wire        _GEN_4565 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_350 & _GEN_4532 : ~(_GEN_1337 & _GEN_350) & _GEN_4532) : _GEN_4532;
  wire        _GEN_4566 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_351 & _GEN_4533 : ~(_GEN_1337 & _GEN_351) & _GEN_4533) : _GEN_4533;
  wire        _GEN_4567 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_352 & _GEN_4534 : ~(_GEN_1337 & _GEN_352) & _GEN_4534) : _GEN_4534;
  wire        _GEN_4568 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_353 & _GEN_4535 : ~(_GEN_1337 & _GEN_353) & _GEN_4535) : _GEN_4535;
  wire        _GEN_4569 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_354 & _GEN_4536 : ~(_GEN_1337 & _GEN_354) & _GEN_4536) : _GEN_4536;
  wire        _GEN_4570 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_355 & _GEN_4537 : ~(_GEN_1337 & _GEN_355) & _GEN_4537) : _GEN_4537;
  wire        _GEN_4571 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_356 & _GEN_4538 : ~(_GEN_1337 & _GEN_356) & _GEN_4538) : _GEN_4538;
  wire        _GEN_4572 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_357 & _GEN_4539 : ~(_GEN_1337 & _GEN_357) & _GEN_4539) : _GEN_4539;
  wire        _GEN_4573 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_358 & _GEN_4540 : ~(_GEN_1337 & _GEN_358) & _GEN_4540) : _GEN_4540;
  wire        _GEN_4574 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_359 & _GEN_4541 : ~(_GEN_1337 & _GEN_359) & _GEN_4541) : _GEN_4541;
  wire        _GEN_4575 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_360 & _GEN_4542 : ~(_GEN_1337 & _GEN_360) & _GEN_4542) : _GEN_4542;
  wire        _GEN_4576 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_361 & _GEN_4543 : ~(_GEN_1337 & _GEN_361) & _GEN_4543) : _GEN_4543;
  wire        _GEN_4577 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_362 & _GEN_4544 : ~(_GEN_1337 & _GEN_362) & _GEN_4544) : _GEN_4544;
  wire        _GEN_4578 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_363 & _GEN_4545 : ~(_GEN_1337 & _GEN_363) & _GEN_4545) : _GEN_4545;
  wire        _GEN_4579 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_364 & _GEN_4546 : ~(_GEN_1337 & _GEN_364) & _GEN_4546) : _GEN_4546;
  wire        _GEN_4580 = _GEN_1339 ? (_GEN_4549 ? ~_GEN_365 & _GEN_4547 : ~(_GEN_1337 & _GEN_365) & _GEN_4547) : _GEN_4547;
  wire        _GEN_4581 = _GEN_1339 ? (_GEN_4549 ? ~(&lcam_ldq_idx_1) & _GEN_4548 : ~(_GEN_1337 & (&lcam_ldq_idx_1)) & _GEN_4548) : _GEN_4548;
  wire        _GEN_4582 = _GEN_1346 | _GEN_1347;
  wire        _GEN_4583 = _GEN_1344 ? (_GEN_4582 ? (|lcam_ldq_idx_0) & _GEN_4550 : ~(_GEN_1348 & ~(|lcam_ldq_idx_0)) & _GEN_4550) : _GEN_4550;
  wire        _GEN_4584 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_296 & _GEN_4551 : ~(_GEN_1348 & _GEN_296) & _GEN_4551) : _GEN_4551;
  wire        _GEN_4585 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_297 & _GEN_4552 : ~(_GEN_1348 & _GEN_297) & _GEN_4552) : _GEN_4552;
  wire        _GEN_4586 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_298 & _GEN_4553 : ~(_GEN_1348 & _GEN_298) & _GEN_4553) : _GEN_4553;
  wire        _GEN_4587 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_299 & _GEN_4554 : ~(_GEN_1348 & _GEN_299) & _GEN_4554) : _GEN_4554;
  wire        _GEN_4588 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_300 & _GEN_4555 : ~(_GEN_1348 & _GEN_300) & _GEN_4555) : _GEN_4555;
  wire        _GEN_4589 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_301 & _GEN_4556 : ~(_GEN_1348 & _GEN_301) & _GEN_4556) : _GEN_4556;
  wire        _GEN_4590 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_302 & _GEN_4557 : ~(_GEN_1348 & _GEN_302) & _GEN_4557) : _GEN_4557;
  wire        _GEN_4591 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_303 & _GEN_4558 : ~(_GEN_1348 & _GEN_303) & _GEN_4558) : _GEN_4558;
  wire        _GEN_4592 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_304 & _GEN_4559 : ~(_GEN_1348 & _GEN_304) & _GEN_4559) : _GEN_4559;
  wire        _GEN_4593 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_305 & _GEN_4560 : ~(_GEN_1348 & _GEN_305) & _GEN_4560) : _GEN_4560;
  wire        _GEN_4594 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_306 & _GEN_4561 : ~(_GEN_1348 & _GEN_306) & _GEN_4561) : _GEN_4561;
  wire        _GEN_4595 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_307 & _GEN_4562 : ~(_GEN_1348 & _GEN_307) & _GEN_4562) : _GEN_4562;
  wire        _GEN_4596 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_308 & _GEN_4563 : ~(_GEN_1348 & _GEN_308) & _GEN_4563) : _GEN_4563;
  wire        _GEN_4597 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_309 & _GEN_4564 : ~(_GEN_1348 & _GEN_309) & _GEN_4564) : _GEN_4564;
  wire        _GEN_4598 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_310 & _GEN_4565 : ~(_GEN_1348 & _GEN_310) & _GEN_4565) : _GEN_4565;
  wire        _GEN_4599 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_311 & _GEN_4566 : ~(_GEN_1348 & _GEN_311) & _GEN_4566) : _GEN_4566;
  wire        _GEN_4600 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_312 & _GEN_4567 : ~(_GEN_1348 & _GEN_312) & _GEN_4567) : _GEN_4567;
  wire        _GEN_4601 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_313 & _GEN_4568 : ~(_GEN_1348 & _GEN_313) & _GEN_4568) : _GEN_4568;
  wire        _GEN_4602 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_314 & _GEN_4569 : ~(_GEN_1348 & _GEN_314) & _GEN_4569) : _GEN_4569;
  wire        _GEN_4603 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_315 & _GEN_4570 : ~(_GEN_1348 & _GEN_315) & _GEN_4570) : _GEN_4570;
  wire        _GEN_4604 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_316 & _GEN_4571 : ~(_GEN_1348 & _GEN_316) & _GEN_4571) : _GEN_4571;
  wire        _GEN_4605 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_317 & _GEN_4572 : ~(_GEN_1348 & _GEN_317) & _GEN_4572) : _GEN_4572;
  wire        _GEN_4606 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_318 & _GEN_4573 : ~(_GEN_1348 & _GEN_318) & _GEN_4573) : _GEN_4573;
  wire        _GEN_4607 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_319 & _GEN_4574 : ~(_GEN_1348 & _GEN_319) & _GEN_4574) : _GEN_4574;
  wire        _GEN_4608 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_320 & _GEN_4575 : ~(_GEN_1348 & _GEN_320) & _GEN_4575) : _GEN_4575;
  wire        _GEN_4609 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_321 & _GEN_4576 : ~(_GEN_1348 & _GEN_321) & _GEN_4576) : _GEN_4576;
  wire        _GEN_4610 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_322 & _GEN_4577 : ~(_GEN_1348 & _GEN_322) & _GEN_4577) : _GEN_4577;
  wire        _GEN_4611 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_323 & _GEN_4578 : ~(_GEN_1348 & _GEN_323) & _GEN_4578) : _GEN_4578;
  wire        _GEN_4612 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_324 & _GEN_4579 : ~(_GEN_1348 & _GEN_324) & _GEN_4579) : _GEN_4579;
  wire        _GEN_4613 = _GEN_1344 ? (_GEN_4582 ? ~_GEN_325 & _GEN_4580 : ~(_GEN_1348 & _GEN_325) & _GEN_4580) : _GEN_4580;
  wire        _GEN_4614 = _GEN_1344 ? (_GEN_4582 ? ~(&lcam_ldq_idx_0) & _GEN_4581 : ~(_GEN_1348 & (&lcam_ldq_idx_0)) & _GEN_4581) : _GEN_4581;
  wire        _GEN_4615 = _GEN_1352 | _GEN_1353;
  wire        _GEN_4616 = _GEN_1350 ? (_GEN_4615 ? (|lcam_ldq_idx_1) & _GEN_4583 : ~(_GEN_1348 & ~(|lcam_ldq_idx_1)) & _GEN_4583) : _GEN_4583;
  wire        _GEN_4617 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_336 & _GEN_4584 : ~(_GEN_1348 & _GEN_336) & _GEN_4584) : _GEN_4584;
  wire        _GEN_4618 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_337 & _GEN_4585 : ~(_GEN_1348 & _GEN_337) & _GEN_4585) : _GEN_4585;
  wire        _GEN_4619 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_338 & _GEN_4586 : ~(_GEN_1348 & _GEN_338) & _GEN_4586) : _GEN_4586;
  wire        _GEN_4620 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_339 & _GEN_4587 : ~(_GEN_1348 & _GEN_339) & _GEN_4587) : _GEN_4587;
  wire        _GEN_4621 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_340 & _GEN_4588 : ~(_GEN_1348 & _GEN_340) & _GEN_4588) : _GEN_4588;
  wire        _GEN_4622 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_341 & _GEN_4589 : ~(_GEN_1348 & _GEN_341) & _GEN_4589) : _GEN_4589;
  wire        _GEN_4623 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_342 & _GEN_4590 : ~(_GEN_1348 & _GEN_342) & _GEN_4590) : _GEN_4590;
  wire        _GEN_4624 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_343 & _GEN_4591 : ~(_GEN_1348 & _GEN_343) & _GEN_4591) : _GEN_4591;
  wire        _GEN_4625 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_344 & _GEN_4592 : ~(_GEN_1348 & _GEN_344) & _GEN_4592) : _GEN_4592;
  wire        _GEN_4626 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_345 & _GEN_4593 : ~(_GEN_1348 & _GEN_345) & _GEN_4593) : _GEN_4593;
  wire        _GEN_4627 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_346 & _GEN_4594 : ~(_GEN_1348 & _GEN_346) & _GEN_4594) : _GEN_4594;
  wire        _GEN_4628 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_347 & _GEN_4595 : ~(_GEN_1348 & _GEN_347) & _GEN_4595) : _GEN_4595;
  wire        _GEN_4629 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_348 & _GEN_4596 : ~(_GEN_1348 & _GEN_348) & _GEN_4596) : _GEN_4596;
  wire        _GEN_4630 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_349 & _GEN_4597 : ~(_GEN_1348 & _GEN_349) & _GEN_4597) : _GEN_4597;
  wire        _GEN_4631 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_350 & _GEN_4598 : ~(_GEN_1348 & _GEN_350) & _GEN_4598) : _GEN_4598;
  wire        _GEN_4632 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_351 & _GEN_4599 : ~(_GEN_1348 & _GEN_351) & _GEN_4599) : _GEN_4599;
  wire        _GEN_4633 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_352 & _GEN_4600 : ~(_GEN_1348 & _GEN_352) & _GEN_4600) : _GEN_4600;
  wire        _GEN_4634 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_353 & _GEN_4601 : ~(_GEN_1348 & _GEN_353) & _GEN_4601) : _GEN_4601;
  wire        _GEN_4635 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_354 & _GEN_4602 : ~(_GEN_1348 & _GEN_354) & _GEN_4602) : _GEN_4602;
  wire        _GEN_4636 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_355 & _GEN_4603 : ~(_GEN_1348 & _GEN_355) & _GEN_4603) : _GEN_4603;
  wire        _GEN_4637 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_356 & _GEN_4604 : ~(_GEN_1348 & _GEN_356) & _GEN_4604) : _GEN_4604;
  wire        _GEN_4638 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_357 & _GEN_4605 : ~(_GEN_1348 & _GEN_357) & _GEN_4605) : _GEN_4605;
  wire        _GEN_4639 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_358 & _GEN_4606 : ~(_GEN_1348 & _GEN_358) & _GEN_4606) : _GEN_4606;
  wire        _GEN_4640 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_359 & _GEN_4607 : ~(_GEN_1348 & _GEN_359) & _GEN_4607) : _GEN_4607;
  wire        _GEN_4641 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_360 & _GEN_4608 : ~(_GEN_1348 & _GEN_360) & _GEN_4608) : _GEN_4608;
  wire        _GEN_4642 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_361 & _GEN_4609 : ~(_GEN_1348 & _GEN_361) & _GEN_4609) : _GEN_4609;
  wire        _GEN_4643 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_362 & _GEN_4610 : ~(_GEN_1348 & _GEN_362) & _GEN_4610) : _GEN_4610;
  wire        _GEN_4644 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_363 & _GEN_4611 : ~(_GEN_1348 & _GEN_363) & _GEN_4611) : _GEN_4611;
  wire        _GEN_4645 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_364 & _GEN_4612 : ~(_GEN_1348 & _GEN_364) & _GEN_4612) : _GEN_4612;
  wire        _GEN_4646 = _GEN_1350 ? (_GEN_4615 ? ~_GEN_365 & _GEN_4613 : ~(_GEN_1348 & _GEN_365) & _GEN_4613) : _GEN_4613;
  wire        _GEN_4647 = _GEN_1350 ? (_GEN_4615 ? ~(&lcam_ldq_idx_1) & _GEN_4614 : ~(_GEN_1348 & (&lcam_ldq_idx_1)) & _GEN_4614) : _GEN_4614;
  wire        _GEN_4648 = _GEN_1357 | _GEN_1358;
  wire        _GEN_4649 = _GEN_1355 ? (_GEN_4648 ? (|lcam_ldq_idx_0) & _GEN_4616 : ~(_GEN_1359 & ~(|lcam_ldq_idx_0)) & _GEN_4616) : _GEN_4616;
  wire        _GEN_4650 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_296 & _GEN_4617 : ~(_GEN_1359 & _GEN_296) & _GEN_4617) : _GEN_4617;
  wire        _GEN_4651 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_297 & _GEN_4618 : ~(_GEN_1359 & _GEN_297) & _GEN_4618) : _GEN_4618;
  wire        _GEN_4652 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_298 & _GEN_4619 : ~(_GEN_1359 & _GEN_298) & _GEN_4619) : _GEN_4619;
  wire        _GEN_4653 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_299 & _GEN_4620 : ~(_GEN_1359 & _GEN_299) & _GEN_4620) : _GEN_4620;
  wire        _GEN_4654 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_300 & _GEN_4621 : ~(_GEN_1359 & _GEN_300) & _GEN_4621) : _GEN_4621;
  wire        _GEN_4655 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_301 & _GEN_4622 : ~(_GEN_1359 & _GEN_301) & _GEN_4622) : _GEN_4622;
  wire        _GEN_4656 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_302 & _GEN_4623 : ~(_GEN_1359 & _GEN_302) & _GEN_4623) : _GEN_4623;
  wire        _GEN_4657 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_303 & _GEN_4624 : ~(_GEN_1359 & _GEN_303) & _GEN_4624) : _GEN_4624;
  wire        _GEN_4658 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_304 & _GEN_4625 : ~(_GEN_1359 & _GEN_304) & _GEN_4625) : _GEN_4625;
  wire        _GEN_4659 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_305 & _GEN_4626 : ~(_GEN_1359 & _GEN_305) & _GEN_4626) : _GEN_4626;
  wire        _GEN_4660 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_306 & _GEN_4627 : ~(_GEN_1359 & _GEN_306) & _GEN_4627) : _GEN_4627;
  wire        _GEN_4661 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_307 & _GEN_4628 : ~(_GEN_1359 & _GEN_307) & _GEN_4628) : _GEN_4628;
  wire        _GEN_4662 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_308 & _GEN_4629 : ~(_GEN_1359 & _GEN_308) & _GEN_4629) : _GEN_4629;
  wire        _GEN_4663 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_309 & _GEN_4630 : ~(_GEN_1359 & _GEN_309) & _GEN_4630) : _GEN_4630;
  wire        _GEN_4664 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_310 & _GEN_4631 : ~(_GEN_1359 & _GEN_310) & _GEN_4631) : _GEN_4631;
  wire        _GEN_4665 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_311 & _GEN_4632 : ~(_GEN_1359 & _GEN_311) & _GEN_4632) : _GEN_4632;
  wire        _GEN_4666 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_312 & _GEN_4633 : ~(_GEN_1359 & _GEN_312) & _GEN_4633) : _GEN_4633;
  wire        _GEN_4667 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_313 & _GEN_4634 : ~(_GEN_1359 & _GEN_313) & _GEN_4634) : _GEN_4634;
  wire        _GEN_4668 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_314 & _GEN_4635 : ~(_GEN_1359 & _GEN_314) & _GEN_4635) : _GEN_4635;
  wire        _GEN_4669 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_315 & _GEN_4636 : ~(_GEN_1359 & _GEN_315) & _GEN_4636) : _GEN_4636;
  wire        _GEN_4670 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_316 & _GEN_4637 : ~(_GEN_1359 & _GEN_316) & _GEN_4637) : _GEN_4637;
  wire        _GEN_4671 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_317 & _GEN_4638 : ~(_GEN_1359 & _GEN_317) & _GEN_4638) : _GEN_4638;
  wire        _GEN_4672 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_318 & _GEN_4639 : ~(_GEN_1359 & _GEN_318) & _GEN_4639) : _GEN_4639;
  wire        _GEN_4673 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_319 & _GEN_4640 : ~(_GEN_1359 & _GEN_319) & _GEN_4640) : _GEN_4640;
  wire        _GEN_4674 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_320 & _GEN_4641 : ~(_GEN_1359 & _GEN_320) & _GEN_4641) : _GEN_4641;
  wire        _GEN_4675 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_321 & _GEN_4642 : ~(_GEN_1359 & _GEN_321) & _GEN_4642) : _GEN_4642;
  wire        _GEN_4676 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_322 & _GEN_4643 : ~(_GEN_1359 & _GEN_322) & _GEN_4643) : _GEN_4643;
  wire        _GEN_4677 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_323 & _GEN_4644 : ~(_GEN_1359 & _GEN_323) & _GEN_4644) : _GEN_4644;
  wire        _GEN_4678 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_324 & _GEN_4645 : ~(_GEN_1359 & _GEN_324) & _GEN_4645) : _GEN_4645;
  wire        _GEN_4679 = _GEN_1355 ? (_GEN_4648 ? ~_GEN_325 & _GEN_4646 : ~(_GEN_1359 & _GEN_325) & _GEN_4646) : _GEN_4646;
  wire        _GEN_4680 = _GEN_1355 ? (_GEN_4648 ? ~(&lcam_ldq_idx_0) & _GEN_4647 : ~(_GEN_1359 & (&lcam_ldq_idx_0)) & _GEN_4647) : _GEN_4647;
  wire        _GEN_4681 = _GEN_1363 | _GEN_1364;
  wire        _GEN_4682 = _GEN_1361 ? (_GEN_4681 ? (|lcam_ldq_idx_1) & _GEN_4649 : ~(_GEN_1359 & ~(|lcam_ldq_idx_1)) & _GEN_4649) : _GEN_4649;
  wire        _GEN_4683 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_336 & _GEN_4650 : ~(_GEN_1359 & _GEN_336) & _GEN_4650) : _GEN_4650;
  wire        _GEN_4684 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_337 & _GEN_4651 : ~(_GEN_1359 & _GEN_337) & _GEN_4651) : _GEN_4651;
  wire        _GEN_4685 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_338 & _GEN_4652 : ~(_GEN_1359 & _GEN_338) & _GEN_4652) : _GEN_4652;
  wire        _GEN_4686 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_339 & _GEN_4653 : ~(_GEN_1359 & _GEN_339) & _GEN_4653) : _GEN_4653;
  wire        _GEN_4687 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_340 & _GEN_4654 : ~(_GEN_1359 & _GEN_340) & _GEN_4654) : _GEN_4654;
  wire        _GEN_4688 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_341 & _GEN_4655 : ~(_GEN_1359 & _GEN_341) & _GEN_4655) : _GEN_4655;
  wire        _GEN_4689 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_342 & _GEN_4656 : ~(_GEN_1359 & _GEN_342) & _GEN_4656) : _GEN_4656;
  wire        _GEN_4690 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_343 & _GEN_4657 : ~(_GEN_1359 & _GEN_343) & _GEN_4657) : _GEN_4657;
  wire        _GEN_4691 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_344 & _GEN_4658 : ~(_GEN_1359 & _GEN_344) & _GEN_4658) : _GEN_4658;
  wire        _GEN_4692 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_345 & _GEN_4659 : ~(_GEN_1359 & _GEN_345) & _GEN_4659) : _GEN_4659;
  wire        _GEN_4693 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_346 & _GEN_4660 : ~(_GEN_1359 & _GEN_346) & _GEN_4660) : _GEN_4660;
  wire        _GEN_4694 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_347 & _GEN_4661 : ~(_GEN_1359 & _GEN_347) & _GEN_4661) : _GEN_4661;
  wire        _GEN_4695 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_348 & _GEN_4662 : ~(_GEN_1359 & _GEN_348) & _GEN_4662) : _GEN_4662;
  wire        _GEN_4696 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_349 & _GEN_4663 : ~(_GEN_1359 & _GEN_349) & _GEN_4663) : _GEN_4663;
  wire        _GEN_4697 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_350 & _GEN_4664 : ~(_GEN_1359 & _GEN_350) & _GEN_4664) : _GEN_4664;
  wire        _GEN_4698 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_351 & _GEN_4665 : ~(_GEN_1359 & _GEN_351) & _GEN_4665) : _GEN_4665;
  wire        _GEN_4699 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_352 & _GEN_4666 : ~(_GEN_1359 & _GEN_352) & _GEN_4666) : _GEN_4666;
  wire        _GEN_4700 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_353 & _GEN_4667 : ~(_GEN_1359 & _GEN_353) & _GEN_4667) : _GEN_4667;
  wire        _GEN_4701 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_354 & _GEN_4668 : ~(_GEN_1359 & _GEN_354) & _GEN_4668) : _GEN_4668;
  wire        _GEN_4702 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_355 & _GEN_4669 : ~(_GEN_1359 & _GEN_355) & _GEN_4669) : _GEN_4669;
  wire        _GEN_4703 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_356 & _GEN_4670 : ~(_GEN_1359 & _GEN_356) & _GEN_4670) : _GEN_4670;
  wire        _GEN_4704 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_357 & _GEN_4671 : ~(_GEN_1359 & _GEN_357) & _GEN_4671) : _GEN_4671;
  wire        _GEN_4705 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_358 & _GEN_4672 : ~(_GEN_1359 & _GEN_358) & _GEN_4672) : _GEN_4672;
  wire        _GEN_4706 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_359 & _GEN_4673 : ~(_GEN_1359 & _GEN_359) & _GEN_4673) : _GEN_4673;
  wire        _GEN_4707 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_360 & _GEN_4674 : ~(_GEN_1359 & _GEN_360) & _GEN_4674) : _GEN_4674;
  wire        _GEN_4708 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_361 & _GEN_4675 : ~(_GEN_1359 & _GEN_361) & _GEN_4675) : _GEN_4675;
  wire        _GEN_4709 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_362 & _GEN_4676 : ~(_GEN_1359 & _GEN_362) & _GEN_4676) : _GEN_4676;
  wire        _GEN_4710 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_363 & _GEN_4677 : ~(_GEN_1359 & _GEN_363) & _GEN_4677) : _GEN_4677;
  wire        _GEN_4711 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_364 & _GEN_4678 : ~(_GEN_1359 & _GEN_364) & _GEN_4678) : _GEN_4678;
  wire        _GEN_4712 = _GEN_1361 ? (_GEN_4681 ? ~_GEN_365 & _GEN_4679 : ~(_GEN_1359 & _GEN_365) & _GEN_4679) : _GEN_4679;
  wire        _GEN_4713 = _GEN_1361 ? (_GEN_4681 ? ~(&lcam_ldq_idx_1) & _GEN_4680 : ~(_GEN_1359 & (&lcam_ldq_idx_1)) & _GEN_4680) : _GEN_4680;
  wire        _GEN_4714 = _GEN_1368 | _GEN_1369;
  wire        _GEN_4715 = _GEN_1366 ? (_GEN_4714 ? (|lcam_ldq_idx_0) & _GEN_4682 : ~(_GEN_1370 & ~(|lcam_ldq_idx_0)) & _GEN_4682) : _GEN_4682;
  wire        _GEN_4716 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_296 & _GEN_4683 : ~(_GEN_1370 & _GEN_296) & _GEN_4683) : _GEN_4683;
  wire        _GEN_4717 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_297 & _GEN_4684 : ~(_GEN_1370 & _GEN_297) & _GEN_4684) : _GEN_4684;
  wire        _GEN_4718 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_298 & _GEN_4685 : ~(_GEN_1370 & _GEN_298) & _GEN_4685) : _GEN_4685;
  wire        _GEN_4719 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_299 & _GEN_4686 : ~(_GEN_1370 & _GEN_299) & _GEN_4686) : _GEN_4686;
  wire        _GEN_4720 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_300 & _GEN_4687 : ~(_GEN_1370 & _GEN_300) & _GEN_4687) : _GEN_4687;
  wire        _GEN_4721 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_301 & _GEN_4688 : ~(_GEN_1370 & _GEN_301) & _GEN_4688) : _GEN_4688;
  wire        _GEN_4722 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_302 & _GEN_4689 : ~(_GEN_1370 & _GEN_302) & _GEN_4689) : _GEN_4689;
  wire        _GEN_4723 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_303 & _GEN_4690 : ~(_GEN_1370 & _GEN_303) & _GEN_4690) : _GEN_4690;
  wire        _GEN_4724 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_304 & _GEN_4691 : ~(_GEN_1370 & _GEN_304) & _GEN_4691) : _GEN_4691;
  wire        _GEN_4725 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_305 & _GEN_4692 : ~(_GEN_1370 & _GEN_305) & _GEN_4692) : _GEN_4692;
  wire        _GEN_4726 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_306 & _GEN_4693 : ~(_GEN_1370 & _GEN_306) & _GEN_4693) : _GEN_4693;
  wire        _GEN_4727 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_307 & _GEN_4694 : ~(_GEN_1370 & _GEN_307) & _GEN_4694) : _GEN_4694;
  wire        _GEN_4728 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_308 & _GEN_4695 : ~(_GEN_1370 & _GEN_308) & _GEN_4695) : _GEN_4695;
  wire        _GEN_4729 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_309 & _GEN_4696 : ~(_GEN_1370 & _GEN_309) & _GEN_4696) : _GEN_4696;
  wire        _GEN_4730 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_310 & _GEN_4697 : ~(_GEN_1370 & _GEN_310) & _GEN_4697) : _GEN_4697;
  wire        _GEN_4731 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_311 & _GEN_4698 : ~(_GEN_1370 & _GEN_311) & _GEN_4698) : _GEN_4698;
  wire        _GEN_4732 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_312 & _GEN_4699 : ~(_GEN_1370 & _GEN_312) & _GEN_4699) : _GEN_4699;
  wire        _GEN_4733 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_313 & _GEN_4700 : ~(_GEN_1370 & _GEN_313) & _GEN_4700) : _GEN_4700;
  wire        _GEN_4734 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_314 & _GEN_4701 : ~(_GEN_1370 & _GEN_314) & _GEN_4701) : _GEN_4701;
  wire        _GEN_4735 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_315 & _GEN_4702 : ~(_GEN_1370 & _GEN_315) & _GEN_4702) : _GEN_4702;
  wire        _GEN_4736 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_316 & _GEN_4703 : ~(_GEN_1370 & _GEN_316) & _GEN_4703) : _GEN_4703;
  wire        _GEN_4737 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_317 & _GEN_4704 : ~(_GEN_1370 & _GEN_317) & _GEN_4704) : _GEN_4704;
  wire        _GEN_4738 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_318 & _GEN_4705 : ~(_GEN_1370 & _GEN_318) & _GEN_4705) : _GEN_4705;
  wire        _GEN_4739 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_319 & _GEN_4706 : ~(_GEN_1370 & _GEN_319) & _GEN_4706) : _GEN_4706;
  wire        _GEN_4740 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_320 & _GEN_4707 : ~(_GEN_1370 & _GEN_320) & _GEN_4707) : _GEN_4707;
  wire        _GEN_4741 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_321 & _GEN_4708 : ~(_GEN_1370 & _GEN_321) & _GEN_4708) : _GEN_4708;
  wire        _GEN_4742 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_322 & _GEN_4709 : ~(_GEN_1370 & _GEN_322) & _GEN_4709) : _GEN_4709;
  wire        _GEN_4743 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_323 & _GEN_4710 : ~(_GEN_1370 & _GEN_323) & _GEN_4710) : _GEN_4710;
  wire        _GEN_4744 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_324 & _GEN_4711 : ~(_GEN_1370 & _GEN_324) & _GEN_4711) : _GEN_4711;
  wire        _GEN_4745 = _GEN_1366 ? (_GEN_4714 ? ~_GEN_325 & _GEN_4712 : ~(_GEN_1370 & _GEN_325) & _GEN_4712) : _GEN_4712;
  wire        _GEN_4746 = _GEN_1366 ? (_GEN_4714 ? ~(&lcam_ldq_idx_0) & _GEN_4713 : ~(_GEN_1370 & (&lcam_ldq_idx_0)) & _GEN_4713) : _GEN_4713;
  wire        _GEN_4747 = _GEN_1374 | _GEN_1375;
  wire        _GEN_4748 = _GEN_1372 ? (_GEN_4747 ? (|lcam_ldq_idx_1) & _GEN_4715 : ~(_GEN_1370 & ~(|lcam_ldq_idx_1)) & _GEN_4715) : _GEN_4715;
  wire        _GEN_4749 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_336 & _GEN_4716 : ~(_GEN_1370 & _GEN_336) & _GEN_4716) : _GEN_4716;
  wire        _GEN_4750 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_337 & _GEN_4717 : ~(_GEN_1370 & _GEN_337) & _GEN_4717) : _GEN_4717;
  wire        _GEN_4751 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_338 & _GEN_4718 : ~(_GEN_1370 & _GEN_338) & _GEN_4718) : _GEN_4718;
  wire        _GEN_4752 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_339 & _GEN_4719 : ~(_GEN_1370 & _GEN_339) & _GEN_4719) : _GEN_4719;
  wire        _GEN_4753 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_340 & _GEN_4720 : ~(_GEN_1370 & _GEN_340) & _GEN_4720) : _GEN_4720;
  wire        _GEN_4754 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_341 & _GEN_4721 : ~(_GEN_1370 & _GEN_341) & _GEN_4721) : _GEN_4721;
  wire        _GEN_4755 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_342 & _GEN_4722 : ~(_GEN_1370 & _GEN_342) & _GEN_4722) : _GEN_4722;
  wire        _GEN_4756 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_343 & _GEN_4723 : ~(_GEN_1370 & _GEN_343) & _GEN_4723) : _GEN_4723;
  wire        _GEN_4757 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_344 & _GEN_4724 : ~(_GEN_1370 & _GEN_344) & _GEN_4724) : _GEN_4724;
  wire        _GEN_4758 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_345 & _GEN_4725 : ~(_GEN_1370 & _GEN_345) & _GEN_4725) : _GEN_4725;
  wire        _GEN_4759 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_346 & _GEN_4726 : ~(_GEN_1370 & _GEN_346) & _GEN_4726) : _GEN_4726;
  wire        _GEN_4760 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_347 & _GEN_4727 : ~(_GEN_1370 & _GEN_347) & _GEN_4727) : _GEN_4727;
  wire        _GEN_4761 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_348 & _GEN_4728 : ~(_GEN_1370 & _GEN_348) & _GEN_4728) : _GEN_4728;
  wire        _GEN_4762 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_349 & _GEN_4729 : ~(_GEN_1370 & _GEN_349) & _GEN_4729) : _GEN_4729;
  wire        _GEN_4763 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_350 & _GEN_4730 : ~(_GEN_1370 & _GEN_350) & _GEN_4730) : _GEN_4730;
  wire        _GEN_4764 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_351 & _GEN_4731 : ~(_GEN_1370 & _GEN_351) & _GEN_4731) : _GEN_4731;
  wire        _GEN_4765 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_352 & _GEN_4732 : ~(_GEN_1370 & _GEN_352) & _GEN_4732) : _GEN_4732;
  wire        _GEN_4766 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_353 & _GEN_4733 : ~(_GEN_1370 & _GEN_353) & _GEN_4733) : _GEN_4733;
  wire        _GEN_4767 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_354 & _GEN_4734 : ~(_GEN_1370 & _GEN_354) & _GEN_4734) : _GEN_4734;
  wire        _GEN_4768 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_355 & _GEN_4735 : ~(_GEN_1370 & _GEN_355) & _GEN_4735) : _GEN_4735;
  wire        _GEN_4769 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_356 & _GEN_4736 : ~(_GEN_1370 & _GEN_356) & _GEN_4736) : _GEN_4736;
  wire        _GEN_4770 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_357 & _GEN_4737 : ~(_GEN_1370 & _GEN_357) & _GEN_4737) : _GEN_4737;
  wire        _GEN_4771 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_358 & _GEN_4738 : ~(_GEN_1370 & _GEN_358) & _GEN_4738) : _GEN_4738;
  wire        _GEN_4772 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_359 & _GEN_4739 : ~(_GEN_1370 & _GEN_359) & _GEN_4739) : _GEN_4739;
  wire        _GEN_4773 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_360 & _GEN_4740 : ~(_GEN_1370 & _GEN_360) & _GEN_4740) : _GEN_4740;
  wire        _GEN_4774 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_361 & _GEN_4741 : ~(_GEN_1370 & _GEN_361) & _GEN_4741) : _GEN_4741;
  wire        _GEN_4775 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_362 & _GEN_4742 : ~(_GEN_1370 & _GEN_362) & _GEN_4742) : _GEN_4742;
  wire        _GEN_4776 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_363 & _GEN_4743 : ~(_GEN_1370 & _GEN_363) & _GEN_4743) : _GEN_4743;
  wire        _GEN_4777 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_364 & _GEN_4744 : ~(_GEN_1370 & _GEN_364) & _GEN_4744) : _GEN_4744;
  wire        _GEN_4778 = _GEN_1372 ? (_GEN_4747 ? ~_GEN_365 & _GEN_4745 : ~(_GEN_1370 & _GEN_365) & _GEN_4745) : _GEN_4745;
  wire        _GEN_4779 = _GEN_1372 ? (_GEN_4747 ? ~(&lcam_ldq_idx_1) & _GEN_4746 : ~(_GEN_1370 & (&lcam_ldq_idx_1)) & _GEN_4746) : _GEN_4746;
  wire        _GEN_4780 = _GEN_1379 | _GEN_1380;
  wire        _GEN_4781 = _GEN_1377 ? (_GEN_4780 ? (|lcam_ldq_idx_0) & _GEN_4748 : ~(_GEN_1381 & ~(|lcam_ldq_idx_0)) & _GEN_4748) : _GEN_4748;
  wire        _GEN_4782 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_296 & _GEN_4749 : ~(_GEN_1381 & _GEN_296) & _GEN_4749) : _GEN_4749;
  wire        _GEN_4783 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_297 & _GEN_4750 : ~(_GEN_1381 & _GEN_297) & _GEN_4750) : _GEN_4750;
  wire        _GEN_4784 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_298 & _GEN_4751 : ~(_GEN_1381 & _GEN_298) & _GEN_4751) : _GEN_4751;
  wire        _GEN_4785 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_299 & _GEN_4752 : ~(_GEN_1381 & _GEN_299) & _GEN_4752) : _GEN_4752;
  wire        _GEN_4786 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_300 & _GEN_4753 : ~(_GEN_1381 & _GEN_300) & _GEN_4753) : _GEN_4753;
  wire        _GEN_4787 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_301 & _GEN_4754 : ~(_GEN_1381 & _GEN_301) & _GEN_4754) : _GEN_4754;
  wire        _GEN_4788 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_302 & _GEN_4755 : ~(_GEN_1381 & _GEN_302) & _GEN_4755) : _GEN_4755;
  wire        _GEN_4789 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_303 & _GEN_4756 : ~(_GEN_1381 & _GEN_303) & _GEN_4756) : _GEN_4756;
  wire        _GEN_4790 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_304 & _GEN_4757 : ~(_GEN_1381 & _GEN_304) & _GEN_4757) : _GEN_4757;
  wire        _GEN_4791 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_305 & _GEN_4758 : ~(_GEN_1381 & _GEN_305) & _GEN_4758) : _GEN_4758;
  wire        _GEN_4792 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_306 & _GEN_4759 : ~(_GEN_1381 & _GEN_306) & _GEN_4759) : _GEN_4759;
  wire        _GEN_4793 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_307 & _GEN_4760 : ~(_GEN_1381 & _GEN_307) & _GEN_4760) : _GEN_4760;
  wire        _GEN_4794 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_308 & _GEN_4761 : ~(_GEN_1381 & _GEN_308) & _GEN_4761) : _GEN_4761;
  wire        _GEN_4795 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_309 & _GEN_4762 : ~(_GEN_1381 & _GEN_309) & _GEN_4762) : _GEN_4762;
  wire        _GEN_4796 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_310 & _GEN_4763 : ~(_GEN_1381 & _GEN_310) & _GEN_4763) : _GEN_4763;
  wire        _GEN_4797 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_311 & _GEN_4764 : ~(_GEN_1381 & _GEN_311) & _GEN_4764) : _GEN_4764;
  wire        _GEN_4798 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_312 & _GEN_4765 : ~(_GEN_1381 & _GEN_312) & _GEN_4765) : _GEN_4765;
  wire        _GEN_4799 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_313 & _GEN_4766 : ~(_GEN_1381 & _GEN_313) & _GEN_4766) : _GEN_4766;
  wire        _GEN_4800 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_314 & _GEN_4767 : ~(_GEN_1381 & _GEN_314) & _GEN_4767) : _GEN_4767;
  wire        _GEN_4801 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_315 & _GEN_4768 : ~(_GEN_1381 & _GEN_315) & _GEN_4768) : _GEN_4768;
  wire        _GEN_4802 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_316 & _GEN_4769 : ~(_GEN_1381 & _GEN_316) & _GEN_4769) : _GEN_4769;
  wire        _GEN_4803 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_317 & _GEN_4770 : ~(_GEN_1381 & _GEN_317) & _GEN_4770) : _GEN_4770;
  wire        _GEN_4804 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_318 & _GEN_4771 : ~(_GEN_1381 & _GEN_318) & _GEN_4771) : _GEN_4771;
  wire        _GEN_4805 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_319 & _GEN_4772 : ~(_GEN_1381 & _GEN_319) & _GEN_4772) : _GEN_4772;
  wire        _GEN_4806 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_320 & _GEN_4773 : ~(_GEN_1381 & _GEN_320) & _GEN_4773) : _GEN_4773;
  wire        _GEN_4807 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_321 & _GEN_4774 : ~(_GEN_1381 & _GEN_321) & _GEN_4774) : _GEN_4774;
  wire        _GEN_4808 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_322 & _GEN_4775 : ~(_GEN_1381 & _GEN_322) & _GEN_4775) : _GEN_4775;
  wire        _GEN_4809 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_323 & _GEN_4776 : ~(_GEN_1381 & _GEN_323) & _GEN_4776) : _GEN_4776;
  wire        _GEN_4810 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_324 & _GEN_4777 : ~(_GEN_1381 & _GEN_324) & _GEN_4777) : _GEN_4777;
  wire        _GEN_4811 = _GEN_1377 ? (_GEN_4780 ? ~_GEN_325 & _GEN_4778 : ~(_GEN_1381 & _GEN_325) & _GEN_4778) : _GEN_4778;
  wire        _GEN_4812 = _GEN_1377 ? (_GEN_4780 ? ~(&lcam_ldq_idx_0) & _GEN_4779 : ~(_GEN_1381 & (&lcam_ldq_idx_0)) & _GEN_4779) : _GEN_4779;
  wire        _GEN_4813 = _GEN_1385 | _GEN_1386;
  wire        _GEN_4814 = _GEN_1383 ? (_GEN_4813 ? (|lcam_ldq_idx_1) & _GEN_4781 : ~(_GEN_1381 & ~(|lcam_ldq_idx_1)) & _GEN_4781) : _GEN_4781;
  wire        _GEN_4815 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_336 & _GEN_4782 : ~(_GEN_1381 & _GEN_336) & _GEN_4782) : _GEN_4782;
  wire        _GEN_4816 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_337 & _GEN_4783 : ~(_GEN_1381 & _GEN_337) & _GEN_4783) : _GEN_4783;
  wire        _GEN_4817 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_338 & _GEN_4784 : ~(_GEN_1381 & _GEN_338) & _GEN_4784) : _GEN_4784;
  wire        _GEN_4818 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_339 & _GEN_4785 : ~(_GEN_1381 & _GEN_339) & _GEN_4785) : _GEN_4785;
  wire        _GEN_4819 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_340 & _GEN_4786 : ~(_GEN_1381 & _GEN_340) & _GEN_4786) : _GEN_4786;
  wire        _GEN_4820 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_341 & _GEN_4787 : ~(_GEN_1381 & _GEN_341) & _GEN_4787) : _GEN_4787;
  wire        _GEN_4821 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_342 & _GEN_4788 : ~(_GEN_1381 & _GEN_342) & _GEN_4788) : _GEN_4788;
  wire        _GEN_4822 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_343 & _GEN_4789 : ~(_GEN_1381 & _GEN_343) & _GEN_4789) : _GEN_4789;
  wire        _GEN_4823 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_344 & _GEN_4790 : ~(_GEN_1381 & _GEN_344) & _GEN_4790) : _GEN_4790;
  wire        _GEN_4824 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_345 & _GEN_4791 : ~(_GEN_1381 & _GEN_345) & _GEN_4791) : _GEN_4791;
  wire        _GEN_4825 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_346 & _GEN_4792 : ~(_GEN_1381 & _GEN_346) & _GEN_4792) : _GEN_4792;
  wire        _GEN_4826 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_347 & _GEN_4793 : ~(_GEN_1381 & _GEN_347) & _GEN_4793) : _GEN_4793;
  wire        _GEN_4827 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_348 & _GEN_4794 : ~(_GEN_1381 & _GEN_348) & _GEN_4794) : _GEN_4794;
  wire        _GEN_4828 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_349 & _GEN_4795 : ~(_GEN_1381 & _GEN_349) & _GEN_4795) : _GEN_4795;
  wire        _GEN_4829 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_350 & _GEN_4796 : ~(_GEN_1381 & _GEN_350) & _GEN_4796) : _GEN_4796;
  wire        _GEN_4830 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_351 & _GEN_4797 : ~(_GEN_1381 & _GEN_351) & _GEN_4797) : _GEN_4797;
  wire        _GEN_4831 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_352 & _GEN_4798 : ~(_GEN_1381 & _GEN_352) & _GEN_4798) : _GEN_4798;
  wire        _GEN_4832 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_353 & _GEN_4799 : ~(_GEN_1381 & _GEN_353) & _GEN_4799) : _GEN_4799;
  wire        _GEN_4833 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_354 & _GEN_4800 : ~(_GEN_1381 & _GEN_354) & _GEN_4800) : _GEN_4800;
  wire        _GEN_4834 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_355 & _GEN_4801 : ~(_GEN_1381 & _GEN_355) & _GEN_4801) : _GEN_4801;
  wire        _GEN_4835 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_356 & _GEN_4802 : ~(_GEN_1381 & _GEN_356) & _GEN_4802) : _GEN_4802;
  wire        _GEN_4836 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_357 & _GEN_4803 : ~(_GEN_1381 & _GEN_357) & _GEN_4803) : _GEN_4803;
  wire        _GEN_4837 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_358 & _GEN_4804 : ~(_GEN_1381 & _GEN_358) & _GEN_4804) : _GEN_4804;
  wire        _GEN_4838 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_359 & _GEN_4805 : ~(_GEN_1381 & _GEN_359) & _GEN_4805) : _GEN_4805;
  wire        _GEN_4839 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_360 & _GEN_4806 : ~(_GEN_1381 & _GEN_360) & _GEN_4806) : _GEN_4806;
  wire        _GEN_4840 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_361 & _GEN_4807 : ~(_GEN_1381 & _GEN_361) & _GEN_4807) : _GEN_4807;
  wire        _GEN_4841 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_362 & _GEN_4808 : ~(_GEN_1381 & _GEN_362) & _GEN_4808) : _GEN_4808;
  wire        _GEN_4842 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_363 & _GEN_4809 : ~(_GEN_1381 & _GEN_363) & _GEN_4809) : _GEN_4809;
  wire        _GEN_4843 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_364 & _GEN_4810 : ~(_GEN_1381 & _GEN_364) & _GEN_4810) : _GEN_4810;
  wire        _GEN_4844 = _GEN_1383 ? (_GEN_4813 ? ~_GEN_365 & _GEN_4811 : ~(_GEN_1381 & _GEN_365) & _GEN_4811) : _GEN_4811;
  wire        _GEN_4845 = _GEN_1383 ? (_GEN_4813 ? ~(&lcam_ldq_idx_1) & _GEN_4812 : ~(_GEN_1381 & (&lcam_ldq_idx_1)) & _GEN_4812) : _GEN_4812;
  wire        _GEN_4846 = _GEN_1390 | _GEN_1391;
  wire        _GEN_4847 = _GEN_1388 ? (_GEN_4846 ? (|lcam_ldq_idx_0) & _GEN_4814 : ~(_GEN_1392 & ~(|lcam_ldq_idx_0)) & _GEN_4814) : _GEN_4814;
  wire        _GEN_4848 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_296 & _GEN_4815 : ~(_GEN_1392 & _GEN_296) & _GEN_4815) : _GEN_4815;
  wire        _GEN_4849 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_297 & _GEN_4816 : ~(_GEN_1392 & _GEN_297) & _GEN_4816) : _GEN_4816;
  wire        _GEN_4850 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_298 & _GEN_4817 : ~(_GEN_1392 & _GEN_298) & _GEN_4817) : _GEN_4817;
  wire        _GEN_4851 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_299 & _GEN_4818 : ~(_GEN_1392 & _GEN_299) & _GEN_4818) : _GEN_4818;
  wire        _GEN_4852 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_300 & _GEN_4819 : ~(_GEN_1392 & _GEN_300) & _GEN_4819) : _GEN_4819;
  wire        _GEN_4853 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_301 & _GEN_4820 : ~(_GEN_1392 & _GEN_301) & _GEN_4820) : _GEN_4820;
  wire        _GEN_4854 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_302 & _GEN_4821 : ~(_GEN_1392 & _GEN_302) & _GEN_4821) : _GEN_4821;
  wire        _GEN_4855 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_303 & _GEN_4822 : ~(_GEN_1392 & _GEN_303) & _GEN_4822) : _GEN_4822;
  wire        _GEN_4856 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_304 & _GEN_4823 : ~(_GEN_1392 & _GEN_304) & _GEN_4823) : _GEN_4823;
  wire        _GEN_4857 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_305 & _GEN_4824 : ~(_GEN_1392 & _GEN_305) & _GEN_4824) : _GEN_4824;
  wire        _GEN_4858 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_306 & _GEN_4825 : ~(_GEN_1392 & _GEN_306) & _GEN_4825) : _GEN_4825;
  wire        _GEN_4859 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_307 & _GEN_4826 : ~(_GEN_1392 & _GEN_307) & _GEN_4826) : _GEN_4826;
  wire        _GEN_4860 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_308 & _GEN_4827 : ~(_GEN_1392 & _GEN_308) & _GEN_4827) : _GEN_4827;
  wire        _GEN_4861 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_309 & _GEN_4828 : ~(_GEN_1392 & _GEN_309) & _GEN_4828) : _GEN_4828;
  wire        _GEN_4862 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_310 & _GEN_4829 : ~(_GEN_1392 & _GEN_310) & _GEN_4829) : _GEN_4829;
  wire        _GEN_4863 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_311 & _GEN_4830 : ~(_GEN_1392 & _GEN_311) & _GEN_4830) : _GEN_4830;
  wire        _GEN_4864 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_312 & _GEN_4831 : ~(_GEN_1392 & _GEN_312) & _GEN_4831) : _GEN_4831;
  wire        _GEN_4865 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_313 & _GEN_4832 : ~(_GEN_1392 & _GEN_313) & _GEN_4832) : _GEN_4832;
  wire        _GEN_4866 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_314 & _GEN_4833 : ~(_GEN_1392 & _GEN_314) & _GEN_4833) : _GEN_4833;
  wire        _GEN_4867 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_315 & _GEN_4834 : ~(_GEN_1392 & _GEN_315) & _GEN_4834) : _GEN_4834;
  wire        _GEN_4868 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_316 & _GEN_4835 : ~(_GEN_1392 & _GEN_316) & _GEN_4835) : _GEN_4835;
  wire        _GEN_4869 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_317 & _GEN_4836 : ~(_GEN_1392 & _GEN_317) & _GEN_4836) : _GEN_4836;
  wire        _GEN_4870 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_318 & _GEN_4837 : ~(_GEN_1392 & _GEN_318) & _GEN_4837) : _GEN_4837;
  wire        _GEN_4871 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_319 & _GEN_4838 : ~(_GEN_1392 & _GEN_319) & _GEN_4838) : _GEN_4838;
  wire        _GEN_4872 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_320 & _GEN_4839 : ~(_GEN_1392 & _GEN_320) & _GEN_4839) : _GEN_4839;
  wire        _GEN_4873 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_321 & _GEN_4840 : ~(_GEN_1392 & _GEN_321) & _GEN_4840) : _GEN_4840;
  wire        _GEN_4874 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_322 & _GEN_4841 : ~(_GEN_1392 & _GEN_322) & _GEN_4841) : _GEN_4841;
  wire        _GEN_4875 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_323 & _GEN_4842 : ~(_GEN_1392 & _GEN_323) & _GEN_4842) : _GEN_4842;
  wire        _GEN_4876 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_324 & _GEN_4843 : ~(_GEN_1392 & _GEN_324) & _GEN_4843) : _GEN_4843;
  wire        _GEN_4877 = _GEN_1388 ? (_GEN_4846 ? ~_GEN_325 & _GEN_4844 : ~(_GEN_1392 & _GEN_325) & _GEN_4844) : _GEN_4844;
  wire        _GEN_4878 = _GEN_1388 ? (_GEN_4846 ? ~(&lcam_ldq_idx_0) & _GEN_4845 : ~(_GEN_1392 & (&lcam_ldq_idx_0)) & _GEN_4845) : _GEN_4845;
  wire        _GEN_4879 = _GEN_1396 | _GEN_1397;
  wire        _GEN_4880 = _GEN_1394 ? (_GEN_4879 ? (|lcam_ldq_idx_1) & _GEN_4847 : ~(_GEN_1392 & ~(|lcam_ldq_idx_1)) & _GEN_4847) : _GEN_4847;
  wire        _GEN_4881 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_336 & _GEN_4848 : ~(_GEN_1392 & _GEN_336) & _GEN_4848) : _GEN_4848;
  wire        _GEN_4882 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_337 & _GEN_4849 : ~(_GEN_1392 & _GEN_337) & _GEN_4849) : _GEN_4849;
  wire        _GEN_4883 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_338 & _GEN_4850 : ~(_GEN_1392 & _GEN_338) & _GEN_4850) : _GEN_4850;
  wire        _GEN_4884 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_339 & _GEN_4851 : ~(_GEN_1392 & _GEN_339) & _GEN_4851) : _GEN_4851;
  wire        _GEN_4885 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_340 & _GEN_4852 : ~(_GEN_1392 & _GEN_340) & _GEN_4852) : _GEN_4852;
  wire        _GEN_4886 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_341 & _GEN_4853 : ~(_GEN_1392 & _GEN_341) & _GEN_4853) : _GEN_4853;
  wire        _GEN_4887 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_342 & _GEN_4854 : ~(_GEN_1392 & _GEN_342) & _GEN_4854) : _GEN_4854;
  wire        _GEN_4888 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_343 & _GEN_4855 : ~(_GEN_1392 & _GEN_343) & _GEN_4855) : _GEN_4855;
  wire        _GEN_4889 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_344 & _GEN_4856 : ~(_GEN_1392 & _GEN_344) & _GEN_4856) : _GEN_4856;
  wire        _GEN_4890 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_345 & _GEN_4857 : ~(_GEN_1392 & _GEN_345) & _GEN_4857) : _GEN_4857;
  wire        _GEN_4891 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_346 & _GEN_4858 : ~(_GEN_1392 & _GEN_346) & _GEN_4858) : _GEN_4858;
  wire        _GEN_4892 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_347 & _GEN_4859 : ~(_GEN_1392 & _GEN_347) & _GEN_4859) : _GEN_4859;
  wire        _GEN_4893 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_348 & _GEN_4860 : ~(_GEN_1392 & _GEN_348) & _GEN_4860) : _GEN_4860;
  wire        _GEN_4894 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_349 & _GEN_4861 : ~(_GEN_1392 & _GEN_349) & _GEN_4861) : _GEN_4861;
  wire        _GEN_4895 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_350 & _GEN_4862 : ~(_GEN_1392 & _GEN_350) & _GEN_4862) : _GEN_4862;
  wire        _GEN_4896 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_351 & _GEN_4863 : ~(_GEN_1392 & _GEN_351) & _GEN_4863) : _GEN_4863;
  wire        _GEN_4897 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_352 & _GEN_4864 : ~(_GEN_1392 & _GEN_352) & _GEN_4864) : _GEN_4864;
  wire        _GEN_4898 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_353 & _GEN_4865 : ~(_GEN_1392 & _GEN_353) & _GEN_4865) : _GEN_4865;
  wire        _GEN_4899 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_354 & _GEN_4866 : ~(_GEN_1392 & _GEN_354) & _GEN_4866) : _GEN_4866;
  wire        _GEN_4900 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_355 & _GEN_4867 : ~(_GEN_1392 & _GEN_355) & _GEN_4867) : _GEN_4867;
  wire        _GEN_4901 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_356 & _GEN_4868 : ~(_GEN_1392 & _GEN_356) & _GEN_4868) : _GEN_4868;
  wire        _GEN_4902 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_357 & _GEN_4869 : ~(_GEN_1392 & _GEN_357) & _GEN_4869) : _GEN_4869;
  wire        _GEN_4903 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_358 & _GEN_4870 : ~(_GEN_1392 & _GEN_358) & _GEN_4870) : _GEN_4870;
  wire        _GEN_4904 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_359 & _GEN_4871 : ~(_GEN_1392 & _GEN_359) & _GEN_4871) : _GEN_4871;
  wire        _GEN_4905 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_360 & _GEN_4872 : ~(_GEN_1392 & _GEN_360) & _GEN_4872) : _GEN_4872;
  wire        _GEN_4906 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_361 & _GEN_4873 : ~(_GEN_1392 & _GEN_361) & _GEN_4873) : _GEN_4873;
  wire        _GEN_4907 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_362 & _GEN_4874 : ~(_GEN_1392 & _GEN_362) & _GEN_4874) : _GEN_4874;
  wire        _GEN_4908 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_363 & _GEN_4875 : ~(_GEN_1392 & _GEN_363) & _GEN_4875) : _GEN_4875;
  wire        _GEN_4909 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_364 & _GEN_4876 : ~(_GEN_1392 & _GEN_364) & _GEN_4876) : _GEN_4876;
  wire        _GEN_4910 = _GEN_1394 ? (_GEN_4879 ? ~_GEN_365 & _GEN_4877 : ~(_GEN_1392 & _GEN_365) & _GEN_4877) : _GEN_4877;
  wire        _GEN_4911 = _GEN_1394 ? (_GEN_4879 ? ~(&lcam_ldq_idx_1) & _GEN_4878 : ~(_GEN_1392 & (&lcam_ldq_idx_1)) & _GEN_4878) : _GEN_4878;
  wire        _GEN_4912 = _GEN_1401 | _GEN_1402;
  wire        _GEN_4913 = _GEN_1399 ? (_GEN_4912 ? (|lcam_ldq_idx_0) & _GEN_4880 : ~(_GEN_1403 & ~(|lcam_ldq_idx_0)) & _GEN_4880) : _GEN_4880;
  wire        _GEN_4914 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_296 & _GEN_4881 : ~(_GEN_1403 & _GEN_296) & _GEN_4881) : _GEN_4881;
  wire        _GEN_4915 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_297 & _GEN_4882 : ~(_GEN_1403 & _GEN_297) & _GEN_4882) : _GEN_4882;
  wire        _GEN_4916 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_298 & _GEN_4883 : ~(_GEN_1403 & _GEN_298) & _GEN_4883) : _GEN_4883;
  wire        _GEN_4917 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_299 & _GEN_4884 : ~(_GEN_1403 & _GEN_299) & _GEN_4884) : _GEN_4884;
  wire        _GEN_4918 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_300 & _GEN_4885 : ~(_GEN_1403 & _GEN_300) & _GEN_4885) : _GEN_4885;
  wire        _GEN_4919 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_301 & _GEN_4886 : ~(_GEN_1403 & _GEN_301) & _GEN_4886) : _GEN_4886;
  wire        _GEN_4920 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_302 & _GEN_4887 : ~(_GEN_1403 & _GEN_302) & _GEN_4887) : _GEN_4887;
  wire        _GEN_4921 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_303 & _GEN_4888 : ~(_GEN_1403 & _GEN_303) & _GEN_4888) : _GEN_4888;
  wire        _GEN_4922 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_304 & _GEN_4889 : ~(_GEN_1403 & _GEN_304) & _GEN_4889) : _GEN_4889;
  wire        _GEN_4923 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_305 & _GEN_4890 : ~(_GEN_1403 & _GEN_305) & _GEN_4890) : _GEN_4890;
  wire        _GEN_4924 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_306 & _GEN_4891 : ~(_GEN_1403 & _GEN_306) & _GEN_4891) : _GEN_4891;
  wire        _GEN_4925 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_307 & _GEN_4892 : ~(_GEN_1403 & _GEN_307) & _GEN_4892) : _GEN_4892;
  wire        _GEN_4926 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_308 & _GEN_4893 : ~(_GEN_1403 & _GEN_308) & _GEN_4893) : _GEN_4893;
  wire        _GEN_4927 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_309 & _GEN_4894 : ~(_GEN_1403 & _GEN_309) & _GEN_4894) : _GEN_4894;
  wire        _GEN_4928 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_310 & _GEN_4895 : ~(_GEN_1403 & _GEN_310) & _GEN_4895) : _GEN_4895;
  wire        _GEN_4929 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_311 & _GEN_4896 : ~(_GEN_1403 & _GEN_311) & _GEN_4896) : _GEN_4896;
  wire        _GEN_4930 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_312 & _GEN_4897 : ~(_GEN_1403 & _GEN_312) & _GEN_4897) : _GEN_4897;
  wire        _GEN_4931 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_313 & _GEN_4898 : ~(_GEN_1403 & _GEN_313) & _GEN_4898) : _GEN_4898;
  wire        _GEN_4932 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_314 & _GEN_4899 : ~(_GEN_1403 & _GEN_314) & _GEN_4899) : _GEN_4899;
  wire        _GEN_4933 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_315 & _GEN_4900 : ~(_GEN_1403 & _GEN_315) & _GEN_4900) : _GEN_4900;
  wire        _GEN_4934 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_316 & _GEN_4901 : ~(_GEN_1403 & _GEN_316) & _GEN_4901) : _GEN_4901;
  wire        _GEN_4935 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_317 & _GEN_4902 : ~(_GEN_1403 & _GEN_317) & _GEN_4902) : _GEN_4902;
  wire        _GEN_4936 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_318 & _GEN_4903 : ~(_GEN_1403 & _GEN_318) & _GEN_4903) : _GEN_4903;
  wire        _GEN_4937 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_319 & _GEN_4904 : ~(_GEN_1403 & _GEN_319) & _GEN_4904) : _GEN_4904;
  wire        _GEN_4938 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_320 & _GEN_4905 : ~(_GEN_1403 & _GEN_320) & _GEN_4905) : _GEN_4905;
  wire        _GEN_4939 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_321 & _GEN_4906 : ~(_GEN_1403 & _GEN_321) & _GEN_4906) : _GEN_4906;
  wire        _GEN_4940 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_322 & _GEN_4907 : ~(_GEN_1403 & _GEN_322) & _GEN_4907) : _GEN_4907;
  wire        _GEN_4941 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_323 & _GEN_4908 : ~(_GEN_1403 & _GEN_323) & _GEN_4908) : _GEN_4908;
  wire        _GEN_4942 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_324 & _GEN_4909 : ~(_GEN_1403 & _GEN_324) & _GEN_4909) : _GEN_4909;
  wire        _GEN_4943 = _GEN_1399 ? (_GEN_4912 ? ~_GEN_325 & _GEN_4910 : ~(_GEN_1403 & _GEN_325) & _GEN_4910) : _GEN_4910;
  wire        _GEN_4944 = _GEN_1399 ? (_GEN_4912 ? ~(&lcam_ldq_idx_0) & _GEN_4911 : ~(_GEN_1403 & (&lcam_ldq_idx_0)) & _GEN_4911) : _GEN_4911;
  wire        _GEN_4945 = _GEN_1407 | _GEN_1408;
  wire        _GEN_4946 = _GEN_1405 ? (_GEN_4945 ? (|lcam_ldq_idx_1) & _GEN_4913 : ~(_GEN_1403 & ~(|lcam_ldq_idx_1)) & _GEN_4913) : _GEN_4913;
  wire        _GEN_4947 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_336 & _GEN_4914 : ~(_GEN_1403 & _GEN_336) & _GEN_4914) : _GEN_4914;
  wire        _GEN_4948 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_337 & _GEN_4915 : ~(_GEN_1403 & _GEN_337) & _GEN_4915) : _GEN_4915;
  wire        _GEN_4949 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_338 & _GEN_4916 : ~(_GEN_1403 & _GEN_338) & _GEN_4916) : _GEN_4916;
  wire        _GEN_4950 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_339 & _GEN_4917 : ~(_GEN_1403 & _GEN_339) & _GEN_4917) : _GEN_4917;
  wire        _GEN_4951 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_340 & _GEN_4918 : ~(_GEN_1403 & _GEN_340) & _GEN_4918) : _GEN_4918;
  wire        _GEN_4952 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_341 & _GEN_4919 : ~(_GEN_1403 & _GEN_341) & _GEN_4919) : _GEN_4919;
  wire        _GEN_4953 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_342 & _GEN_4920 : ~(_GEN_1403 & _GEN_342) & _GEN_4920) : _GEN_4920;
  wire        _GEN_4954 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_343 & _GEN_4921 : ~(_GEN_1403 & _GEN_343) & _GEN_4921) : _GEN_4921;
  wire        _GEN_4955 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_344 & _GEN_4922 : ~(_GEN_1403 & _GEN_344) & _GEN_4922) : _GEN_4922;
  wire        _GEN_4956 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_345 & _GEN_4923 : ~(_GEN_1403 & _GEN_345) & _GEN_4923) : _GEN_4923;
  wire        _GEN_4957 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_346 & _GEN_4924 : ~(_GEN_1403 & _GEN_346) & _GEN_4924) : _GEN_4924;
  wire        _GEN_4958 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_347 & _GEN_4925 : ~(_GEN_1403 & _GEN_347) & _GEN_4925) : _GEN_4925;
  wire        _GEN_4959 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_348 & _GEN_4926 : ~(_GEN_1403 & _GEN_348) & _GEN_4926) : _GEN_4926;
  wire        _GEN_4960 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_349 & _GEN_4927 : ~(_GEN_1403 & _GEN_349) & _GEN_4927) : _GEN_4927;
  wire        _GEN_4961 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_350 & _GEN_4928 : ~(_GEN_1403 & _GEN_350) & _GEN_4928) : _GEN_4928;
  wire        _GEN_4962 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_351 & _GEN_4929 : ~(_GEN_1403 & _GEN_351) & _GEN_4929) : _GEN_4929;
  wire        _GEN_4963 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_352 & _GEN_4930 : ~(_GEN_1403 & _GEN_352) & _GEN_4930) : _GEN_4930;
  wire        _GEN_4964 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_353 & _GEN_4931 : ~(_GEN_1403 & _GEN_353) & _GEN_4931) : _GEN_4931;
  wire        _GEN_4965 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_354 & _GEN_4932 : ~(_GEN_1403 & _GEN_354) & _GEN_4932) : _GEN_4932;
  wire        _GEN_4966 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_355 & _GEN_4933 : ~(_GEN_1403 & _GEN_355) & _GEN_4933) : _GEN_4933;
  wire        _GEN_4967 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_356 & _GEN_4934 : ~(_GEN_1403 & _GEN_356) & _GEN_4934) : _GEN_4934;
  wire        _GEN_4968 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_357 & _GEN_4935 : ~(_GEN_1403 & _GEN_357) & _GEN_4935) : _GEN_4935;
  wire        _GEN_4969 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_358 & _GEN_4936 : ~(_GEN_1403 & _GEN_358) & _GEN_4936) : _GEN_4936;
  wire        _GEN_4970 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_359 & _GEN_4937 : ~(_GEN_1403 & _GEN_359) & _GEN_4937) : _GEN_4937;
  wire        _GEN_4971 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_360 & _GEN_4938 : ~(_GEN_1403 & _GEN_360) & _GEN_4938) : _GEN_4938;
  wire        _GEN_4972 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_361 & _GEN_4939 : ~(_GEN_1403 & _GEN_361) & _GEN_4939) : _GEN_4939;
  wire        _GEN_4973 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_362 & _GEN_4940 : ~(_GEN_1403 & _GEN_362) & _GEN_4940) : _GEN_4940;
  wire        _GEN_4974 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_363 & _GEN_4941 : ~(_GEN_1403 & _GEN_363) & _GEN_4941) : _GEN_4941;
  wire        _GEN_4975 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_364 & _GEN_4942 : ~(_GEN_1403 & _GEN_364) & _GEN_4942) : _GEN_4942;
  wire        _GEN_4976 = _GEN_1405 ? (_GEN_4945 ? ~_GEN_365 & _GEN_4943 : ~(_GEN_1403 & _GEN_365) & _GEN_4943) : _GEN_4943;
  wire        _GEN_4977 = _GEN_1405 ? (_GEN_4945 ? ~(&lcam_ldq_idx_1) & _GEN_4944 : ~(_GEN_1403 & (&lcam_ldq_idx_1)) & _GEN_4944) : _GEN_4944;
  wire        _GEN_4978 = _GEN_1412 | _GEN_1413;
  wire        _GEN_4979 = _GEN_1410 ? (_GEN_4978 ? (|lcam_ldq_idx_0) & _GEN_4946 : ~(_GEN_1414 & ~(|lcam_ldq_idx_0)) & _GEN_4946) : _GEN_4946;
  wire        _GEN_4980 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_296 & _GEN_4947 : ~(_GEN_1414 & _GEN_296) & _GEN_4947) : _GEN_4947;
  wire        _GEN_4981 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_297 & _GEN_4948 : ~(_GEN_1414 & _GEN_297) & _GEN_4948) : _GEN_4948;
  wire        _GEN_4982 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_298 & _GEN_4949 : ~(_GEN_1414 & _GEN_298) & _GEN_4949) : _GEN_4949;
  wire        _GEN_4983 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_299 & _GEN_4950 : ~(_GEN_1414 & _GEN_299) & _GEN_4950) : _GEN_4950;
  wire        _GEN_4984 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_300 & _GEN_4951 : ~(_GEN_1414 & _GEN_300) & _GEN_4951) : _GEN_4951;
  wire        _GEN_4985 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_301 & _GEN_4952 : ~(_GEN_1414 & _GEN_301) & _GEN_4952) : _GEN_4952;
  wire        _GEN_4986 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_302 & _GEN_4953 : ~(_GEN_1414 & _GEN_302) & _GEN_4953) : _GEN_4953;
  wire        _GEN_4987 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_303 & _GEN_4954 : ~(_GEN_1414 & _GEN_303) & _GEN_4954) : _GEN_4954;
  wire        _GEN_4988 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_304 & _GEN_4955 : ~(_GEN_1414 & _GEN_304) & _GEN_4955) : _GEN_4955;
  wire        _GEN_4989 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_305 & _GEN_4956 : ~(_GEN_1414 & _GEN_305) & _GEN_4956) : _GEN_4956;
  wire        _GEN_4990 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_306 & _GEN_4957 : ~(_GEN_1414 & _GEN_306) & _GEN_4957) : _GEN_4957;
  wire        _GEN_4991 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_307 & _GEN_4958 : ~(_GEN_1414 & _GEN_307) & _GEN_4958) : _GEN_4958;
  wire        _GEN_4992 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_308 & _GEN_4959 : ~(_GEN_1414 & _GEN_308) & _GEN_4959) : _GEN_4959;
  wire        _GEN_4993 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_309 & _GEN_4960 : ~(_GEN_1414 & _GEN_309) & _GEN_4960) : _GEN_4960;
  wire        _GEN_4994 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_310 & _GEN_4961 : ~(_GEN_1414 & _GEN_310) & _GEN_4961) : _GEN_4961;
  wire        _GEN_4995 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_311 & _GEN_4962 : ~(_GEN_1414 & _GEN_311) & _GEN_4962) : _GEN_4962;
  wire        _GEN_4996 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_312 & _GEN_4963 : ~(_GEN_1414 & _GEN_312) & _GEN_4963) : _GEN_4963;
  wire        _GEN_4997 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_313 & _GEN_4964 : ~(_GEN_1414 & _GEN_313) & _GEN_4964) : _GEN_4964;
  wire        _GEN_4998 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_314 & _GEN_4965 : ~(_GEN_1414 & _GEN_314) & _GEN_4965) : _GEN_4965;
  wire        _GEN_4999 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_315 & _GEN_4966 : ~(_GEN_1414 & _GEN_315) & _GEN_4966) : _GEN_4966;
  wire        _GEN_5000 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_316 & _GEN_4967 : ~(_GEN_1414 & _GEN_316) & _GEN_4967) : _GEN_4967;
  wire        _GEN_5001 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_317 & _GEN_4968 : ~(_GEN_1414 & _GEN_317) & _GEN_4968) : _GEN_4968;
  wire        _GEN_5002 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_318 & _GEN_4969 : ~(_GEN_1414 & _GEN_318) & _GEN_4969) : _GEN_4969;
  wire        _GEN_5003 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_319 & _GEN_4970 : ~(_GEN_1414 & _GEN_319) & _GEN_4970) : _GEN_4970;
  wire        _GEN_5004 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_320 & _GEN_4971 : ~(_GEN_1414 & _GEN_320) & _GEN_4971) : _GEN_4971;
  wire        _GEN_5005 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_321 & _GEN_4972 : ~(_GEN_1414 & _GEN_321) & _GEN_4972) : _GEN_4972;
  wire        _GEN_5006 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_322 & _GEN_4973 : ~(_GEN_1414 & _GEN_322) & _GEN_4973) : _GEN_4973;
  wire        _GEN_5007 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_323 & _GEN_4974 : ~(_GEN_1414 & _GEN_323) & _GEN_4974) : _GEN_4974;
  wire        _GEN_5008 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_324 & _GEN_4975 : ~(_GEN_1414 & _GEN_324) & _GEN_4975) : _GEN_4975;
  wire        _GEN_5009 = _GEN_1410 ? (_GEN_4978 ? ~_GEN_325 & _GEN_4976 : ~(_GEN_1414 & _GEN_325) & _GEN_4976) : _GEN_4976;
  wire        _GEN_5010 = _GEN_1410 ? (_GEN_4978 ? ~(&lcam_ldq_idx_0) & _GEN_4977 : ~(_GEN_1414 & (&lcam_ldq_idx_0)) & _GEN_4977) : _GEN_4977;
  wire        _GEN_5011 = _GEN_1418 | _GEN_1419;
  wire        _GEN_5012 = _GEN_1416 ? (_GEN_5011 ? (|lcam_ldq_idx_1) & _GEN_4979 : ~(_GEN_1414 & ~(|lcam_ldq_idx_1)) & _GEN_4979) : _GEN_4979;
  wire        _GEN_5013 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_336 & _GEN_4980 : ~(_GEN_1414 & _GEN_336) & _GEN_4980) : _GEN_4980;
  wire        _GEN_5014 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_337 & _GEN_4981 : ~(_GEN_1414 & _GEN_337) & _GEN_4981) : _GEN_4981;
  wire        _GEN_5015 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_338 & _GEN_4982 : ~(_GEN_1414 & _GEN_338) & _GEN_4982) : _GEN_4982;
  wire        _GEN_5016 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_339 & _GEN_4983 : ~(_GEN_1414 & _GEN_339) & _GEN_4983) : _GEN_4983;
  wire        _GEN_5017 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_340 & _GEN_4984 : ~(_GEN_1414 & _GEN_340) & _GEN_4984) : _GEN_4984;
  wire        _GEN_5018 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_341 & _GEN_4985 : ~(_GEN_1414 & _GEN_341) & _GEN_4985) : _GEN_4985;
  wire        _GEN_5019 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_342 & _GEN_4986 : ~(_GEN_1414 & _GEN_342) & _GEN_4986) : _GEN_4986;
  wire        _GEN_5020 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_343 & _GEN_4987 : ~(_GEN_1414 & _GEN_343) & _GEN_4987) : _GEN_4987;
  wire        _GEN_5021 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_344 & _GEN_4988 : ~(_GEN_1414 & _GEN_344) & _GEN_4988) : _GEN_4988;
  wire        _GEN_5022 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_345 & _GEN_4989 : ~(_GEN_1414 & _GEN_345) & _GEN_4989) : _GEN_4989;
  wire        _GEN_5023 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_346 & _GEN_4990 : ~(_GEN_1414 & _GEN_346) & _GEN_4990) : _GEN_4990;
  wire        _GEN_5024 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_347 & _GEN_4991 : ~(_GEN_1414 & _GEN_347) & _GEN_4991) : _GEN_4991;
  wire        _GEN_5025 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_348 & _GEN_4992 : ~(_GEN_1414 & _GEN_348) & _GEN_4992) : _GEN_4992;
  wire        _GEN_5026 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_349 & _GEN_4993 : ~(_GEN_1414 & _GEN_349) & _GEN_4993) : _GEN_4993;
  wire        _GEN_5027 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_350 & _GEN_4994 : ~(_GEN_1414 & _GEN_350) & _GEN_4994) : _GEN_4994;
  wire        _GEN_5028 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_351 & _GEN_4995 : ~(_GEN_1414 & _GEN_351) & _GEN_4995) : _GEN_4995;
  wire        _GEN_5029 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_352 & _GEN_4996 : ~(_GEN_1414 & _GEN_352) & _GEN_4996) : _GEN_4996;
  wire        _GEN_5030 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_353 & _GEN_4997 : ~(_GEN_1414 & _GEN_353) & _GEN_4997) : _GEN_4997;
  wire        _GEN_5031 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_354 & _GEN_4998 : ~(_GEN_1414 & _GEN_354) & _GEN_4998) : _GEN_4998;
  wire        _GEN_5032 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_355 & _GEN_4999 : ~(_GEN_1414 & _GEN_355) & _GEN_4999) : _GEN_4999;
  wire        _GEN_5033 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_356 & _GEN_5000 : ~(_GEN_1414 & _GEN_356) & _GEN_5000) : _GEN_5000;
  wire        _GEN_5034 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_357 & _GEN_5001 : ~(_GEN_1414 & _GEN_357) & _GEN_5001) : _GEN_5001;
  wire        _GEN_5035 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_358 & _GEN_5002 : ~(_GEN_1414 & _GEN_358) & _GEN_5002) : _GEN_5002;
  wire        _GEN_5036 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_359 & _GEN_5003 : ~(_GEN_1414 & _GEN_359) & _GEN_5003) : _GEN_5003;
  wire        _GEN_5037 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_360 & _GEN_5004 : ~(_GEN_1414 & _GEN_360) & _GEN_5004) : _GEN_5004;
  wire        _GEN_5038 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_361 & _GEN_5005 : ~(_GEN_1414 & _GEN_361) & _GEN_5005) : _GEN_5005;
  wire        _GEN_5039 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_362 & _GEN_5006 : ~(_GEN_1414 & _GEN_362) & _GEN_5006) : _GEN_5006;
  wire        _GEN_5040 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_363 & _GEN_5007 : ~(_GEN_1414 & _GEN_363) & _GEN_5007) : _GEN_5007;
  wire        _GEN_5041 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_364 & _GEN_5008 : ~(_GEN_1414 & _GEN_364) & _GEN_5008) : _GEN_5008;
  wire        _GEN_5042 = _GEN_1416 ? (_GEN_5011 ? ~_GEN_365 & _GEN_5009 : ~(_GEN_1414 & _GEN_365) & _GEN_5009) : _GEN_5009;
  wire        _GEN_5043 = _GEN_1416 ? (_GEN_5011 ? ~(&lcam_ldq_idx_1) & _GEN_5010 : ~(_GEN_1414 & (&lcam_ldq_idx_1)) & _GEN_5010) : _GEN_5010;
  wire        _GEN_5044 = _GEN_1423 | _GEN_1424;
  wire        _GEN_5045 = _GEN_1421 ? (_GEN_5044 ? (|lcam_ldq_idx_0) & _GEN_5012 : ~(_GEN_1425 & ~(|lcam_ldq_idx_0)) & _GEN_5012) : _GEN_5012;
  wire        _GEN_5046 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_296 & _GEN_5013 : ~(_GEN_1425 & _GEN_296) & _GEN_5013) : _GEN_5013;
  wire        _GEN_5047 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_297 & _GEN_5014 : ~(_GEN_1425 & _GEN_297) & _GEN_5014) : _GEN_5014;
  wire        _GEN_5048 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_298 & _GEN_5015 : ~(_GEN_1425 & _GEN_298) & _GEN_5015) : _GEN_5015;
  wire        _GEN_5049 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_299 & _GEN_5016 : ~(_GEN_1425 & _GEN_299) & _GEN_5016) : _GEN_5016;
  wire        _GEN_5050 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_300 & _GEN_5017 : ~(_GEN_1425 & _GEN_300) & _GEN_5017) : _GEN_5017;
  wire        _GEN_5051 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_301 & _GEN_5018 : ~(_GEN_1425 & _GEN_301) & _GEN_5018) : _GEN_5018;
  wire        _GEN_5052 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_302 & _GEN_5019 : ~(_GEN_1425 & _GEN_302) & _GEN_5019) : _GEN_5019;
  wire        _GEN_5053 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_303 & _GEN_5020 : ~(_GEN_1425 & _GEN_303) & _GEN_5020) : _GEN_5020;
  wire        _GEN_5054 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_304 & _GEN_5021 : ~(_GEN_1425 & _GEN_304) & _GEN_5021) : _GEN_5021;
  wire        _GEN_5055 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_305 & _GEN_5022 : ~(_GEN_1425 & _GEN_305) & _GEN_5022) : _GEN_5022;
  wire        _GEN_5056 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_306 & _GEN_5023 : ~(_GEN_1425 & _GEN_306) & _GEN_5023) : _GEN_5023;
  wire        _GEN_5057 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_307 & _GEN_5024 : ~(_GEN_1425 & _GEN_307) & _GEN_5024) : _GEN_5024;
  wire        _GEN_5058 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_308 & _GEN_5025 : ~(_GEN_1425 & _GEN_308) & _GEN_5025) : _GEN_5025;
  wire        _GEN_5059 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_309 & _GEN_5026 : ~(_GEN_1425 & _GEN_309) & _GEN_5026) : _GEN_5026;
  wire        _GEN_5060 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_310 & _GEN_5027 : ~(_GEN_1425 & _GEN_310) & _GEN_5027) : _GEN_5027;
  wire        _GEN_5061 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_311 & _GEN_5028 : ~(_GEN_1425 & _GEN_311) & _GEN_5028) : _GEN_5028;
  wire        _GEN_5062 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_312 & _GEN_5029 : ~(_GEN_1425 & _GEN_312) & _GEN_5029) : _GEN_5029;
  wire        _GEN_5063 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_313 & _GEN_5030 : ~(_GEN_1425 & _GEN_313) & _GEN_5030) : _GEN_5030;
  wire        _GEN_5064 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_314 & _GEN_5031 : ~(_GEN_1425 & _GEN_314) & _GEN_5031) : _GEN_5031;
  wire        _GEN_5065 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_315 & _GEN_5032 : ~(_GEN_1425 & _GEN_315) & _GEN_5032) : _GEN_5032;
  wire        _GEN_5066 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_316 & _GEN_5033 : ~(_GEN_1425 & _GEN_316) & _GEN_5033) : _GEN_5033;
  wire        _GEN_5067 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_317 & _GEN_5034 : ~(_GEN_1425 & _GEN_317) & _GEN_5034) : _GEN_5034;
  wire        _GEN_5068 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_318 & _GEN_5035 : ~(_GEN_1425 & _GEN_318) & _GEN_5035) : _GEN_5035;
  wire        _GEN_5069 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_319 & _GEN_5036 : ~(_GEN_1425 & _GEN_319) & _GEN_5036) : _GEN_5036;
  wire        _GEN_5070 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_320 & _GEN_5037 : ~(_GEN_1425 & _GEN_320) & _GEN_5037) : _GEN_5037;
  wire        _GEN_5071 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_321 & _GEN_5038 : ~(_GEN_1425 & _GEN_321) & _GEN_5038) : _GEN_5038;
  wire        _GEN_5072 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_322 & _GEN_5039 : ~(_GEN_1425 & _GEN_322) & _GEN_5039) : _GEN_5039;
  wire        _GEN_5073 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_323 & _GEN_5040 : ~(_GEN_1425 & _GEN_323) & _GEN_5040) : _GEN_5040;
  wire        _GEN_5074 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_324 & _GEN_5041 : ~(_GEN_1425 & _GEN_324) & _GEN_5041) : _GEN_5041;
  wire        _GEN_5075 = _GEN_1421 ? (_GEN_5044 ? ~_GEN_325 & _GEN_5042 : ~(_GEN_1425 & _GEN_325) & _GEN_5042) : _GEN_5042;
  wire        _GEN_5076 = _GEN_1421 ? (_GEN_5044 ? ~(&lcam_ldq_idx_0) & _GEN_5043 : ~(_GEN_1425 & (&lcam_ldq_idx_0)) & _GEN_5043) : _GEN_5043;
  wire        _GEN_5077 = _GEN_1428 | _GEN_1429;
  wire        ld_xcpt_valid = _temp_bits_WIRE_1_32 | _temp_bits_WIRE_1_33 | _temp_bits_WIRE_1_34 | _temp_bits_WIRE_1_35 | _temp_bits_WIRE_1_36 | _temp_bits_WIRE_1_37 | _temp_bits_WIRE_1_38 | _temp_bits_WIRE_1_39 | _temp_bits_WIRE_1_40 | _temp_bits_WIRE_1_41 | _temp_bits_WIRE_1_42 | _temp_bits_WIRE_1_43 | _temp_bits_WIRE_1_44 | _temp_bits_WIRE_1_45 | _temp_bits_WIRE_1_46 | _temp_bits_WIRE_1_47 | _temp_bits_WIRE_1_48 | _temp_bits_WIRE_1_49 | _temp_bits_WIRE_1_50 | _temp_bits_WIRE_1_51 | _temp_bits_WIRE_1_52 | _temp_bits_WIRE_1_53 | _temp_bits_WIRE_1_54 | _temp_bits_WIRE_1_55 | _temp_bits_WIRE_1_56 | _temp_bits_WIRE_1_57 | _temp_bits_WIRE_1_58 | _temp_bits_WIRE_1_59 | _temp_bits_WIRE_1_60 | _temp_bits_WIRE_1_61 | _temp_bits_WIRE_1_62 | _temp_bits_WIRE_1_63;
  wire        use_mem_xcpt = mem_xcpt_valid & (mem_xcpt_uop_rob_idx < casez_tmp_458 ^ mem_xcpt_uop_rob_idx < io_core_rob_head_idx ^ casez_tmp_458 < io_core_rob_head_idx) | ~ld_xcpt_valid;
  wire [19:0] xcpt_uop_br_mask = use_mem_xcpt ? (_GEN_2550 ? mem_xcpt_uops_1_br_mask : mem_xcpt_uops_0_br_mask) : casez_tmp_457;
  wire        _ldq_bits_succeeded_T = _io_core_exe_0_iresp_valid_output | _io_core_exe_0_fresp_valid_output;
  wire        _GEN_5078 = casez_tmp_490 & live;
  wire        _GEN_5079 = _GEN_1469 & _GEN_5078 & ~(|wb_forward_ldq_idx_0);
  wire        _GEN_5080 = _GEN_1468 | ~_GEN_5079;
  wire        _GEN_5081 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h1;
  wire        _GEN_5082 = _GEN_1468 | ~_GEN_5081;
  wire        _GEN_5083 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h2;
  wire        _GEN_5084 = _GEN_1468 | ~_GEN_5083;
  wire        _GEN_5085 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h3;
  wire        _GEN_5086 = _GEN_1468 | ~_GEN_5085;
  wire        _GEN_5087 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h4;
  wire        _GEN_5088 = _GEN_1468 | ~_GEN_5087;
  wire        _GEN_5089 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h5;
  wire        _GEN_5090 = _GEN_1468 | ~_GEN_5089;
  wire        _GEN_5091 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h6;
  wire        _GEN_5092 = _GEN_1468 | ~_GEN_5091;
  wire        _GEN_5093 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h7;
  wire        _GEN_5094 = _GEN_1468 | ~_GEN_5093;
  wire        _GEN_5095 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h8;
  wire        _GEN_5096 = _GEN_1468 | ~_GEN_5095;
  wire        _GEN_5097 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h9;
  wire        _GEN_5098 = _GEN_1468 | ~_GEN_5097;
  wire        _GEN_5099 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'hA;
  wire        _GEN_5100 = _GEN_1468 | ~_GEN_5099;
  wire        _GEN_5101 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'hB;
  wire        _GEN_5102 = _GEN_1468 | ~_GEN_5101;
  wire        _GEN_5103 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'hC;
  wire        _GEN_5104 = _GEN_1468 | ~_GEN_5103;
  wire        _GEN_5105 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'hD;
  wire        _GEN_5106 = _GEN_1468 | ~_GEN_5105;
  wire        _GEN_5107 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'hE;
  wire        _GEN_5108 = _GEN_1468 | ~_GEN_5107;
  wire        _GEN_5109 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'hF;
  wire        _GEN_5110 = _GEN_1468 | ~_GEN_5109;
  wire        _GEN_5111 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h10;
  wire        _GEN_5112 = _GEN_1468 | ~_GEN_5111;
  wire        _GEN_5113 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h11;
  wire        _GEN_5114 = _GEN_1468 | ~_GEN_5113;
  wire        _GEN_5115 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h12;
  wire        _GEN_5116 = _GEN_1468 | ~_GEN_5115;
  wire        _GEN_5117 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h13;
  wire        _GEN_5118 = _GEN_1468 | ~_GEN_5117;
  wire        _GEN_5119 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h14;
  wire        _GEN_5120 = _GEN_1468 | ~_GEN_5119;
  wire        _GEN_5121 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h15;
  wire        _GEN_5122 = _GEN_1468 | ~_GEN_5121;
  wire        _GEN_5123 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h16;
  wire        _GEN_5124 = _GEN_1468 | ~_GEN_5123;
  wire        _GEN_5125 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h17;
  wire        _GEN_5126 = _GEN_1468 | ~_GEN_5125;
  wire        _GEN_5127 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h18;
  wire        _GEN_5128 = _GEN_1468 | ~_GEN_5127;
  wire        _GEN_5129 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h19;
  wire        _GEN_5130 = _GEN_1468 | ~_GEN_5129;
  wire        _GEN_5131 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h1A;
  wire        _GEN_5132 = _GEN_1468 | ~_GEN_5131;
  wire        _GEN_5133 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h1B;
  wire        _GEN_5134 = _GEN_1468 | ~_GEN_5133;
  wire        _GEN_5135 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h1C;
  wire        _GEN_5136 = _GEN_1468 | ~_GEN_5135;
  wire        _GEN_5137 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h1D;
  wire        _GEN_5138 = _GEN_1468 | ~_GEN_5137;
  wire        _GEN_5139 = _GEN_1469 & _GEN_5078 & wb_forward_ldq_idx_0 == 5'h1E;
  wire        _GEN_5140 = _GEN_1468 | ~_GEN_5139;
  wire        _GEN_5141 = _GEN_1469 & _GEN_5078 & (&wb_forward_ldq_idx_0);
  wire        _GEN_5142 = _GEN_1468 | ~_GEN_5141;
  wire        _ldq_bits_succeeded_T_1 = _io_core_exe_1_iresp_valid_output | _io_core_exe_1_fresp_valid_output;
  wire        _GEN_5143 = casez_tmp_524 & live_1;
  wire        _GEN_5144 = _GEN_1509 & _GEN_5143 & ~(|wb_forward_ldq_idx_1);
  wire        _GEN_5145 = _GEN_1508 | ~_GEN_5144;
  wire        _GEN_5146 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h1;
  wire        _GEN_5147 = _GEN_1508 | ~_GEN_5146;
  wire        _GEN_5148 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h2;
  wire        _GEN_5149 = _GEN_1508 | ~_GEN_5148;
  wire        _GEN_5150 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h3;
  wire        _GEN_5151 = _GEN_1508 | ~_GEN_5150;
  wire        _GEN_5152 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h4;
  wire        _GEN_5153 = _GEN_1508 | ~_GEN_5152;
  wire        _GEN_5154 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h5;
  wire        _GEN_5155 = _GEN_1508 | ~_GEN_5154;
  wire        _GEN_5156 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h6;
  wire        _GEN_5157 = _GEN_1508 | ~_GEN_5156;
  wire        _GEN_5158 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h7;
  wire        _GEN_5159 = _GEN_1508 | ~_GEN_5158;
  wire        _GEN_5160 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h8;
  wire        _GEN_5161 = _GEN_1508 | ~_GEN_5160;
  wire        _GEN_5162 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h9;
  wire        _GEN_5163 = _GEN_1508 | ~_GEN_5162;
  wire        _GEN_5164 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'hA;
  wire        _GEN_5165 = _GEN_1508 | ~_GEN_5164;
  wire        _GEN_5166 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'hB;
  wire        _GEN_5167 = _GEN_1508 | ~_GEN_5166;
  wire        _GEN_5168 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'hC;
  wire        _GEN_5169 = _GEN_1508 | ~_GEN_5168;
  wire        _GEN_5170 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'hD;
  wire        _GEN_5171 = _GEN_1508 | ~_GEN_5170;
  wire        _GEN_5172 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'hE;
  wire        _GEN_5173 = _GEN_1508 | ~_GEN_5172;
  wire        _GEN_5174 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'hF;
  wire        _GEN_5175 = _GEN_1508 | ~_GEN_5174;
  wire        _GEN_5176 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h10;
  wire        _GEN_5177 = _GEN_1508 | ~_GEN_5176;
  wire        _GEN_5178 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h11;
  wire        _GEN_5179 = _GEN_1508 | ~_GEN_5178;
  wire        _GEN_5180 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h12;
  wire        _GEN_5181 = _GEN_1508 | ~_GEN_5180;
  wire        _GEN_5182 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h13;
  wire        _GEN_5183 = _GEN_1508 | ~_GEN_5182;
  wire        _GEN_5184 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h14;
  wire        _GEN_5185 = _GEN_1508 | ~_GEN_5184;
  wire        _GEN_5186 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h15;
  wire        _GEN_5187 = _GEN_1508 | ~_GEN_5186;
  wire        _GEN_5188 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h16;
  wire        _GEN_5189 = _GEN_1508 | ~_GEN_5188;
  wire        _GEN_5190 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h17;
  wire        _GEN_5191 = _GEN_1508 | ~_GEN_5190;
  wire        _GEN_5192 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h18;
  wire        _GEN_5193 = _GEN_1508 | ~_GEN_5192;
  wire        _GEN_5194 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h19;
  wire        _GEN_5195 = _GEN_1508 | ~_GEN_5194;
  wire        _GEN_5196 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h1A;
  wire        _GEN_5197 = _GEN_1508 | ~_GEN_5196;
  wire        _GEN_5198 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h1B;
  wire        _GEN_5199 = _GEN_1508 | ~_GEN_5198;
  wire        _GEN_5200 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h1C;
  wire        _GEN_5201 = _GEN_1508 | ~_GEN_5200;
  wire        _GEN_5202 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h1D;
  wire        _GEN_5203 = _GEN_1508 | ~_GEN_5202;
  wire        _GEN_5204 = _GEN_1509 & _GEN_5143 & wb_forward_ldq_idx_1 == 5'h1E;
  wire        _GEN_5205 = _GEN_1508 | ~_GEN_5204;
  wire        _GEN_5206 = _GEN_1509 & _GEN_5143 & (&wb_forward_ldq_idx_1);
  wire        _GEN_5207 = _GEN_1508 | ~_GEN_5206;
  wire        _GEN_5208 = stq_0_valid & (|_GEN_1511);
  wire        _GEN_5209 = stq_1_valid & (|_GEN_1512);
  wire        _GEN_5210 = stq_2_valid & (|_GEN_1513);
  wire        _GEN_5211 = stq_3_valid & (|_GEN_1514);
  wire        _GEN_5212 = stq_4_valid & (|_GEN_1515);
  wire        _GEN_5213 = stq_5_valid & (|_GEN_1516);
  wire        _GEN_5214 = stq_6_valid & (|_GEN_1517);
  wire        _GEN_5215 = stq_7_valid & (|_GEN_1518);
  wire        _GEN_5216 = stq_8_valid & (|_GEN_1519);
  wire        _GEN_5217 = stq_9_valid & (|_GEN_1520);
  wire        _GEN_5218 = stq_10_valid & (|_GEN_1521);
  wire        _GEN_5219 = stq_11_valid & (|_GEN_1522);
  wire        _GEN_5220 = stq_12_valid & (|_GEN_1523);
  wire        _GEN_5221 = stq_13_valid & (|_GEN_1524);
  wire        _GEN_5222 = stq_14_valid & (|_GEN_1525);
  wire        _GEN_5223 = stq_15_valid & (|_GEN_1526);
  wire        _GEN_5224 = stq_16_valid & (|_GEN_1527);
  wire        _GEN_5225 = stq_17_valid & (|_GEN_1528);
  wire        _GEN_5226 = stq_18_valid & (|_GEN_1529);
  wire        _GEN_5227 = stq_19_valid & (|_GEN_1530);
  wire        _GEN_5228 = stq_20_valid & (|_GEN_1531);
  wire        _GEN_5229 = stq_21_valid & (|_GEN_1532);
  wire        _GEN_5230 = stq_22_valid & (|_GEN_1533);
  wire        _GEN_5231 = stq_23_valid & (|_GEN_1534);
  wire        _GEN_5232 = stq_24_valid & (|_GEN_1535);
  wire        _GEN_5233 = stq_25_valid & (|_GEN_1536);
  wire        _GEN_5234 = stq_26_valid & (|_GEN_1537);
  wire        _GEN_5235 = stq_27_valid & (|_GEN_1538);
  wire        _GEN_5236 = stq_28_valid & (|_GEN_1539);
  wire        _GEN_5237 = stq_29_valid & (|_GEN_1540);
  wire        _GEN_5238 = stq_30_valid & (|_GEN_1541);
  wire        _GEN_5239 = stq_31_valid & (|_GEN_1542);
  wire        _GEN_5240 = ldq_0_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_0_bits_uop_br_mask));
  wire        _GEN_5241 = ldq_1_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_1_bits_uop_br_mask));
  wire        _GEN_5242 = ldq_2_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_2_bits_uop_br_mask));
  wire        _GEN_5243 = ldq_3_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_3_bits_uop_br_mask));
  wire        _GEN_5244 = ldq_4_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_4_bits_uop_br_mask));
  wire        _GEN_5245 = ldq_5_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_5_bits_uop_br_mask));
  wire        _GEN_5246 = ldq_6_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_6_bits_uop_br_mask));
  wire        _GEN_5247 = ldq_7_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_7_bits_uop_br_mask));
  wire        _GEN_5248 = ldq_8_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_8_bits_uop_br_mask));
  wire        _GEN_5249 = ldq_9_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_9_bits_uop_br_mask));
  wire        _GEN_5250 = ldq_10_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_10_bits_uop_br_mask));
  wire        _GEN_5251 = ldq_11_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_11_bits_uop_br_mask));
  wire        _GEN_5252 = ldq_12_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_12_bits_uop_br_mask));
  wire        _GEN_5253 = ldq_13_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_13_bits_uop_br_mask));
  wire        _GEN_5254 = ldq_14_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_14_bits_uop_br_mask));
  wire        _GEN_5255 = ldq_15_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_15_bits_uop_br_mask));
  wire        _GEN_5256 = ldq_16_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_16_bits_uop_br_mask));
  wire        _GEN_5257 = ldq_17_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_17_bits_uop_br_mask));
  wire        _GEN_5258 = ldq_18_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_18_bits_uop_br_mask));
  wire        _GEN_5259 = ldq_19_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_19_bits_uop_br_mask));
  wire        _GEN_5260 = ldq_20_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_20_bits_uop_br_mask));
  wire        _GEN_5261 = ldq_21_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_21_bits_uop_br_mask));
  wire        _GEN_5262 = ldq_22_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_22_bits_uop_br_mask));
  wire        _GEN_5263 = ldq_23_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_23_bits_uop_br_mask));
  wire        _GEN_5264 = ldq_24_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_24_bits_uop_br_mask));
  wire        _GEN_5265 = ldq_25_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_25_bits_uop_br_mask));
  wire        _GEN_5266 = ldq_26_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_26_bits_uop_br_mask));
  wire        _GEN_5267 = ldq_27_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_27_bits_uop_br_mask));
  wire        _GEN_5268 = ldq_28_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_28_bits_uop_br_mask));
  wire        _GEN_5269 = ldq_29_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_29_bits_uop_br_mask));
  wire        _GEN_5270 = ldq_30_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_30_bits_uop_br_mask));
  wire        _GEN_5271 = ldq_31_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_31_bits_uop_br_mask));
  wire        _GEN_5272 = idx == 5'h0;
  wire        _GEN_5273 = commit_store & _GEN_5272;
  wire        _GEN_5274 = idx == 5'h1;
  wire        _GEN_5275 = commit_store & _GEN_5274;
  wire        _GEN_5276 = idx == 5'h2;
  wire        _GEN_5277 = commit_store & _GEN_5276;
  wire        _GEN_5278 = idx == 5'h3;
  wire        _GEN_5279 = commit_store & _GEN_5278;
  wire        _GEN_5280 = idx == 5'h4;
  wire        _GEN_5281 = commit_store & _GEN_5280;
  wire        _GEN_5282 = idx == 5'h5;
  wire        _GEN_5283 = commit_store & _GEN_5282;
  wire        _GEN_5284 = idx == 5'h6;
  wire        _GEN_5285 = commit_store & _GEN_5284;
  wire        _GEN_5286 = idx == 5'h7;
  wire        _GEN_5287 = commit_store & _GEN_5286;
  wire        _GEN_5288 = idx == 5'h8;
  wire        _GEN_5289 = commit_store & _GEN_5288;
  wire        _GEN_5290 = idx == 5'h9;
  wire        _GEN_5291 = commit_store & _GEN_5290;
  wire        _GEN_5292 = idx == 5'hA;
  wire        _GEN_5293 = commit_store & _GEN_5292;
  wire        _GEN_5294 = idx == 5'hB;
  wire        _GEN_5295 = commit_store & _GEN_5294;
  wire        _GEN_5296 = idx == 5'hC;
  wire        _GEN_5297 = commit_store & _GEN_5296;
  wire        _GEN_5298 = idx == 5'hD;
  wire        _GEN_5299 = commit_store & _GEN_5298;
  wire        _GEN_5300 = idx == 5'hE;
  wire        _GEN_5301 = commit_store & _GEN_5300;
  wire        _GEN_5302 = idx == 5'hF;
  wire        _GEN_5303 = commit_store & _GEN_5302;
  wire        _GEN_5304 = idx == 5'h10;
  wire        _GEN_5305 = commit_store & _GEN_5304;
  wire        _GEN_5306 = idx == 5'h11;
  wire        _GEN_5307 = commit_store & _GEN_5306;
  wire        _GEN_5308 = idx == 5'h12;
  wire        _GEN_5309 = commit_store & _GEN_5308;
  wire        _GEN_5310 = idx == 5'h13;
  wire        _GEN_5311 = commit_store & _GEN_5310;
  wire        _GEN_5312 = idx == 5'h14;
  wire        _GEN_5313 = commit_store & _GEN_5312;
  wire        _GEN_5314 = idx == 5'h15;
  wire        _GEN_5315 = commit_store & _GEN_5314;
  wire        _GEN_5316 = idx == 5'h16;
  wire        _GEN_5317 = commit_store & _GEN_5316;
  wire        _GEN_5318 = idx == 5'h17;
  wire        _GEN_5319 = commit_store & _GEN_5318;
  wire        _GEN_5320 = idx == 5'h18;
  wire        _GEN_5321 = commit_store & _GEN_5320;
  wire        _GEN_5322 = idx == 5'h19;
  wire        _GEN_5323 = commit_store & _GEN_5322;
  wire        _GEN_5324 = idx == 5'h1A;
  wire        _GEN_5325 = commit_store & _GEN_5324;
  wire        _GEN_5326 = idx == 5'h1B;
  wire        _GEN_5327 = commit_store & _GEN_5326;
  wire        _GEN_5328 = idx == 5'h1C;
  wire        _GEN_5329 = commit_store & _GEN_5328;
  wire        _GEN_5330 = idx == 5'h1D;
  wire        _GEN_5331 = commit_store & _GEN_5330;
  wire        _GEN_5332 = idx == 5'h1E;
  wire        _GEN_5333 = commit_store & _GEN_5332;
  wire        _GEN_5334 = commit_store & (&idx);
  wire        _GEN_5335 = _GEN_5272 | _GEN_5240;
  wire        _GEN_5336 = commit_store | ~commit_load;
  wire        _GEN_5337 = _GEN_5274 | _GEN_5241;
  wire        _GEN_5338 = _GEN_5276 | _GEN_5242;
  wire        _GEN_5339 = _GEN_5278 | _GEN_5243;
  wire        _GEN_5340 = _GEN_5280 | _GEN_5244;
  wire        _GEN_5341 = _GEN_5282 | _GEN_5245;
  wire        _GEN_5342 = _GEN_5284 | _GEN_5246;
  wire        _GEN_5343 = _GEN_5286 | _GEN_5247;
  wire        _GEN_5344 = _GEN_5288 | _GEN_5248;
  wire        _GEN_5345 = _GEN_5290 | _GEN_5249;
  wire        _GEN_5346 = _GEN_5292 | _GEN_5250;
  wire        _GEN_5347 = _GEN_5294 | _GEN_5251;
  wire        _GEN_5348 = _GEN_5296 | _GEN_5252;
  wire        _GEN_5349 = _GEN_5298 | _GEN_5253;
  wire        _GEN_5350 = _GEN_5300 | _GEN_5254;
  wire        _GEN_5351 = _GEN_5302 | _GEN_5255;
  wire        _GEN_5352 = _GEN_5304 | _GEN_5256;
  wire        _GEN_5353 = _GEN_5306 | _GEN_5257;
  wire        _GEN_5354 = _GEN_5308 | _GEN_5258;
  wire        _GEN_5355 = _GEN_5310 | _GEN_5259;
  wire        _GEN_5356 = _GEN_5312 | _GEN_5260;
  wire        _GEN_5357 = _GEN_5314 | _GEN_5261;
  wire        _GEN_5358 = _GEN_5316 | _GEN_5262;
  wire        _GEN_5359 = _GEN_5318 | _GEN_5263;
  wire        _GEN_5360 = _GEN_5320 | _GEN_5264;
  wire        _GEN_5361 = _GEN_5322 | _GEN_5265;
  wire        _GEN_5362 = _GEN_5324 | _GEN_5266;
  wire        _GEN_5363 = _GEN_5326 | _GEN_5267;
  wire        _GEN_5364 = _GEN_5328 | _GEN_5268;
  wire        _GEN_5365 = _GEN_5330 | _GEN_5269;
  wire        _GEN_5366 = _GEN_5332 | _GEN_5270;
  wire        _GEN_5367 = (&idx) | _GEN_5271;
  wire        _GEN_5368 = commit_store | ~(commit_load & _GEN_5272);
  wire        _GEN_5369 = commit_store | ~(commit_load & _GEN_5274);
  wire        _GEN_5370 = commit_store | ~(commit_load & _GEN_5276);
  wire        _GEN_5371 = commit_store | ~(commit_load & _GEN_5278);
  wire        _GEN_5372 = commit_store | ~(commit_load & _GEN_5280);
  wire        _GEN_5373 = commit_store | ~(commit_load & _GEN_5282);
  wire        _GEN_5374 = commit_store | ~(commit_load & _GEN_5284);
  wire        _GEN_5375 = commit_store | ~(commit_load & _GEN_5286);
  wire        _GEN_5376 = commit_store | ~(commit_load & _GEN_5288);
  wire        _GEN_5377 = commit_store | ~(commit_load & _GEN_5290);
  wire        _GEN_5378 = commit_store | ~(commit_load & _GEN_5292);
  wire        _GEN_5379 = commit_store | ~(commit_load & _GEN_5294);
  wire        _GEN_5380 = commit_store | ~(commit_load & _GEN_5296);
  wire        _GEN_5381 = commit_store | ~(commit_load & _GEN_5298);
  wire        _GEN_5382 = commit_store | ~(commit_load & _GEN_5300);
  wire        _GEN_5383 = commit_store | ~(commit_load & _GEN_5302);
  wire        _GEN_5384 = commit_store | ~(commit_load & _GEN_5304);
  wire        _GEN_5385 = commit_store | ~(commit_load & _GEN_5306);
  wire        _GEN_5386 = commit_store | ~(commit_load & _GEN_5308);
  wire        _GEN_5387 = commit_store | ~(commit_load & _GEN_5310);
  wire        _GEN_5388 = commit_store | ~(commit_load & _GEN_5312);
  wire        _GEN_5389 = commit_store | ~(commit_load & _GEN_5314);
  wire        _GEN_5390 = commit_store | ~(commit_load & _GEN_5316);
  wire        _GEN_5391 = commit_store | ~(commit_load & _GEN_5318);
  wire        _GEN_5392 = commit_store | ~(commit_load & _GEN_5320);
  wire        _GEN_5393 = commit_store | ~(commit_load & _GEN_5322);
  wire        _GEN_5394 = commit_store | ~(commit_load & _GEN_5324);
  wire        _GEN_5395 = commit_store | ~(commit_load & _GEN_5326);
  wire        _GEN_5396 = commit_store | ~(commit_load & _GEN_5328);
  wire        _GEN_5397 = commit_store | ~(commit_load & _GEN_5330);
  wire        _GEN_5398 = commit_store | ~(commit_load & _GEN_5332);
  wire        _GEN_5399 = commit_store | ~(commit_load & (&idx));
  wire        _GEN_5400 = idx_1 == 5'h0;
  wire        _GEN_5401 = commit_store_1 ? _GEN_5400 | _GEN_5273 | _GEN_2518 : _GEN_5273 | _GEN_2518;
  wire        _GEN_5402 = idx_1 == 5'h1;
  wire        _GEN_5403 = commit_store_1 ? _GEN_5402 | _GEN_5275 | _GEN_2519 : _GEN_5275 | _GEN_2519;
  wire        _GEN_5404 = idx_1 == 5'h2;
  wire        _GEN_5405 = commit_store_1 ? _GEN_5404 | _GEN_5277 | _GEN_2520 : _GEN_5277 | _GEN_2520;
  wire        _GEN_5406 = idx_1 == 5'h3;
  wire        _GEN_5407 = commit_store_1 ? _GEN_5406 | _GEN_5279 | _GEN_2521 : _GEN_5279 | _GEN_2521;
  wire        _GEN_5408 = idx_1 == 5'h4;
  wire        _GEN_5409 = commit_store_1 ? _GEN_5408 | _GEN_5281 | _GEN_2522 : _GEN_5281 | _GEN_2522;
  wire        _GEN_5410 = idx_1 == 5'h5;
  wire        _GEN_5411 = commit_store_1 ? _GEN_5410 | _GEN_5283 | _GEN_2523 : _GEN_5283 | _GEN_2523;
  wire        _GEN_5412 = idx_1 == 5'h6;
  wire        _GEN_5413 = commit_store_1 ? _GEN_5412 | _GEN_5285 | _GEN_2524 : _GEN_5285 | _GEN_2524;
  wire        _GEN_5414 = idx_1 == 5'h7;
  wire        _GEN_5415 = commit_store_1 ? _GEN_5414 | _GEN_5287 | _GEN_2525 : _GEN_5287 | _GEN_2525;
  wire        _GEN_5416 = idx_1 == 5'h8;
  wire        _GEN_5417 = commit_store_1 ? _GEN_5416 | _GEN_5289 | _GEN_2526 : _GEN_5289 | _GEN_2526;
  wire        _GEN_5418 = idx_1 == 5'h9;
  wire        _GEN_5419 = commit_store_1 ? _GEN_5418 | _GEN_5291 | _GEN_2527 : _GEN_5291 | _GEN_2527;
  wire        _GEN_5420 = idx_1 == 5'hA;
  wire        _GEN_5421 = commit_store_1 ? _GEN_5420 | _GEN_5293 | _GEN_2528 : _GEN_5293 | _GEN_2528;
  wire        _GEN_5422 = idx_1 == 5'hB;
  wire        _GEN_5423 = commit_store_1 ? _GEN_5422 | _GEN_5295 | _GEN_2529 : _GEN_5295 | _GEN_2529;
  wire        _GEN_5424 = idx_1 == 5'hC;
  wire        _GEN_5425 = commit_store_1 ? _GEN_5424 | _GEN_5297 | _GEN_2530 : _GEN_5297 | _GEN_2530;
  wire        _GEN_5426 = idx_1 == 5'hD;
  wire        _GEN_5427 = commit_store_1 ? _GEN_5426 | _GEN_5299 | _GEN_2531 : _GEN_5299 | _GEN_2531;
  wire        _GEN_5428 = idx_1 == 5'hE;
  wire        _GEN_5429 = commit_store_1 ? _GEN_5428 | _GEN_5301 | _GEN_2532 : _GEN_5301 | _GEN_2532;
  wire        _GEN_5430 = idx_1 == 5'hF;
  wire        _GEN_5431 = commit_store_1 ? _GEN_5430 | _GEN_5303 | _GEN_2533 : _GEN_5303 | _GEN_2533;
  wire        _GEN_5432 = idx_1 == 5'h10;
  wire        _GEN_5433 = commit_store_1 ? _GEN_5432 | _GEN_5305 | _GEN_2534 : _GEN_5305 | _GEN_2534;
  wire        _GEN_5434 = idx_1 == 5'h11;
  wire        _GEN_5435 = commit_store_1 ? _GEN_5434 | _GEN_5307 | _GEN_2535 : _GEN_5307 | _GEN_2535;
  wire        _GEN_5436 = idx_1 == 5'h12;
  wire        _GEN_5437 = commit_store_1 ? _GEN_5436 | _GEN_5309 | _GEN_2536 : _GEN_5309 | _GEN_2536;
  wire        _GEN_5438 = idx_1 == 5'h13;
  wire        _GEN_5439 = commit_store_1 ? _GEN_5438 | _GEN_5311 | _GEN_2537 : _GEN_5311 | _GEN_2537;
  wire        _GEN_5440 = idx_1 == 5'h14;
  wire        _GEN_5441 = commit_store_1 ? _GEN_5440 | _GEN_5313 | _GEN_2538 : _GEN_5313 | _GEN_2538;
  wire        _GEN_5442 = idx_1 == 5'h15;
  wire        _GEN_5443 = commit_store_1 ? _GEN_5442 | _GEN_5315 | _GEN_2539 : _GEN_5315 | _GEN_2539;
  wire        _GEN_5444 = idx_1 == 5'h16;
  wire        _GEN_5445 = commit_store_1 ? _GEN_5444 | _GEN_5317 | _GEN_2540 : _GEN_5317 | _GEN_2540;
  wire        _GEN_5446 = idx_1 == 5'h17;
  wire        _GEN_5447 = commit_store_1 ? _GEN_5446 | _GEN_5319 | _GEN_2541 : _GEN_5319 | _GEN_2541;
  wire        _GEN_5448 = idx_1 == 5'h18;
  wire        _GEN_5449 = commit_store_1 ? _GEN_5448 | _GEN_5321 | _GEN_2542 : _GEN_5321 | _GEN_2542;
  wire        _GEN_5450 = idx_1 == 5'h19;
  wire        _GEN_5451 = commit_store_1 ? _GEN_5450 | _GEN_5323 | _GEN_2543 : _GEN_5323 | _GEN_2543;
  wire        _GEN_5452 = idx_1 == 5'h1A;
  wire        _GEN_5453 = commit_store_1 ? _GEN_5452 | _GEN_5325 | _GEN_2544 : _GEN_5325 | _GEN_2544;
  wire        _GEN_5454 = idx_1 == 5'h1B;
  wire        _GEN_5455 = commit_store_1 ? _GEN_5454 | _GEN_5327 | _GEN_2545 : _GEN_5327 | _GEN_2545;
  wire        _GEN_5456 = idx_1 == 5'h1C;
  wire        _GEN_5457 = commit_store_1 ? _GEN_5456 | _GEN_5329 | _GEN_2546 : _GEN_5329 | _GEN_2546;
  wire        _GEN_5458 = idx_1 == 5'h1D;
  wire        _GEN_5459 = commit_store_1 ? _GEN_5458 | _GEN_5331 | _GEN_2547 : _GEN_5331 | _GEN_2547;
  wire        _GEN_5460 = idx_1 == 5'h1E;
  wire        _GEN_5461 = commit_store_1 ? _GEN_5460 | _GEN_5333 | _GEN_2548 : _GEN_5333 | _GEN_2548;
  wire        _GEN_5462 = commit_store_1 ? (&idx_1) | _GEN_5334 | _GEN_2549 : _GEN_5334 | _GEN_2549;
  wire        _GEN_5463 = commit_store_1 | ~(commit_load_1 & _GEN_5400);
  wire        _GEN_5464 = commit_store_1 | ~(commit_load_1 & _GEN_5402);
  wire        _GEN_5465 = commit_store_1 | ~(commit_load_1 & _GEN_5404);
  wire        _GEN_5466 = commit_store_1 | ~(commit_load_1 & _GEN_5406);
  wire        _GEN_5467 = commit_store_1 | ~(commit_load_1 & _GEN_5408);
  wire        _GEN_5468 = commit_store_1 | ~(commit_load_1 & _GEN_5410);
  wire        _GEN_5469 = commit_store_1 | ~(commit_load_1 & _GEN_5412);
  wire        _GEN_5470 = commit_store_1 | ~(commit_load_1 & _GEN_5414);
  wire        _GEN_5471 = commit_store_1 | ~(commit_load_1 & _GEN_5416);
  wire        _GEN_5472 = commit_store_1 | ~(commit_load_1 & _GEN_5418);
  wire        _GEN_5473 = commit_store_1 | ~(commit_load_1 & _GEN_5420);
  wire        _GEN_5474 = commit_store_1 | ~(commit_load_1 & _GEN_5422);
  wire        _GEN_5475 = commit_store_1 | ~(commit_load_1 & _GEN_5424);
  wire        _GEN_5476 = commit_store_1 | ~(commit_load_1 & _GEN_5426);
  wire        _GEN_5477 = commit_store_1 | ~(commit_load_1 & _GEN_5428);
  wire        _GEN_5478 = commit_store_1 | ~(commit_load_1 & _GEN_5430);
  wire        _GEN_5479 = commit_store_1 | ~(commit_load_1 & _GEN_5432);
  wire        _GEN_5480 = commit_store_1 | ~(commit_load_1 & _GEN_5434);
  wire        _GEN_5481 = commit_store_1 | ~(commit_load_1 & _GEN_5436);
  wire        _GEN_5482 = commit_store_1 | ~(commit_load_1 & _GEN_5438);
  wire        _GEN_5483 = commit_store_1 | ~(commit_load_1 & _GEN_5440);
  wire        _GEN_5484 = commit_store_1 | ~(commit_load_1 & _GEN_5442);
  wire        _GEN_5485 = commit_store_1 | ~(commit_load_1 & _GEN_5444);
  wire        _GEN_5486 = commit_store_1 | ~(commit_load_1 & _GEN_5446);
  wire        _GEN_5487 = commit_store_1 | ~(commit_load_1 & _GEN_5448);
  wire        _GEN_5488 = commit_store_1 | ~(commit_load_1 & _GEN_5450);
  wire        _GEN_5489 = commit_store_1 | ~(commit_load_1 & _GEN_5452);
  wire        _GEN_5490 = commit_store_1 | ~(commit_load_1 & _GEN_5454);
  wire        _GEN_5491 = commit_store_1 | ~(commit_load_1 & _GEN_5456);
  wire        _GEN_5492 = commit_store_1 | ~(commit_load_1 & _GEN_5458);
  wire        _GEN_5493 = commit_store_1 | ~(commit_load_1 & _GEN_5460);
  wire        _GEN_5494 = commit_store_1 | ~(commit_load_1 & (&idx_1));
  wire        _GEN_5495 = idx_2 == 5'h0;
  wire        _GEN_5496 = commit_store_2 & _GEN_5495;
  wire        _GEN_5497 = idx_2 == 5'h1;
  wire        _GEN_5498 = commit_store_2 & _GEN_5497;
  wire        _GEN_5499 = idx_2 == 5'h2;
  wire        _GEN_5500 = commit_store_2 & _GEN_5499;
  wire        _GEN_5501 = idx_2 == 5'h3;
  wire        _GEN_5502 = commit_store_2 & _GEN_5501;
  wire        _GEN_5503 = idx_2 == 5'h4;
  wire        _GEN_5504 = commit_store_2 & _GEN_5503;
  wire        _GEN_5505 = idx_2 == 5'h5;
  wire        _GEN_5506 = commit_store_2 & _GEN_5505;
  wire        _GEN_5507 = idx_2 == 5'h6;
  wire        _GEN_5508 = commit_store_2 & _GEN_5507;
  wire        _GEN_5509 = idx_2 == 5'h7;
  wire        _GEN_5510 = commit_store_2 & _GEN_5509;
  wire        _GEN_5511 = idx_2 == 5'h8;
  wire        _GEN_5512 = commit_store_2 & _GEN_5511;
  wire        _GEN_5513 = idx_2 == 5'h9;
  wire        _GEN_5514 = commit_store_2 & _GEN_5513;
  wire        _GEN_5515 = idx_2 == 5'hA;
  wire        _GEN_5516 = commit_store_2 & _GEN_5515;
  wire        _GEN_5517 = idx_2 == 5'hB;
  wire        _GEN_5518 = commit_store_2 & _GEN_5517;
  wire        _GEN_5519 = idx_2 == 5'hC;
  wire        _GEN_5520 = commit_store_2 & _GEN_5519;
  wire        _GEN_5521 = idx_2 == 5'hD;
  wire        _GEN_5522 = commit_store_2 & _GEN_5521;
  wire        _GEN_5523 = idx_2 == 5'hE;
  wire        _GEN_5524 = commit_store_2 & _GEN_5523;
  wire        _GEN_5525 = idx_2 == 5'hF;
  wire        _GEN_5526 = commit_store_2 & _GEN_5525;
  wire        _GEN_5527 = idx_2 == 5'h10;
  wire        _GEN_5528 = commit_store_2 & _GEN_5527;
  wire        _GEN_5529 = idx_2 == 5'h11;
  wire        _GEN_5530 = commit_store_2 & _GEN_5529;
  wire        _GEN_5531 = idx_2 == 5'h12;
  wire        _GEN_5532 = commit_store_2 & _GEN_5531;
  wire        _GEN_5533 = idx_2 == 5'h13;
  wire        _GEN_5534 = commit_store_2 & _GEN_5533;
  wire        _GEN_5535 = idx_2 == 5'h14;
  wire        _GEN_5536 = commit_store_2 & _GEN_5535;
  wire        _GEN_5537 = idx_2 == 5'h15;
  wire        _GEN_5538 = commit_store_2 & _GEN_5537;
  wire        _GEN_5539 = idx_2 == 5'h16;
  wire        _GEN_5540 = commit_store_2 & _GEN_5539;
  wire        _GEN_5541 = idx_2 == 5'h17;
  wire        _GEN_5542 = commit_store_2 & _GEN_5541;
  wire        _GEN_5543 = idx_2 == 5'h18;
  wire        _GEN_5544 = commit_store_2 & _GEN_5543;
  wire        _GEN_5545 = idx_2 == 5'h19;
  wire        _GEN_5546 = commit_store_2 & _GEN_5545;
  wire        _GEN_5547 = idx_2 == 5'h1A;
  wire        _GEN_5548 = commit_store_2 & _GEN_5547;
  wire        _GEN_5549 = idx_2 == 5'h1B;
  wire        _GEN_5550 = commit_store_2 & _GEN_5549;
  wire        _GEN_5551 = idx_2 == 5'h1C;
  wire        _GEN_5552 = commit_store_2 & _GEN_5551;
  wire        _GEN_5553 = idx_2 == 5'h1D;
  wire        _GEN_5554 = commit_store_2 & _GEN_5553;
  wire        _GEN_5555 = idx_2 == 5'h1E;
  wire        _GEN_5556 = commit_store_2 & _GEN_5555;
  wire        _GEN_5557 = commit_store_2 & (&idx_2);
  wire        _GEN_5558 = commit_store_2 | ~(commit_load_2 & _GEN_5495);
  wire        _GEN_5559 = commit_store_2 | ~(commit_load_2 & _GEN_5497);
  wire        _GEN_5560 = commit_store_2 | ~(commit_load_2 & _GEN_5499);
  wire        _GEN_5561 = commit_store_2 | ~(commit_load_2 & _GEN_5501);
  wire        _GEN_5562 = commit_store_2 | ~(commit_load_2 & _GEN_5503);
  wire        _GEN_5563 = commit_store_2 | ~(commit_load_2 & _GEN_5505);
  wire        _GEN_5564 = commit_store_2 | ~(commit_load_2 & _GEN_5507);
  wire        _GEN_5565 = commit_store_2 | ~(commit_load_2 & _GEN_5509);
  wire        _GEN_5566 = commit_store_2 | ~(commit_load_2 & _GEN_5511);
  wire        _GEN_5567 = commit_store_2 | ~(commit_load_2 & _GEN_5513);
  wire        _GEN_5568 = commit_store_2 | ~(commit_load_2 & _GEN_5515);
  wire        _GEN_5569 = commit_store_2 | ~(commit_load_2 & _GEN_5517);
  wire        _GEN_5570 = commit_store_2 | ~(commit_load_2 & _GEN_5519);
  wire        _GEN_5571 = commit_store_2 | ~(commit_load_2 & _GEN_5521);
  wire        _GEN_5572 = commit_store_2 | ~(commit_load_2 & _GEN_5523);
  wire        _GEN_5573 = commit_store_2 | ~(commit_load_2 & _GEN_5525);
  wire        _GEN_5574 = commit_store_2 | ~(commit_load_2 & _GEN_5527);
  wire        _GEN_5575 = commit_store_2 | ~(commit_load_2 & _GEN_5529);
  wire        _GEN_5576 = commit_store_2 | ~(commit_load_2 & _GEN_5531);
  wire        _GEN_5577 = commit_store_2 | ~(commit_load_2 & _GEN_5533);
  wire        _GEN_5578 = commit_store_2 | ~(commit_load_2 & _GEN_5535);
  wire        _GEN_5579 = commit_store_2 | ~(commit_load_2 & _GEN_5537);
  wire        _GEN_5580 = commit_store_2 | ~(commit_load_2 & _GEN_5539);
  wire        _GEN_5581 = commit_store_2 | ~(commit_load_2 & _GEN_5541);
  wire        _GEN_5582 = commit_store_2 | ~(commit_load_2 & _GEN_5543);
  wire        _GEN_5583 = commit_store_2 | ~(commit_load_2 & _GEN_5545);
  wire        _GEN_5584 = commit_store_2 | ~(commit_load_2 & _GEN_5547);
  wire        _GEN_5585 = commit_store_2 | ~(commit_load_2 & _GEN_5549);
  wire        _GEN_5586 = commit_store_2 | ~(commit_load_2 & _GEN_5551);
  wire        _GEN_5587 = commit_store_2 | ~(commit_load_2 & _GEN_5553);
  wire        _GEN_5588 = commit_store_2 | ~(commit_load_2 & _GEN_5555);
  wire        _GEN_5589 = commit_store_2 | ~(commit_load_2 & (&idx_2));
  wire        _GEN_5590 = idx_3 == 5'h0;
  wire        _GEN_5591 = idx_3 == 5'h1;
  wire        _GEN_5592 = idx_3 == 5'h2;
  wire        _GEN_5593 = idx_3 == 5'h3;
  wire        _GEN_5594 = idx_3 == 5'h4;
  wire        _GEN_5595 = idx_3 == 5'h5;
  wire        _GEN_5596 = idx_3 == 5'h6;
  wire        _GEN_5597 = idx_3 == 5'h7;
  wire        _GEN_5598 = idx_3 == 5'h8;
  wire        _GEN_5599 = idx_3 == 5'h9;
  wire        _GEN_5600 = idx_3 == 5'hA;
  wire        _GEN_5601 = idx_3 == 5'hB;
  wire        _GEN_5602 = idx_3 == 5'hC;
  wire        _GEN_5603 = idx_3 == 5'hD;
  wire        _GEN_5604 = idx_3 == 5'hE;
  wire        _GEN_5605 = idx_3 == 5'hF;
  wire        _GEN_5606 = idx_3 == 5'h10;
  wire        _GEN_5607 = idx_3 == 5'h11;
  wire        _GEN_5608 = idx_3 == 5'h12;
  wire        _GEN_5609 = idx_3 == 5'h13;
  wire        _GEN_5610 = idx_3 == 5'h14;
  wire        _GEN_5611 = idx_3 == 5'h15;
  wire        _GEN_5612 = idx_3 == 5'h16;
  wire        _GEN_5613 = idx_3 == 5'h17;
  wire        _GEN_5614 = idx_3 == 5'h18;
  wire        _GEN_5615 = idx_3 == 5'h19;
  wire        _GEN_5616 = idx_3 == 5'h1A;
  wire        _GEN_5617 = idx_3 == 5'h1B;
  wire        _GEN_5618 = idx_3 == 5'h1C;
  wire        _GEN_5619 = idx_3 == 5'h1D;
  wire        _GEN_5620 = idx_3 == 5'h1E;
  wire        _GEN_5621 = commit_store_3 | ~(commit_load_3 & _GEN_5590);
  wire        _GEN_5622 = commit_store_3 | ~(commit_load_3 & _GEN_5591);
  wire        _GEN_5623 = commit_store_3 | ~(commit_load_3 & _GEN_5592);
  wire        _GEN_5624 = commit_store_3 | ~(commit_load_3 & _GEN_5593);
  wire        _GEN_5625 = commit_store_3 | ~(commit_load_3 & _GEN_5594);
  wire        _GEN_5626 = commit_store_3 | ~(commit_load_3 & _GEN_5595);
  wire        _GEN_5627 = commit_store_3 | ~(commit_load_3 & _GEN_5596);
  wire        _GEN_5628 = commit_store_3 | ~(commit_load_3 & _GEN_5597);
  wire        _GEN_5629 = commit_store_3 | ~(commit_load_3 & _GEN_5598);
  wire        _GEN_5630 = commit_store_3 | ~(commit_load_3 & _GEN_5599);
  wire        _GEN_5631 = commit_store_3 | ~(commit_load_3 & _GEN_5600);
  wire        _GEN_5632 = commit_store_3 | ~(commit_load_3 & _GEN_5601);
  wire        _GEN_5633 = commit_store_3 | ~(commit_load_3 & _GEN_5602);
  wire        _GEN_5634 = commit_store_3 | ~(commit_load_3 & _GEN_5603);
  wire        _GEN_5635 = commit_store_3 | ~(commit_load_3 & _GEN_5604);
  wire        _GEN_5636 = commit_store_3 | ~(commit_load_3 & _GEN_5605);
  wire        _GEN_5637 = commit_store_3 | ~(commit_load_3 & _GEN_5606);
  wire        _GEN_5638 = commit_store_3 | ~(commit_load_3 & _GEN_5607);
  wire        _GEN_5639 = commit_store_3 | ~(commit_load_3 & _GEN_5608);
  wire        _GEN_5640 = commit_store_3 | ~(commit_load_3 & _GEN_5609);
  wire        _GEN_5641 = commit_store_3 | ~(commit_load_3 & _GEN_5610);
  wire        _GEN_5642 = commit_store_3 | ~(commit_load_3 & _GEN_5611);
  wire        _GEN_5643 = commit_store_3 | ~(commit_load_3 & _GEN_5612);
  wire        _GEN_5644 = commit_store_3 | ~(commit_load_3 & _GEN_5613);
  wire        _GEN_5645 = commit_store_3 | ~(commit_load_3 & _GEN_5614);
  wire        _GEN_5646 = commit_store_3 | ~(commit_load_3 & _GEN_5615);
  wire        _GEN_5647 = commit_store_3 | ~(commit_load_3 & _GEN_5616);
  wire        _GEN_5648 = commit_store_3 | ~(commit_load_3 & _GEN_5617);
  wire        _GEN_5649 = commit_store_3 | ~(commit_load_3 & _GEN_5618);
  wire        _GEN_5650 = commit_store_3 | ~(commit_load_3 & _GEN_5619);
  wire        _GEN_5651 = commit_store_3 | ~(commit_load_3 & _GEN_5620);
  wire        _GEN_5652 = commit_store_3 | ~(commit_load_3 & (&idx_3));
  wire        _GEN_5653 = stq_head == 5'h0;
  wire        _GEN_5654 = _GEN_5653 | _GEN_5208;
  wire        _GEN_5655 = stq_head == 5'h1;
  wire        _GEN_5656 = _GEN_5655 | _GEN_5209;
  wire        _GEN_5657 = stq_head == 5'h2;
  wire        _GEN_5658 = _GEN_5657 | _GEN_5210;
  wire        _GEN_5659 = stq_head == 5'h3;
  wire        _GEN_5660 = _GEN_5659 | _GEN_5211;
  wire        _GEN_5661 = stq_head == 5'h4;
  wire        _GEN_5662 = _GEN_5661 | _GEN_5212;
  wire        _GEN_5663 = stq_head == 5'h5;
  wire        _GEN_5664 = _GEN_5663 | _GEN_5213;
  wire        _GEN_5665 = stq_head == 5'h6;
  wire        _GEN_5666 = _GEN_5665 | _GEN_5214;
  wire        _GEN_5667 = stq_head == 5'h7;
  wire        _GEN_5668 = _GEN_5667 | _GEN_5215;
  wire        _GEN_5669 = stq_head == 5'h8;
  wire        _GEN_5670 = _GEN_5669 | _GEN_5216;
  wire        _GEN_5671 = stq_head == 5'h9;
  wire        _GEN_5672 = _GEN_5671 | _GEN_5217;
  wire        _GEN_5673 = stq_head == 5'hA;
  wire        _GEN_5674 = _GEN_5673 | _GEN_5218;
  wire        _GEN_5675 = stq_head == 5'hB;
  wire        _GEN_5676 = _GEN_5675 | _GEN_5219;
  wire        _GEN_5677 = stq_head == 5'hC;
  wire        _GEN_5678 = _GEN_5677 | _GEN_5220;
  wire        _GEN_5679 = stq_head == 5'hD;
  wire        _GEN_5680 = _GEN_5679 | _GEN_5221;
  wire        _GEN_5681 = stq_head == 5'hE;
  wire        _GEN_5682 = _GEN_5681 | _GEN_5222;
  wire        _GEN_5683 = stq_head == 5'hF;
  wire        _GEN_5684 = _GEN_5683 | _GEN_5223;
  wire        _GEN_5685 = stq_head == 5'h10;
  wire        _GEN_5686 = _GEN_5685 | _GEN_5224;
  wire        _GEN_5687 = stq_head == 5'h11;
  wire        _GEN_5688 = _GEN_5687 | _GEN_5225;
  wire        _GEN_5689 = stq_head == 5'h12;
  wire        _GEN_5690 = _GEN_5689 | _GEN_5226;
  wire        _GEN_5691 = stq_head == 5'h13;
  wire        _GEN_5692 = _GEN_5691 | _GEN_5227;
  wire        _GEN_5693 = stq_head == 5'h14;
  wire        _GEN_5694 = _GEN_5693 | _GEN_5228;
  wire        _GEN_5695 = stq_head == 5'h15;
  wire        _GEN_5696 = _GEN_5695 | _GEN_5229;
  wire        _GEN_5697 = stq_head == 5'h16;
  wire        _GEN_5698 = _GEN_5697 | _GEN_5230;
  wire        _GEN_5699 = stq_head == 5'h17;
  wire        _GEN_5700 = _GEN_5699 | _GEN_5231;
  wire        _GEN_5701 = stq_head == 5'h18;
  wire        _GEN_5702 = _GEN_5701 | _GEN_5232;
  wire        _GEN_5703 = stq_head == 5'h19;
  wire        _GEN_5704 = _GEN_5703 | _GEN_5233;
  wire        _GEN_5705 = stq_head == 5'h1A;
  wire        _GEN_5706 = _GEN_5705 | _GEN_5234;
  wire        _GEN_5707 = stq_head == 5'h1B;
  wire        _GEN_5708 = _GEN_5707 | _GEN_5235;
  wire        _GEN_5709 = stq_head == 5'h1C;
  wire        _GEN_5710 = _GEN_5709 | _GEN_5236;
  wire        _GEN_5711 = stq_head == 5'h1D;
  wire        _GEN_5712 = _GEN_5711 | _GEN_5237;
  wire        _GEN_5713 = stq_head == 5'h1E;
  wire        _GEN_5714 = _GEN_5713 | _GEN_5238;
  wire        _GEN_5715 = (&stq_head) | _GEN_5239;
  wire        _GEN_5716 = clear_store & _GEN_5653;
  wire        _GEN_5717 = clear_store & _GEN_5655;
  wire        _GEN_5718 = clear_store & _GEN_5657;
  wire        _GEN_5719 = clear_store & _GEN_5659;
  wire        _GEN_5720 = clear_store & _GEN_5661;
  wire        _GEN_5721 = clear_store & _GEN_5663;
  wire        _GEN_5722 = clear_store & _GEN_5665;
  wire        _GEN_5723 = clear_store & _GEN_5667;
  wire        _GEN_5724 = clear_store & _GEN_5669;
  wire        _GEN_5725 = clear_store & _GEN_5671;
  wire        _GEN_5726 = clear_store & _GEN_5673;
  wire        _GEN_5727 = clear_store & _GEN_5675;
  wire        _GEN_5728 = clear_store & _GEN_5677;
  wire        _GEN_5729 = clear_store & _GEN_5679;
  wire        _GEN_5730 = clear_store & _GEN_5681;
  wire        _GEN_5731 = clear_store & _GEN_5683;
  wire        _GEN_5732 = clear_store & _GEN_5685;
  wire        _GEN_5733 = clear_store & _GEN_5687;
  wire        _GEN_5734 = clear_store & _GEN_5689;
  wire        _GEN_5735 = clear_store & _GEN_5691;
  wire        _GEN_5736 = clear_store & _GEN_5693;
  wire        _GEN_5737 = clear_store & _GEN_5695;
  wire        _GEN_5738 = clear_store & _GEN_5697;
  wire        _GEN_5739 = clear_store & _GEN_5699;
  wire        _GEN_5740 = clear_store & _GEN_5701;
  wire        _GEN_5741 = clear_store & _GEN_5703;
  wire        _GEN_5742 = clear_store & _GEN_5705;
  wire        _GEN_5743 = clear_store & _GEN_5707;
  wire        _GEN_5744 = clear_store & _GEN_5709;
  wire        _GEN_5745 = clear_store & _GEN_5711;
  wire        _GEN_5746 = clear_store & _GEN_5713;
  wire        _GEN_5747 = clear_store & (&stq_head);
  wire        _GEN_5748 = _io_hellacache_req_ready_output | ~_GEN_2;
  wire        _GEN_5749 = reset | io_core_exception;
  wire        _GEN_5750 = _GEN_5749 & reset;
  wire        _GEN_5751 = ~stq_0_bits_committed & ~stq_0_bits_succeeded;
  wire        _GEN_5752 = _GEN_5749 & (reset | _GEN_5751);
  wire        _GEN_5753 = ~stq_1_bits_committed & ~stq_1_bits_succeeded;
  wire        _GEN_5754 = _GEN_5749 & (reset | _GEN_5753);
  wire        _GEN_5755 = ~stq_2_bits_committed & ~stq_2_bits_succeeded;
  wire        _GEN_5756 = _GEN_5749 & (reset | _GEN_5755);
  wire        _GEN_5757 = ~stq_3_bits_committed & ~stq_3_bits_succeeded;
  wire        _GEN_5758 = _GEN_5749 & (reset | _GEN_5757);
  wire        _GEN_5759 = ~stq_4_bits_committed & ~stq_4_bits_succeeded;
  wire        _GEN_5760 = _GEN_5749 & (reset | _GEN_5759);
  wire        _GEN_5761 = ~stq_5_bits_committed & ~stq_5_bits_succeeded;
  wire        _GEN_5762 = _GEN_5749 & (reset | _GEN_5761);
  wire        _GEN_5763 = ~stq_6_bits_committed & ~stq_6_bits_succeeded;
  wire        _GEN_5764 = _GEN_5749 & (reset | _GEN_5763);
  wire        _GEN_5765 = ~stq_7_bits_committed & ~stq_7_bits_succeeded;
  wire        _GEN_5766 = _GEN_5749 & (reset | _GEN_5765);
  wire        _GEN_5767 = ~stq_8_bits_committed & ~stq_8_bits_succeeded;
  wire        _GEN_5768 = _GEN_5749 & (reset | _GEN_5767);
  wire        _GEN_5769 = ~stq_9_bits_committed & ~stq_9_bits_succeeded;
  wire        _GEN_5770 = _GEN_5749 & (reset | _GEN_5769);
  wire        _GEN_5771 = ~stq_10_bits_committed & ~stq_10_bits_succeeded;
  wire        _GEN_5772 = _GEN_5749 & (reset | _GEN_5771);
  wire        _GEN_5773 = ~stq_11_bits_committed & ~stq_11_bits_succeeded;
  wire        _GEN_5774 = _GEN_5749 & (reset | _GEN_5773);
  wire        _GEN_5775 = ~stq_12_bits_committed & ~stq_12_bits_succeeded;
  wire        _GEN_5776 = _GEN_5749 & (reset | _GEN_5775);
  wire        _GEN_5777 = ~stq_13_bits_committed & ~stq_13_bits_succeeded;
  wire        _GEN_5778 = _GEN_5749 & (reset | _GEN_5777);
  wire        _GEN_5779 = ~stq_14_bits_committed & ~stq_14_bits_succeeded;
  wire        _GEN_5780 = _GEN_5749 & (reset | _GEN_5779);
  wire        _GEN_5781 = ~stq_15_bits_committed & ~stq_15_bits_succeeded;
  wire        _GEN_5782 = _GEN_5749 & (reset | _GEN_5781);
  wire        _GEN_5783 = ~stq_16_bits_committed & ~stq_16_bits_succeeded;
  wire        _GEN_5784 = _GEN_5749 & (reset | _GEN_5783);
  wire        _GEN_5785 = ~stq_17_bits_committed & ~stq_17_bits_succeeded;
  wire        _GEN_5786 = _GEN_5749 & (reset | _GEN_5785);
  wire        _GEN_5787 = ~stq_18_bits_committed & ~stq_18_bits_succeeded;
  wire        _GEN_5788 = _GEN_5749 & (reset | _GEN_5787);
  wire        _GEN_5789 = ~stq_19_bits_committed & ~stq_19_bits_succeeded;
  wire        _GEN_5790 = _GEN_5749 & (reset | _GEN_5789);
  wire        _GEN_5791 = ~stq_20_bits_committed & ~stq_20_bits_succeeded;
  wire        _GEN_5792 = _GEN_5749 & (reset | _GEN_5791);
  wire        _GEN_5793 = ~stq_21_bits_committed & ~stq_21_bits_succeeded;
  wire        _GEN_5794 = _GEN_5749 & (reset | _GEN_5793);
  wire        _GEN_5795 = ~stq_22_bits_committed & ~stq_22_bits_succeeded;
  wire        _GEN_5796 = _GEN_5749 & (reset | _GEN_5795);
  wire        _GEN_5797 = ~stq_23_bits_committed & ~stq_23_bits_succeeded;
  wire        _GEN_5798 = _GEN_5749 & (reset | _GEN_5797);
  wire        _GEN_5799 = ~stq_24_bits_committed & ~stq_24_bits_succeeded;
  wire        _GEN_5800 = _GEN_5749 & (reset | _GEN_5799);
  wire        _GEN_5801 = ~stq_25_bits_committed & ~stq_25_bits_succeeded;
  wire        _GEN_5802 = _GEN_5749 & (reset | _GEN_5801);
  wire        _GEN_5803 = ~stq_26_bits_committed & ~stq_26_bits_succeeded;
  wire        _GEN_5804 = _GEN_5749 & (reset | _GEN_5803);
  wire        _GEN_5805 = ~stq_27_bits_committed & ~stq_27_bits_succeeded;
  wire        _GEN_5806 = _GEN_5749 & (reset | _GEN_5805);
  wire        _GEN_5807 = ~stq_28_bits_committed & ~stq_28_bits_succeeded;
  wire        _GEN_5808 = _GEN_5749 & (reset | _GEN_5807);
  wire        _GEN_5809 = ~stq_29_bits_committed & ~stq_29_bits_succeeded;
  wire        _GEN_5810 = _GEN_5749 & (reset | _GEN_5809);
  wire        _GEN_5811 = ~stq_30_bits_committed & ~stq_30_bits_succeeded;
  wire        _GEN_5812 = _GEN_5749 & (reset | _GEN_5811);
  wire        _GEN_5813 = ~stq_31_bits_committed & ~stq_31_bits_succeeded;
  wire        _GEN_5814 = _GEN_5749 & (reset | _GEN_5813);
  wire        _GEN_5815 = _GEN_2005 | ~_GEN_1653;
  wire        _GEN_5816 = _GEN_2006 | ~_GEN_1654;
  wire        _GEN_5817 = _GEN_2007 | ~_GEN_1655;
  wire        _GEN_5818 = _GEN_2008 | ~_GEN_1656;
  wire        _GEN_5819 = _GEN_2009 | ~_GEN_1657;
  wire        _GEN_5820 = _GEN_2010 | ~_GEN_1658;
  wire        _GEN_5821 = _GEN_2011 | ~_GEN_1659;
  wire        _GEN_5822 = _GEN_2012 | ~_GEN_1660;
  wire        _GEN_5823 = _GEN_2013 | ~_GEN_1661;
  wire        _GEN_5824 = _GEN_2014 | ~_GEN_1662;
  wire        _GEN_5825 = _GEN_2015 | ~_GEN_1663;
  wire        _GEN_5826 = _GEN_2016 | ~_GEN_1664;
  wire        _GEN_5827 = _GEN_2017 | ~_GEN_1665;
  wire        _GEN_5828 = _GEN_2018 | ~_GEN_1666;
  wire        _GEN_5829 = _GEN_2019 | ~_GEN_1667;
  wire        _GEN_5830 = _GEN_2020 | ~_GEN_1668;
  wire        _GEN_5831 = _GEN_2021 | ~_GEN_1669;
  wire        _GEN_5832 = _GEN_2022 | ~_GEN_1670;
  wire        _GEN_5833 = _GEN_2023 | ~_GEN_1671;
  wire        _GEN_5834 = _GEN_2024 | ~_GEN_1672;
  wire        _GEN_5835 = _GEN_2025 | ~_GEN_1673;
  wire        _GEN_5836 = _GEN_2026 | ~_GEN_1674;
  wire        _GEN_5837 = _GEN_2027 | ~_GEN_1675;
  wire        _GEN_5838 = _GEN_2028 | ~_GEN_1676;
  wire        _GEN_5839 = _GEN_2029 | ~_GEN_1677;
  wire        _GEN_5840 = _GEN_2030 | ~_GEN_1678;
  wire        _GEN_5841 = _GEN_2031 | ~_GEN_1679;
  wire        _GEN_5842 = _GEN_2032 | ~_GEN_1680;
  wire        _GEN_5843 = _GEN_2033 | ~_GEN_1681;
  wire        _GEN_5844 = _GEN_2034 | ~_GEN_1682;
  wire        _GEN_5845 = _GEN_2035 | ~_GEN_1683;
  wire        _GEN_5846 = _GEN_2036 | ~_GEN_1684;
  wire [5:0]  _ldq_retry_idx_idx_T_42 = _ldq_retry_idx_T_62 & _temp_bits_T_40 ? 6'h14 : _ldq_retry_idx_T_65 & _temp_bits_T_42 ? 6'h15 : _ldq_retry_idx_T_68 & _temp_bits_T_44 ? 6'h16 : _ldq_retry_idx_T_71 & _temp_bits_T_46 ? 6'h17 : _ldq_retry_idx_T_74 & _temp_bits_T_48 ? 6'h18 : _ldq_retry_idx_T_77 & _temp_bits_T_50 ? 6'h19 : _ldq_retry_idx_T_80 & _temp_bits_T_52 ? 6'h1A : _ldq_retry_idx_T_83 & _temp_bits_T_54 ? 6'h1B : _ldq_retry_idx_T_86 & _temp_bits_T_56 ? 6'h1C : _ldq_retry_idx_T_89 & _temp_bits_T_58 ? 6'h1D : _ldq_retry_idx_T_92 & _temp_bits_T_60 ? 6'h1E : ldq_31_bits_addr_valid & ldq_31_bits_addr_is_virtual & ~ldq_retry_idx_block_31 ? 6'h1F : _ldq_retry_idx_T_2 ? 6'h20 : _ldq_retry_idx_T_5 ? 6'h21 : _ldq_retry_idx_T_8 ? 6'h22 : _ldq_retry_idx_T_11 ? 6'h23 : _ldq_retry_idx_T_14 ? 6'h24 : _ldq_retry_idx_T_17 ? 6'h25 : _ldq_retry_idx_T_20 ? 6'h26 : _ldq_retry_idx_T_23 ? 6'h27 : _ldq_retry_idx_T_26 ? 6'h28 : _ldq_retry_idx_T_29 ? 6'h29 : _ldq_retry_idx_T_32 ? 6'h2A : _ldq_retry_idx_T_35 ? 6'h2B : _ldq_retry_idx_T_38 ? 6'h2C : _ldq_retry_idx_T_41 ? 6'h2D : _ldq_retry_idx_T_44 ? 6'h2E : _ldq_retry_idx_T_47 ? 6'h2F : _ldq_retry_idx_T_50 ? 6'h30 : _ldq_retry_idx_T_53 ? 6'h31 : _ldq_retry_idx_T_56 ? 6'h32 : _ldq_retry_idx_T_59 ? 6'h33 : _ldq_retry_idx_T_62 ? 6'h34 : _ldq_retry_idx_T_65 ? 6'h35 : _ldq_retry_idx_T_68 ? 6'h36 : _ldq_retry_idx_T_71 ? 6'h37 : _ldq_retry_idx_T_74 ? 6'h38 : _ldq_retry_idx_T_77 ? 6'h39 : _ldq_retry_idx_T_80 ? 6'h3A : _ldq_retry_idx_T_83 ? 6'h3B : _ldq_retry_idx_T_86 ? 6'h3C : _ldq_retry_idx_T_89 ? 6'h3D : {5'h1F, ~_ldq_retry_idx_T_92};
  wire [5:0]  _stq_retry_idx_idx_T_42 = _stq_retry_idx_T_20 & stq_commit_head < 5'h15 ? 6'h14 : _stq_retry_idx_T_21 & stq_commit_head < 5'h16 ? 6'h15 : _stq_retry_idx_T_22 & stq_commit_head < 5'h17 ? 6'h16 : _stq_retry_idx_T_23 & stq_commit_head[4:3] != 2'h3 ? 6'h17 : _stq_retry_idx_T_24 & stq_commit_head < 5'h19 ? 6'h18 : _stq_retry_idx_T_25 & stq_commit_head < 5'h1A ? 6'h19 : _stq_retry_idx_T_26 & stq_commit_head < 5'h1B ? 6'h1A : _stq_retry_idx_T_27 & stq_commit_head[4:2] != 3'h7 ? 6'h1B : _stq_retry_idx_T_28 & stq_commit_head < 5'h1D ? 6'h1C : _stq_retry_idx_T_29 & stq_commit_head[4:1] != 4'hF ? 6'h1D : _stq_retry_idx_T_30 & stq_commit_head != 5'h1F ? 6'h1E : stq_31_bits_addr_valid & stq_31_bits_addr_is_virtual ? 6'h1F : _stq_retry_idx_T ? 6'h20 : _stq_retry_idx_T_1 ? 6'h21 : _stq_retry_idx_T_2 ? 6'h22 : _stq_retry_idx_T_3 ? 6'h23 : _stq_retry_idx_T_4 ? 6'h24 : _stq_retry_idx_T_5 ? 6'h25 : _stq_retry_idx_T_6 ? 6'h26 : _stq_retry_idx_T_7 ? 6'h27 : _stq_retry_idx_T_8 ? 6'h28 : _stq_retry_idx_T_9 ? 6'h29 : _stq_retry_idx_T_10 ? 6'h2A : _stq_retry_idx_T_11 ? 6'h2B : _stq_retry_idx_T_12 ? 6'h2C : _stq_retry_idx_T_13 ? 6'h2D : _stq_retry_idx_T_14 ? 6'h2E : _stq_retry_idx_T_15 ? 6'h2F : _stq_retry_idx_T_16 ? 6'h30 : _stq_retry_idx_T_17 ? 6'h31 : _stq_retry_idx_T_18 ? 6'h32 : _stq_retry_idx_T_19 ? 6'h33 : _stq_retry_idx_T_20 ? 6'h34 : _stq_retry_idx_T_21 ? 6'h35 : _stq_retry_idx_T_22 ? 6'h36 : _stq_retry_idx_T_23 ? 6'h37 : _stq_retry_idx_T_24 ? 6'h38 : _stq_retry_idx_T_25 ? 6'h39 : _stq_retry_idx_T_26 ? 6'h3A : _stq_retry_idx_T_27 ? 6'h3B : _stq_retry_idx_T_28 ? 6'h3C : _stq_retry_idx_T_29 ? 6'h3D : {5'h1F, ~_stq_retry_idx_T_30};
  wire [5:0]  _ldq_wakeup_idx_idx_T_42 = _ldq_wakeup_idx_T_167 & _temp_bits_T_40 ? 6'h14 : _ldq_wakeup_idx_T_175 & _temp_bits_T_42 ? 6'h15 : _ldq_wakeup_idx_T_183 & _temp_bits_T_44 ? 6'h16 : _ldq_wakeup_idx_T_191 & _temp_bits_T_46 ? 6'h17 : _ldq_wakeup_idx_T_199 & _temp_bits_T_48 ? 6'h18 : _ldq_wakeup_idx_T_207 & _temp_bits_T_50 ? 6'h19 : _ldq_wakeup_idx_T_215 & _temp_bits_T_52 ? 6'h1A : _ldq_wakeup_idx_T_223 & _temp_bits_T_54 ? 6'h1B : _ldq_wakeup_idx_T_231 & _temp_bits_T_56 ? 6'h1C : _ldq_wakeup_idx_T_239 & _temp_bits_T_58 ? 6'h1D : _ldq_wakeup_idx_T_247 & _temp_bits_T_60 ? 6'h1E : ldq_31_bits_addr_valid & ~ldq_31_bits_executed & ~ldq_31_bits_succeeded & ~ldq_31_bits_addr_is_virtual & ~ldq_retry_idx_block_31 ? 6'h1F : _ldq_wakeup_idx_T_7 ? 6'h20 : _ldq_wakeup_idx_T_15 ? 6'h21 : _ldq_wakeup_idx_T_23 ? 6'h22 : _ldq_wakeup_idx_T_31 ? 6'h23 : _ldq_wakeup_idx_T_39 ? 6'h24 : _ldq_wakeup_idx_T_47 ? 6'h25 : _ldq_wakeup_idx_T_55 ? 6'h26 : _ldq_wakeup_idx_T_63 ? 6'h27 : _ldq_wakeup_idx_T_71 ? 6'h28 : _ldq_wakeup_idx_T_79 ? 6'h29 : _ldq_wakeup_idx_T_87 ? 6'h2A : _ldq_wakeup_idx_T_95 ? 6'h2B : _ldq_wakeup_idx_T_103 ? 6'h2C : _ldq_wakeup_idx_T_111 ? 6'h2D : _ldq_wakeup_idx_T_119 ? 6'h2E : _ldq_wakeup_idx_T_127 ? 6'h2F : _ldq_wakeup_idx_T_135 ? 6'h30 : _ldq_wakeup_idx_T_143 ? 6'h31 : _ldq_wakeup_idx_T_151 ? 6'h32 : _ldq_wakeup_idx_T_159 ? 6'h33 : _ldq_wakeup_idx_T_167 ? 6'h34 : _ldq_wakeup_idx_T_175 ? 6'h35 : _ldq_wakeup_idx_T_183 ? 6'h36 : _ldq_wakeup_idx_T_191 ? 6'h37 : _ldq_wakeup_idx_T_199 ? 6'h38 : _ldq_wakeup_idx_T_207 ? 6'h39 : _ldq_wakeup_idx_T_215 ? 6'h3A : _ldq_wakeup_idx_T_223 ? 6'h3B : _ldq_wakeup_idx_T_231 ? 6'h3C : _ldq_wakeup_idx_T_239 ? 6'h3D : {5'h1F, ~_ldq_wakeup_idx_T_247};
  always @(posedge clock) begin
    if (_GEN_1434)
      assert__assert_52: assert(casez_tmp_459);
    if (_GEN_1473)
      assert__assert_58: assert(casez_tmp_493);
    if (_GEN_1543)
      assert__assert_95: assert(casez_tmp_527);
    if (_GEN_1548)
      assert__assert_97: assert(casez_tmp_531);
    if (_GEN_1553)
      assert__assert_99: assert(casez_tmp_535);
    if (_GEN_1558)
      assert__assert_101: assert(casez_tmp_539);
    ldq_0_valid <= ~_GEN_5749 & _GEN_5621 & _GEN_5558 & _GEN_5463 & (_GEN_5336 ? ~_GEN_5240 & _GEN_2169 : ~_GEN_5335 & _GEN_2169);
    if (_GEN_2262) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_0_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_0_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_0_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_0_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_0_bits_st_dep_mask <= _GEN_2166;
      ldq_0_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2070) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_0_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_0_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_0_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_0_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_0_bits_st_dep_mask <= _GEN_2069;
      ldq_0_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1781) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_0_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_0_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_0_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_0_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_0_bits_st_dep_mask <= _GEN_1685;
      ldq_0_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1589) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_0_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_0_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_0_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_0_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_0_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_0_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_0_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_0_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_0_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_0_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_0_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_0_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_0_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_0_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_0_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_0_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_0_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_0_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_0_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_0_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_0_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_0_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_0_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_0_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_0_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_0_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_0_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_0_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_0_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_0_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_0_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_0_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_0_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_0_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_0_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_0_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_0_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_0_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_0_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_0_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_0_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_0_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_0_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_0_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_0_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_0_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_0_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_0_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_0_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_0_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_0_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_0_bits_st_dep_mask <= next_live_store_mask;
      ldq_0_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_0_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_0_bits_st_dep_mask;
    if (ldq_0_valid)
      ldq_0_bits_uop_br_mask <= ldq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2262)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2070)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1781)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1589)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2742) begin
      if (_exe_tlb_uop_T_9)
        ldq_0_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_0_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_0_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_0_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_0_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_0_bits_addr_bits <= casez_tmp_202;
        else
          ldq_0_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_0_bits_addr_bits <= _GEN_280;
      ldq_0_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_0_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2646) begin
      if (_exe_tlb_uop_T_2)
        ldq_0_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_0_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_0_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_0_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_0_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_0_bits_addr_bits <= casez_tmp_202;
        else
          ldq_0_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_0_bits_addr_bits <= _GEN_274;
      ldq_0_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_0_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2262)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2070)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1781)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1589)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    if (mem_xcpt_valids_1 & mem_xcpt_uops_1_uses_ldq) begin
      ldq_0_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h0 | _GEN_2551 | _GEN_2263;
      ldq_1_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h1 | _GEN_2552 | _GEN_2265;
      ldq_2_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h2 | _GEN_2553 | _GEN_2267;
      ldq_3_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h3 | _GEN_2554 | _GEN_2269;
      ldq_4_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h4 | _GEN_2555 | _GEN_2271;
      ldq_5_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h5 | _GEN_2556 | _GEN_2273;
      ldq_6_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h6 | _GEN_2557 | _GEN_2275;
      ldq_7_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h7 | _GEN_2558 | _GEN_2277;
      ldq_8_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h8 | _GEN_2559 | _GEN_2279;
      ldq_9_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h9 | _GEN_2560 | _GEN_2281;
      ldq_10_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'hA | _GEN_2561 | _GEN_2283;
      ldq_11_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'hB | _GEN_2562 | _GEN_2285;
      ldq_12_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'hC | _GEN_2563 | _GEN_2287;
      ldq_13_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'hD | _GEN_2564 | _GEN_2289;
      ldq_14_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'hE | _GEN_2565 | _GEN_2291;
      ldq_15_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'hF | _GEN_2566 | _GEN_2293;
      ldq_16_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h10 | _GEN_2567 | _GEN_2295;
      ldq_17_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h11 | _GEN_2568 | _GEN_2297;
      ldq_18_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h12 | _GEN_2569 | _GEN_2299;
      ldq_19_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h13 | _GEN_2570 | _GEN_2301;
      ldq_20_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h14 | _GEN_2571 | _GEN_2303;
      ldq_21_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h15 | _GEN_2572 | _GEN_2305;
      ldq_22_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h16 | _GEN_2573 | _GEN_2307;
      ldq_23_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h17 | _GEN_2574 | _GEN_2309;
      ldq_24_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h18 | _GEN_2575 | _GEN_2311;
      ldq_25_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h19 | _GEN_2576 | _GEN_2313;
      ldq_26_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h1A | _GEN_2577 | _GEN_2315;
      ldq_27_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h1B | _GEN_2578 | _GEN_2317;
      ldq_28_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h1C | _GEN_2579 | _GEN_2319;
      ldq_29_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h1D | _GEN_2580 | _GEN_2321;
      ldq_30_bits_uop_exception <= mem_xcpt_uops_1_ldq_idx == 5'h1E | _GEN_2581 | _GEN_2323;
      ldq_31_bits_uop_exception <= (&mem_xcpt_uops_1_ldq_idx) | _GEN_2582 | _GEN_2325;
    end
    else begin
      ldq_0_bits_uop_exception <= _GEN_2551 | _GEN_2263;
      ldq_1_bits_uop_exception <= _GEN_2552 | _GEN_2265;
      ldq_2_bits_uop_exception <= _GEN_2553 | _GEN_2267;
      ldq_3_bits_uop_exception <= _GEN_2554 | _GEN_2269;
      ldq_4_bits_uop_exception <= _GEN_2555 | _GEN_2271;
      ldq_5_bits_uop_exception <= _GEN_2556 | _GEN_2273;
      ldq_6_bits_uop_exception <= _GEN_2557 | _GEN_2275;
      ldq_7_bits_uop_exception <= _GEN_2558 | _GEN_2277;
      ldq_8_bits_uop_exception <= _GEN_2559 | _GEN_2279;
      ldq_9_bits_uop_exception <= _GEN_2560 | _GEN_2281;
      ldq_10_bits_uop_exception <= _GEN_2561 | _GEN_2283;
      ldq_11_bits_uop_exception <= _GEN_2562 | _GEN_2285;
      ldq_12_bits_uop_exception <= _GEN_2563 | _GEN_2287;
      ldq_13_bits_uop_exception <= _GEN_2564 | _GEN_2289;
      ldq_14_bits_uop_exception <= _GEN_2565 | _GEN_2291;
      ldq_15_bits_uop_exception <= _GEN_2566 | _GEN_2293;
      ldq_16_bits_uop_exception <= _GEN_2567 | _GEN_2295;
      ldq_17_bits_uop_exception <= _GEN_2568 | _GEN_2297;
      ldq_18_bits_uop_exception <= _GEN_2569 | _GEN_2299;
      ldq_19_bits_uop_exception <= _GEN_2570 | _GEN_2301;
      ldq_20_bits_uop_exception <= _GEN_2571 | _GEN_2303;
      ldq_21_bits_uop_exception <= _GEN_2572 | _GEN_2305;
      ldq_22_bits_uop_exception <= _GEN_2573 | _GEN_2307;
      ldq_23_bits_uop_exception <= _GEN_2574 | _GEN_2309;
      ldq_24_bits_uop_exception <= _GEN_2575 | _GEN_2311;
      ldq_25_bits_uop_exception <= _GEN_2576 | _GEN_2313;
      ldq_26_bits_uop_exception <= _GEN_2577 | _GEN_2315;
      ldq_27_bits_uop_exception <= _GEN_2578 | _GEN_2317;
      ldq_28_bits_uop_exception <= _GEN_2579 | _GEN_2319;
      ldq_29_bits_uop_exception <= _GEN_2580 | _GEN_2321;
      ldq_30_bits_uop_exception <= _GEN_2581 | _GEN_2323;
      ldq_31_bits_uop_exception <= _GEN_2582 | _GEN_2325;
    end
    ldq_0_bits_addr_valid <= ~_GEN_5749 & _GEN_5621 & _GEN_5558 & _GEN_5463 & (_GEN_5336 ? ~_GEN_5240 & _GEN_2743 : ~_GEN_5335 & _GEN_2743);
    ldq_0_bits_executed <= ~_GEN_5749 & _GEN_5621 & _GEN_5558 & _GEN_5463 & _GEN_5368 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1474) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1435)) & ((_GEN_1426 ? (_GEN_5077 ? (|lcam_ldq_idx_1) & _GEN_5045 : ~(_GEN_1425 & ~(|lcam_ldq_idx_1)) & _GEN_5045) : _GEN_5045) | (dis_ld_val_3 ? ~_GEN_2168 & _GEN_1845 : ~_GEN_2070 & _GEN_1845));
    ldq_0_bits_succeeded <= _GEN_5621 & _GEN_5558 & _GEN_5463 & _GEN_5368 & (_GEN_5145 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h0 ? _ldq_bits_succeeded_T_1 : _GEN_5080 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h0 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2168 & _GEN_1877 : ~_GEN_2070 & _GEN_1877) : casez_tmp_490) : casez_tmp_524);
    ldq_0_bits_order_fail <= _GEN_5621 & _GEN_5558 & _GEN_5463 & _GEN_5368 & (_GEN_327 ? _GEN_2932 : _GEN_330 ? _GEN_331 | _GEN_2932 : _GEN_333 | _GEN_2932);
    ldq_0_bits_observed <= _GEN_327 | _GEN_284 | (dis_ld_val_3 ? ~_GEN_2168 & _GEN_1941 : ~_GEN_2070 & _GEN_1941);
    ldq_0_bits_forward_std_val <= _GEN_5621 & _GEN_5558 & _GEN_5463 & _GEN_5368 & (~_GEN_1508 & _GEN_5144 | ~_GEN_1468 & _GEN_5079 | (dis_ld_val_3 ? ~_GEN_2168 & _GEN_1973 : ~_GEN_2070 & _GEN_1973));
    if (_GEN_5145) begin
      if (_GEN_5080) begin
      end
      else
        ldq_0_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_0_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_1_valid <= ~_GEN_5749 & _GEN_5622 & _GEN_5559 & _GEN_5464 & (_GEN_5336 ? ~_GEN_5241 & _GEN_2172 : ~_GEN_5337 & _GEN_2172);
    if (_GEN_2264) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_1_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_1_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_1_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_1_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_1_bits_st_dep_mask <= _GEN_2166;
      ldq_1_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2071) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_1_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_1_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_1_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_1_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_1_bits_st_dep_mask <= _GEN_2069;
      ldq_1_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1782) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_1_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_1_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_1_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_1_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_1_bits_st_dep_mask <= _GEN_1685;
      ldq_1_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1590) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_1_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_1_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_1_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_1_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_1_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_1_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_1_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_1_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_1_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_1_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_1_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_1_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_1_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_1_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_1_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_1_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_1_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_1_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_1_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_1_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_1_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_1_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_1_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_1_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_1_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_1_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_1_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_1_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_1_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_1_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_1_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_1_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_1_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_1_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_1_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_1_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_1_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_1_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_1_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_1_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_1_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_1_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_1_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_1_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_1_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_1_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_1_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_1_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_1_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_1_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_1_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_1_bits_st_dep_mask <= next_live_store_mask;
      ldq_1_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_1_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_1_bits_st_dep_mask;
    if (ldq_1_valid)
      ldq_1_bits_uop_br_mask <= ldq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2264)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2071)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1782)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1590)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2744) begin
      if (_exe_tlb_uop_T_9)
        ldq_1_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_1_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_1_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_1_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_1_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_1_bits_addr_bits <= casez_tmp_202;
        else
          ldq_1_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_1_bits_addr_bits <= _GEN_280;
      ldq_1_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_1_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2647) begin
      if (_exe_tlb_uop_T_2)
        ldq_1_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_1_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_1_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_1_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_1_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_1_bits_addr_bits <= casez_tmp_202;
        else
          ldq_1_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_1_bits_addr_bits <= _GEN_274;
      ldq_1_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_1_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2264)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2071)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1782)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1590)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_1_bits_addr_valid <= ~_GEN_5749 & _GEN_5622 & _GEN_5559 & _GEN_5464 & (_GEN_5336 ? ~_GEN_5241 & _GEN_2745 : ~_GEN_5337 & _GEN_2745);
    ldq_1_bits_executed <= ~_GEN_5749 & _GEN_5622 & _GEN_5559 & _GEN_5464 & _GEN_5369 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1475) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1436)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_336 & _GEN_5046 : ~(_GEN_1425 & _GEN_336) & _GEN_5046) : _GEN_5046) | (dis_ld_val_3 ? ~_GEN_2171 & _GEN_1846 : ~_GEN_2071 & _GEN_1846));
    ldq_1_bits_succeeded <= _GEN_5622 & _GEN_5559 & _GEN_5464 & _GEN_5369 & (_GEN_5147 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1 ? _ldq_bits_succeeded_T_1 : _GEN_5082 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2171 & _GEN_1878 : ~_GEN_2071 & _GEN_1878) : casez_tmp_490) : casez_tmp_524);
    ldq_1_bits_order_fail <= _GEN_5622 & _GEN_5559 & _GEN_5464 & _GEN_5369 & (_GEN_380 ? _GEN_2933 : _GEN_382 ? _GEN_383 | _GEN_2933 : _GEN_385 | _GEN_2933);
    ldq_1_bits_observed <= _GEN_380 | _GEN_367 | (dis_ld_val_3 ? ~_GEN_2171 & _GEN_1942 : ~_GEN_2071 & _GEN_1942);
    ldq_1_bits_forward_std_val <= _GEN_5622 & _GEN_5559 & _GEN_5464 & _GEN_5369 & (~_GEN_1508 & _GEN_5146 | ~_GEN_1468 & _GEN_5081 | (dis_ld_val_3 ? ~_GEN_2171 & _GEN_1974 : ~_GEN_2071 & _GEN_1974));
    if (_GEN_5147) begin
      if (_GEN_5082) begin
      end
      else
        ldq_1_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_1_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_2_valid <= ~_GEN_5749 & _GEN_5623 & _GEN_5560 & _GEN_5465 & (_GEN_5336 ? ~_GEN_5242 & _GEN_2175 : ~_GEN_5338 & _GEN_2175);
    if (_GEN_2266) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_2_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_2_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_2_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_2_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_2_bits_st_dep_mask <= _GEN_2166;
      ldq_2_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2072) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_2_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_2_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_2_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_2_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_2_bits_st_dep_mask <= _GEN_2069;
      ldq_2_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1783) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_2_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_2_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_2_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_2_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_2_bits_st_dep_mask <= _GEN_1685;
      ldq_2_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1591) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_2_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_2_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_2_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_2_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_2_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_2_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_2_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_2_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_2_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_2_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_2_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_2_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_2_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_2_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_2_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_2_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_2_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_2_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_2_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_2_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_2_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_2_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_2_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_2_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_2_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_2_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_2_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_2_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_2_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_2_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_2_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_2_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_2_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_2_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_2_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_2_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_2_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_2_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_2_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_2_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_2_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_2_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_2_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_2_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_2_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_2_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_2_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_2_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_2_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_2_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_2_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_2_bits_st_dep_mask <= next_live_store_mask;
      ldq_2_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_2_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_2_bits_st_dep_mask;
    if (ldq_2_valid)
      ldq_2_bits_uop_br_mask <= ldq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2266)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2072)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1783)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1591)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2746) begin
      if (_exe_tlb_uop_T_9)
        ldq_2_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_2_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_2_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_2_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_2_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_2_bits_addr_bits <= casez_tmp_202;
        else
          ldq_2_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_2_bits_addr_bits <= _GEN_280;
      ldq_2_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_2_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2648) begin
      if (_exe_tlb_uop_T_2)
        ldq_2_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_2_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_2_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_2_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_2_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_2_bits_addr_bits <= casez_tmp_202;
        else
          ldq_2_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_2_bits_addr_bits <= _GEN_274;
      ldq_2_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_2_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2266)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2072)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1783)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1591)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_2_bits_addr_valid <= ~_GEN_5749 & _GEN_5623 & _GEN_5560 & _GEN_5465 & (_GEN_5336 ? ~_GEN_5242 & _GEN_2747 : ~_GEN_5338 & _GEN_2747);
    ldq_2_bits_executed <= ~_GEN_5749 & _GEN_5623 & _GEN_5560 & _GEN_5465 & _GEN_5370 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1476) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1437)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_337 & _GEN_5047 : ~(_GEN_1425 & _GEN_337) & _GEN_5047) : _GEN_5047) | (dis_ld_val_3 ? ~_GEN_2174 & _GEN_1847 : ~_GEN_2072 & _GEN_1847));
    ldq_2_bits_succeeded <= _GEN_5623 & _GEN_5560 & _GEN_5465 & _GEN_5370 & (_GEN_5149 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h2 ? _ldq_bits_succeeded_T_1 : _GEN_5084 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h2 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2174 & _GEN_1879 : ~_GEN_2072 & _GEN_1879) : casez_tmp_490) : casez_tmp_524);
    ldq_2_bits_order_fail <= _GEN_5623 & _GEN_5560 & _GEN_5465 & _GEN_5370 & (_GEN_403 ? _GEN_2934 : _GEN_405 ? _GEN_406 | _GEN_2934 : _GEN_408 | _GEN_2934);
    ldq_2_bits_observed <= _GEN_403 | _GEN_390 | (dis_ld_val_3 ? ~_GEN_2174 & _GEN_1943 : ~_GEN_2072 & _GEN_1943);
    ldq_2_bits_forward_std_val <= _GEN_5623 & _GEN_5560 & _GEN_5465 & _GEN_5370 & (~_GEN_1508 & _GEN_5148 | ~_GEN_1468 & _GEN_5083 | (dis_ld_val_3 ? ~_GEN_2174 & _GEN_1975 : ~_GEN_2072 & _GEN_1975));
    if (_GEN_5149) begin
      if (_GEN_5084) begin
      end
      else
        ldq_2_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_2_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_3_valid <= ~_GEN_5749 & _GEN_5624 & _GEN_5561 & _GEN_5466 & (_GEN_5336 ? ~_GEN_5243 & _GEN_2178 : ~_GEN_5339 & _GEN_2178);
    if (_GEN_2268) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_3_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_3_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_3_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_3_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_3_bits_st_dep_mask <= _GEN_2166;
      ldq_3_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2073) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_3_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_3_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_3_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_3_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_3_bits_st_dep_mask <= _GEN_2069;
      ldq_3_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1784) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_3_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_3_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_3_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_3_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_3_bits_st_dep_mask <= _GEN_1685;
      ldq_3_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1592) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_3_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_3_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_3_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_3_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_3_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_3_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_3_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_3_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_3_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_3_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_3_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_3_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_3_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_3_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_3_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_3_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_3_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_3_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_3_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_3_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_3_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_3_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_3_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_3_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_3_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_3_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_3_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_3_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_3_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_3_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_3_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_3_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_3_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_3_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_3_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_3_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_3_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_3_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_3_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_3_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_3_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_3_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_3_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_3_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_3_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_3_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_3_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_3_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_3_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_3_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_3_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_3_bits_st_dep_mask <= next_live_store_mask;
      ldq_3_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_3_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_3_bits_st_dep_mask;
    if (ldq_3_valid)
      ldq_3_bits_uop_br_mask <= ldq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2268)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2073)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1784)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1592)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2748) begin
      if (_exe_tlb_uop_T_9)
        ldq_3_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_3_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_3_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_3_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_3_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_3_bits_addr_bits <= casez_tmp_202;
        else
          ldq_3_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_3_bits_addr_bits <= _GEN_280;
      ldq_3_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_3_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2649) begin
      if (_exe_tlb_uop_T_2)
        ldq_3_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_3_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_3_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_3_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_3_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_3_bits_addr_bits <= casez_tmp_202;
        else
          ldq_3_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_3_bits_addr_bits <= _GEN_274;
      ldq_3_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_3_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2268)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2073)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1784)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1592)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_3_bits_addr_valid <= ~_GEN_5749 & _GEN_5624 & _GEN_5561 & _GEN_5466 & (_GEN_5336 ? ~_GEN_5243 & _GEN_2749 : ~_GEN_5339 & _GEN_2749);
    ldq_3_bits_executed <= ~_GEN_5749 & _GEN_5624 & _GEN_5561 & _GEN_5466 & _GEN_5371 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1477) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1438)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_338 & _GEN_5048 : ~(_GEN_1425 & _GEN_338) & _GEN_5048) : _GEN_5048) | (dis_ld_val_3 ? ~_GEN_2177 & _GEN_1848 : ~_GEN_2073 & _GEN_1848));
    ldq_3_bits_succeeded <= _GEN_5624 & _GEN_5561 & _GEN_5466 & _GEN_5371 & (_GEN_5151 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h3 ? _ldq_bits_succeeded_T_1 : _GEN_5086 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h3 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2177 & _GEN_1880 : ~_GEN_2073 & _GEN_1880) : casez_tmp_490) : casez_tmp_524);
    ldq_3_bits_order_fail <= _GEN_5624 & _GEN_5561 & _GEN_5466 & _GEN_5371 & (_GEN_426 ? _GEN_2935 : _GEN_428 ? _GEN_429 | _GEN_2935 : _GEN_431 | _GEN_2935);
    ldq_3_bits_observed <= _GEN_426 | _GEN_413 | (dis_ld_val_3 ? ~_GEN_2177 & _GEN_1944 : ~_GEN_2073 & _GEN_1944);
    ldq_3_bits_forward_std_val <= _GEN_5624 & _GEN_5561 & _GEN_5466 & _GEN_5371 & (~_GEN_1508 & _GEN_5150 | ~_GEN_1468 & _GEN_5085 | (dis_ld_val_3 ? ~_GEN_2177 & _GEN_1976 : ~_GEN_2073 & _GEN_1976));
    if (_GEN_5151) begin
      if (_GEN_5086) begin
      end
      else
        ldq_3_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_3_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_4_valid <= ~_GEN_5749 & _GEN_5625 & _GEN_5562 & _GEN_5467 & (_GEN_5336 ? ~_GEN_5244 & _GEN_2181 : ~_GEN_5340 & _GEN_2181);
    if (_GEN_2270) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_4_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_4_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_4_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_4_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_4_bits_st_dep_mask <= _GEN_2166;
      ldq_4_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2074) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_4_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_4_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_4_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_4_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_4_bits_st_dep_mask <= _GEN_2069;
      ldq_4_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1785) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_4_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_4_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_4_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_4_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_4_bits_st_dep_mask <= _GEN_1685;
      ldq_4_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1593) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_4_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_4_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_4_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_4_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_4_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_4_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_4_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_4_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_4_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_4_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_4_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_4_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_4_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_4_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_4_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_4_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_4_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_4_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_4_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_4_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_4_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_4_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_4_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_4_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_4_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_4_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_4_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_4_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_4_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_4_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_4_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_4_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_4_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_4_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_4_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_4_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_4_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_4_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_4_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_4_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_4_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_4_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_4_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_4_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_4_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_4_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_4_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_4_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_4_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_4_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_4_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_4_bits_st_dep_mask <= next_live_store_mask;
      ldq_4_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_4_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_4_bits_st_dep_mask;
    if (ldq_4_valid)
      ldq_4_bits_uop_br_mask <= ldq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2270)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2074)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1785)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1593)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2750) begin
      if (_exe_tlb_uop_T_9)
        ldq_4_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_4_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_4_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_4_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_4_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_4_bits_addr_bits <= casez_tmp_202;
        else
          ldq_4_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_4_bits_addr_bits <= _GEN_280;
      ldq_4_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_4_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2650) begin
      if (_exe_tlb_uop_T_2)
        ldq_4_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_4_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_4_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_4_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_4_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_4_bits_addr_bits <= casez_tmp_202;
        else
          ldq_4_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_4_bits_addr_bits <= _GEN_274;
      ldq_4_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_4_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2270)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2074)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1785)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1593)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_4_bits_addr_valid <= ~_GEN_5749 & _GEN_5625 & _GEN_5562 & _GEN_5467 & (_GEN_5336 ? ~_GEN_5244 & _GEN_2751 : ~_GEN_5340 & _GEN_2751);
    ldq_4_bits_executed <= ~_GEN_5749 & _GEN_5625 & _GEN_5562 & _GEN_5467 & _GEN_5372 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1478) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1439)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_339 & _GEN_5049 : ~(_GEN_1425 & _GEN_339) & _GEN_5049) : _GEN_5049) | (dis_ld_val_3 ? ~_GEN_2180 & _GEN_1849 : ~_GEN_2074 & _GEN_1849));
    ldq_4_bits_succeeded <= _GEN_5625 & _GEN_5562 & _GEN_5467 & _GEN_5372 & (_GEN_5153 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h4 ? _ldq_bits_succeeded_T_1 : _GEN_5088 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h4 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2180 & _GEN_1881 : ~_GEN_2074 & _GEN_1881) : casez_tmp_490) : casez_tmp_524);
    ldq_4_bits_order_fail <= _GEN_5625 & _GEN_5562 & _GEN_5467 & _GEN_5372 & (_GEN_449 ? _GEN_2936 : _GEN_451 ? _GEN_452 | _GEN_2936 : _GEN_454 | _GEN_2936);
    ldq_4_bits_observed <= _GEN_449 | _GEN_436 | (dis_ld_val_3 ? ~_GEN_2180 & _GEN_1945 : ~_GEN_2074 & _GEN_1945);
    ldq_4_bits_forward_std_val <= _GEN_5625 & _GEN_5562 & _GEN_5467 & _GEN_5372 & (~_GEN_1508 & _GEN_5152 | ~_GEN_1468 & _GEN_5087 | (dis_ld_val_3 ? ~_GEN_2180 & _GEN_1977 : ~_GEN_2074 & _GEN_1977));
    if (_GEN_5153) begin
      if (_GEN_5088) begin
      end
      else
        ldq_4_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_4_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_5_valid <= ~_GEN_5749 & _GEN_5626 & _GEN_5563 & _GEN_5468 & (_GEN_5336 ? ~_GEN_5245 & _GEN_2184 : ~_GEN_5341 & _GEN_2184);
    if (_GEN_2272) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_5_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_5_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_5_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_5_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_5_bits_st_dep_mask <= _GEN_2166;
      ldq_5_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2075) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_5_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_5_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_5_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_5_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_5_bits_st_dep_mask <= _GEN_2069;
      ldq_5_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1786) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_5_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_5_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_5_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_5_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_5_bits_st_dep_mask <= _GEN_1685;
      ldq_5_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1594) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_5_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_5_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_5_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_5_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_5_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_5_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_5_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_5_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_5_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_5_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_5_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_5_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_5_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_5_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_5_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_5_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_5_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_5_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_5_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_5_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_5_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_5_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_5_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_5_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_5_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_5_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_5_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_5_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_5_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_5_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_5_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_5_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_5_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_5_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_5_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_5_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_5_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_5_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_5_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_5_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_5_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_5_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_5_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_5_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_5_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_5_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_5_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_5_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_5_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_5_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_5_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_5_bits_st_dep_mask <= next_live_store_mask;
      ldq_5_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_5_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_5_bits_st_dep_mask;
    if (ldq_5_valid)
      ldq_5_bits_uop_br_mask <= ldq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2272)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2075)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1786)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1594)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2752) begin
      if (_exe_tlb_uop_T_9)
        ldq_5_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_5_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_5_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_5_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_5_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_5_bits_addr_bits <= casez_tmp_202;
        else
          ldq_5_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_5_bits_addr_bits <= _GEN_280;
      ldq_5_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_5_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2651) begin
      if (_exe_tlb_uop_T_2)
        ldq_5_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_5_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_5_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_5_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_5_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_5_bits_addr_bits <= casez_tmp_202;
        else
          ldq_5_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_5_bits_addr_bits <= _GEN_274;
      ldq_5_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_5_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2272)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2075)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1786)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1594)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_5_bits_addr_valid <= ~_GEN_5749 & _GEN_5626 & _GEN_5563 & _GEN_5468 & (_GEN_5336 ? ~_GEN_5245 & _GEN_2753 : ~_GEN_5341 & _GEN_2753);
    ldq_5_bits_executed <= ~_GEN_5749 & _GEN_5626 & _GEN_5563 & _GEN_5468 & _GEN_5373 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1479) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1440)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_340 & _GEN_5050 : ~(_GEN_1425 & _GEN_340) & _GEN_5050) : _GEN_5050) | (dis_ld_val_3 ? ~_GEN_2183 & _GEN_1850 : ~_GEN_2075 & _GEN_1850));
    ldq_5_bits_succeeded <= _GEN_5626 & _GEN_5563 & _GEN_5468 & _GEN_5373 & (_GEN_5155 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h5 ? _ldq_bits_succeeded_T_1 : _GEN_5090 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h5 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2183 & _GEN_1882 : ~_GEN_2075 & _GEN_1882) : casez_tmp_490) : casez_tmp_524);
    ldq_5_bits_order_fail <= _GEN_5626 & _GEN_5563 & _GEN_5468 & _GEN_5373 & (_GEN_472 ? _GEN_2937 : _GEN_474 ? _GEN_475 | _GEN_2937 : _GEN_477 | _GEN_2937);
    ldq_5_bits_observed <= _GEN_472 | _GEN_459 | (dis_ld_val_3 ? ~_GEN_2183 & _GEN_1946 : ~_GEN_2075 & _GEN_1946);
    ldq_5_bits_forward_std_val <= _GEN_5626 & _GEN_5563 & _GEN_5468 & _GEN_5373 & (~_GEN_1508 & _GEN_5154 | ~_GEN_1468 & _GEN_5089 | (dis_ld_val_3 ? ~_GEN_2183 & _GEN_1978 : ~_GEN_2075 & _GEN_1978));
    if (_GEN_5155) begin
      if (_GEN_5090) begin
      end
      else
        ldq_5_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_5_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_6_valid <= ~_GEN_5749 & _GEN_5627 & _GEN_5564 & _GEN_5469 & (_GEN_5336 ? ~_GEN_5246 & _GEN_2187 : ~_GEN_5342 & _GEN_2187);
    if (_GEN_2274) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_6_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_6_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_6_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_6_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_6_bits_st_dep_mask <= _GEN_2166;
      ldq_6_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2076) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_6_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_6_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_6_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_6_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_6_bits_st_dep_mask <= _GEN_2069;
      ldq_6_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1787) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_6_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_6_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_6_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_6_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_6_bits_st_dep_mask <= _GEN_1685;
      ldq_6_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1595) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_6_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_6_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_6_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_6_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_6_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_6_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_6_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_6_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_6_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_6_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_6_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_6_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_6_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_6_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_6_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_6_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_6_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_6_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_6_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_6_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_6_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_6_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_6_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_6_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_6_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_6_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_6_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_6_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_6_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_6_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_6_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_6_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_6_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_6_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_6_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_6_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_6_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_6_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_6_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_6_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_6_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_6_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_6_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_6_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_6_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_6_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_6_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_6_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_6_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_6_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_6_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_6_bits_st_dep_mask <= next_live_store_mask;
      ldq_6_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_6_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_6_bits_st_dep_mask;
    if (ldq_6_valid)
      ldq_6_bits_uop_br_mask <= ldq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2274)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2076)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1787)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1595)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2754) begin
      if (_exe_tlb_uop_T_9)
        ldq_6_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_6_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_6_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_6_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_6_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_6_bits_addr_bits <= casez_tmp_202;
        else
          ldq_6_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_6_bits_addr_bits <= _GEN_280;
      ldq_6_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_6_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2652) begin
      if (_exe_tlb_uop_T_2)
        ldq_6_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_6_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_6_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_6_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_6_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_6_bits_addr_bits <= casez_tmp_202;
        else
          ldq_6_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_6_bits_addr_bits <= _GEN_274;
      ldq_6_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_6_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2274)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2076)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1787)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1595)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_6_bits_addr_valid <= ~_GEN_5749 & _GEN_5627 & _GEN_5564 & _GEN_5469 & (_GEN_5336 ? ~_GEN_5246 & _GEN_2755 : ~_GEN_5342 & _GEN_2755);
    ldq_6_bits_executed <= ~_GEN_5749 & _GEN_5627 & _GEN_5564 & _GEN_5469 & _GEN_5374 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1480) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1441)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_341 & _GEN_5051 : ~(_GEN_1425 & _GEN_341) & _GEN_5051) : _GEN_5051) | (dis_ld_val_3 ? ~_GEN_2186 & _GEN_1851 : ~_GEN_2076 & _GEN_1851));
    ldq_6_bits_succeeded <= _GEN_5627 & _GEN_5564 & _GEN_5469 & _GEN_5374 & (_GEN_5157 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h6 ? _ldq_bits_succeeded_T_1 : _GEN_5092 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h6 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2186 & _GEN_1883 : ~_GEN_2076 & _GEN_1883) : casez_tmp_490) : casez_tmp_524);
    ldq_6_bits_order_fail <= _GEN_5627 & _GEN_5564 & _GEN_5469 & _GEN_5374 & (_GEN_495 ? _GEN_2938 : _GEN_497 ? _GEN_498 | _GEN_2938 : _GEN_500 | _GEN_2938);
    ldq_6_bits_observed <= _GEN_495 | _GEN_482 | (dis_ld_val_3 ? ~_GEN_2186 & _GEN_1947 : ~_GEN_2076 & _GEN_1947);
    ldq_6_bits_forward_std_val <= _GEN_5627 & _GEN_5564 & _GEN_5469 & _GEN_5374 & (~_GEN_1508 & _GEN_5156 | ~_GEN_1468 & _GEN_5091 | (dis_ld_val_3 ? ~_GEN_2186 & _GEN_1979 : ~_GEN_2076 & _GEN_1979));
    if (_GEN_5157) begin
      if (_GEN_5092) begin
      end
      else
        ldq_6_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_6_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_7_valid <= ~_GEN_5749 & _GEN_5628 & _GEN_5565 & _GEN_5470 & (_GEN_5336 ? ~_GEN_5247 & _GEN_2190 : ~_GEN_5343 & _GEN_2190);
    if (_GEN_2276) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_7_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_7_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_7_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_7_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_7_bits_st_dep_mask <= _GEN_2166;
      ldq_7_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2077) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_7_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_7_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_7_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_7_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_7_bits_st_dep_mask <= _GEN_2069;
      ldq_7_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1788) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_7_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_7_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_7_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_7_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_7_bits_st_dep_mask <= _GEN_1685;
      ldq_7_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1596) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_7_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_7_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_7_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_7_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_7_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_7_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_7_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_7_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_7_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_7_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_7_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_7_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_7_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_7_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_7_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_7_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_7_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_7_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_7_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_7_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_7_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_7_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_7_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_7_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_7_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_7_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_7_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_7_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_7_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_7_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_7_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_7_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_7_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_7_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_7_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_7_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_7_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_7_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_7_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_7_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_7_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_7_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_7_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_7_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_7_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_7_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_7_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_7_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_7_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_7_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_7_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_7_bits_st_dep_mask <= next_live_store_mask;
      ldq_7_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_7_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_7_bits_st_dep_mask;
    if (ldq_7_valid)
      ldq_7_bits_uop_br_mask <= ldq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2276)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2077)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1788)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1596)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2756) begin
      if (_exe_tlb_uop_T_9)
        ldq_7_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_7_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_7_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_7_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_7_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_7_bits_addr_bits <= casez_tmp_202;
        else
          ldq_7_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_7_bits_addr_bits <= _GEN_280;
      ldq_7_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_7_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2653) begin
      if (_exe_tlb_uop_T_2)
        ldq_7_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_7_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_7_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_7_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_7_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_7_bits_addr_bits <= casez_tmp_202;
        else
          ldq_7_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_7_bits_addr_bits <= _GEN_274;
      ldq_7_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_7_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2276)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2077)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1788)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1596)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_7_bits_addr_valid <= ~_GEN_5749 & _GEN_5628 & _GEN_5565 & _GEN_5470 & (_GEN_5336 ? ~_GEN_5247 & _GEN_2757 : ~_GEN_5343 & _GEN_2757);
    ldq_7_bits_executed <= ~_GEN_5749 & _GEN_5628 & _GEN_5565 & _GEN_5470 & _GEN_5375 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1481) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1442)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_342 & _GEN_5052 : ~(_GEN_1425 & _GEN_342) & _GEN_5052) : _GEN_5052) | (dis_ld_val_3 ? ~_GEN_2189 & _GEN_1852 : ~_GEN_2077 & _GEN_1852));
    ldq_7_bits_succeeded <= _GEN_5628 & _GEN_5565 & _GEN_5470 & _GEN_5375 & (_GEN_5159 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h7 ? _ldq_bits_succeeded_T_1 : _GEN_5094 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h7 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2189 & _GEN_1884 : ~_GEN_2077 & _GEN_1884) : casez_tmp_490) : casez_tmp_524);
    ldq_7_bits_order_fail <= _GEN_5628 & _GEN_5565 & _GEN_5470 & _GEN_5375 & (_GEN_518 ? _GEN_2939 : _GEN_520 ? _GEN_521 | _GEN_2939 : _GEN_523 | _GEN_2939);
    ldq_7_bits_observed <= _GEN_518 | _GEN_505 | (dis_ld_val_3 ? ~_GEN_2189 & _GEN_1948 : ~_GEN_2077 & _GEN_1948);
    ldq_7_bits_forward_std_val <= _GEN_5628 & _GEN_5565 & _GEN_5470 & _GEN_5375 & (~_GEN_1508 & _GEN_5158 | ~_GEN_1468 & _GEN_5093 | (dis_ld_val_3 ? ~_GEN_2189 & _GEN_1980 : ~_GEN_2077 & _GEN_1980));
    if (_GEN_5159) begin
      if (_GEN_5094) begin
      end
      else
        ldq_7_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_7_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_8_valid <= ~_GEN_5749 & _GEN_5629 & _GEN_5566 & _GEN_5471 & (_GEN_5336 ? ~_GEN_5248 & _GEN_2193 : ~_GEN_5344 & _GEN_2193);
    if (_GEN_2278) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_8_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_8_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_8_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_8_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_8_bits_st_dep_mask <= _GEN_2166;
      ldq_8_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2078) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_8_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_8_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_8_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_8_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_8_bits_st_dep_mask <= _GEN_2069;
      ldq_8_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1789) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_8_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_8_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_8_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_8_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_8_bits_st_dep_mask <= _GEN_1685;
      ldq_8_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1597) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_8_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_8_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_8_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_8_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_8_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_8_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_8_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_8_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_8_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_8_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_8_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_8_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_8_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_8_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_8_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_8_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_8_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_8_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_8_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_8_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_8_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_8_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_8_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_8_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_8_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_8_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_8_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_8_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_8_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_8_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_8_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_8_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_8_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_8_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_8_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_8_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_8_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_8_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_8_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_8_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_8_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_8_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_8_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_8_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_8_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_8_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_8_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_8_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_8_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_8_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_8_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_8_bits_st_dep_mask <= next_live_store_mask;
      ldq_8_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_8_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_8_bits_st_dep_mask;
    if (ldq_8_valid)
      ldq_8_bits_uop_br_mask <= ldq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2278)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2078)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1789)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1597)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2758) begin
      if (_exe_tlb_uop_T_9)
        ldq_8_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_8_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_8_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_8_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_8_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_8_bits_addr_bits <= casez_tmp_202;
        else
          ldq_8_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_8_bits_addr_bits <= _GEN_280;
      ldq_8_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_8_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2654) begin
      if (_exe_tlb_uop_T_2)
        ldq_8_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_8_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_8_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_8_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_8_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_8_bits_addr_bits <= casez_tmp_202;
        else
          ldq_8_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_8_bits_addr_bits <= _GEN_274;
      ldq_8_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_8_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2278)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2078)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1789)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1597)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_8_bits_addr_valid <= ~_GEN_5749 & _GEN_5629 & _GEN_5566 & _GEN_5471 & (_GEN_5336 ? ~_GEN_5248 & _GEN_2759 : ~_GEN_5344 & _GEN_2759);
    ldq_8_bits_executed <= ~_GEN_5749 & _GEN_5629 & _GEN_5566 & _GEN_5471 & _GEN_5376 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1482) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1443)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_343 & _GEN_5053 : ~(_GEN_1425 & _GEN_343) & _GEN_5053) : _GEN_5053) | (dis_ld_val_3 ? ~_GEN_2192 & _GEN_1853 : ~_GEN_2078 & _GEN_1853));
    ldq_8_bits_succeeded <= _GEN_5629 & _GEN_5566 & _GEN_5471 & _GEN_5376 & (_GEN_5161 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h8 ? _ldq_bits_succeeded_T_1 : _GEN_5096 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h8 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2192 & _GEN_1885 : ~_GEN_2078 & _GEN_1885) : casez_tmp_490) : casez_tmp_524);
    ldq_8_bits_order_fail <= _GEN_5629 & _GEN_5566 & _GEN_5471 & _GEN_5376 & (_GEN_541 ? _GEN_2940 : _GEN_543 ? _GEN_544 | _GEN_2940 : _GEN_546 | _GEN_2940);
    ldq_8_bits_observed <= _GEN_541 | _GEN_528 | (dis_ld_val_3 ? ~_GEN_2192 & _GEN_1949 : ~_GEN_2078 & _GEN_1949);
    ldq_8_bits_forward_std_val <= _GEN_5629 & _GEN_5566 & _GEN_5471 & _GEN_5376 & (~_GEN_1508 & _GEN_5160 | ~_GEN_1468 & _GEN_5095 | (dis_ld_val_3 ? ~_GEN_2192 & _GEN_1981 : ~_GEN_2078 & _GEN_1981));
    if (_GEN_5161) begin
      if (_GEN_5096) begin
      end
      else
        ldq_8_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_8_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_9_valid <= ~_GEN_5749 & _GEN_5630 & _GEN_5567 & _GEN_5472 & (_GEN_5336 ? ~_GEN_5249 & _GEN_2196 : ~_GEN_5345 & _GEN_2196);
    if (_GEN_2280) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_9_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_9_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_9_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_9_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_9_bits_st_dep_mask <= _GEN_2166;
      ldq_9_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2079) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_9_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_9_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_9_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_9_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_9_bits_st_dep_mask <= _GEN_2069;
      ldq_9_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1790) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_9_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_9_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_9_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_9_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_9_bits_st_dep_mask <= _GEN_1685;
      ldq_9_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1598) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_9_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_9_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_9_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_9_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_9_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_9_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_9_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_9_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_9_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_9_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_9_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_9_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_9_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_9_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_9_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_9_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_9_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_9_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_9_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_9_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_9_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_9_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_9_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_9_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_9_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_9_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_9_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_9_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_9_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_9_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_9_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_9_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_9_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_9_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_9_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_9_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_9_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_9_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_9_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_9_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_9_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_9_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_9_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_9_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_9_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_9_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_9_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_9_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_9_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_9_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_9_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_9_bits_st_dep_mask <= next_live_store_mask;
      ldq_9_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_9_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_9_bits_st_dep_mask;
    if (ldq_9_valid)
      ldq_9_bits_uop_br_mask <= ldq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2280)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2079)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1790)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1598)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2760) begin
      if (_exe_tlb_uop_T_9)
        ldq_9_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_9_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_9_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_9_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_9_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_9_bits_addr_bits <= casez_tmp_202;
        else
          ldq_9_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_9_bits_addr_bits <= _GEN_280;
      ldq_9_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_9_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2655) begin
      if (_exe_tlb_uop_T_2)
        ldq_9_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_9_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_9_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_9_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_9_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_9_bits_addr_bits <= casez_tmp_202;
        else
          ldq_9_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_9_bits_addr_bits <= _GEN_274;
      ldq_9_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_9_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2280)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2079)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1790)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1598)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_9_bits_addr_valid <= ~_GEN_5749 & _GEN_5630 & _GEN_5567 & _GEN_5472 & (_GEN_5336 ? ~_GEN_5249 & _GEN_2761 : ~_GEN_5345 & _GEN_2761);
    ldq_9_bits_executed <= ~_GEN_5749 & _GEN_5630 & _GEN_5567 & _GEN_5472 & _GEN_5377 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1483) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1444)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_344 & _GEN_5054 : ~(_GEN_1425 & _GEN_344) & _GEN_5054) : _GEN_5054) | (dis_ld_val_3 ? ~_GEN_2195 & _GEN_1854 : ~_GEN_2079 & _GEN_1854));
    ldq_9_bits_succeeded <= _GEN_5630 & _GEN_5567 & _GEN_5472 & _GEN_5377 & (_GEN_5163 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h9 ? _ldq_bits_succeeded_T_1 : _GEN_5098 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h9 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2195 & _GEN_1886 : ~_GEN_2079 & _GEN_1886) : casez_tmp_490) : casez_tmp_524);
    ldq_9_bits_order_fail <= _GEN_5630 & _GEN_5567 & _GEN_5472 & _GEN_5377 & (_GEN_564 ? _GEN_2941 : _GEN_566 ? _GEN_567 | _GEN_2941 : _GEN_569 | _GEN_2941);
    ldq_9_bits_observed <= _GEN_564 | _GEN_551 | (dis_ld_val_3 ? ~_GEN_2195 & _GEN_1950 : ~_GEN_2079 & _GEN_1950);
    ldq_9_bits_forward_std_val <= _GEN_5630 & _GEN_5567 & _GEN_5472 & _GEN_5377 & (~_GEN_1508 & _GEN_5162 | ~_GEN_1468 & _GEN_5097 | (dis_ld_val_3 ? ~_GEN_2195 & _GEN_1982 : ~_GEN_2079 & _GEN_1982));
    if (_GEN_5163) begin
      if (_GEN_5098) begin
      end
      else
        ldq_9_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_9_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_10_valid <= ~_GEN_5749 & _GEN_5631 & _GEN_5568 & _GEN_5473 & (_GEN_5336 ? ~_GEN_5250 & _GEN_2199 : ~_GEN_5346 & _GEN_2199);
    if (_GEN_2282) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_10_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_10_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_10_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_10_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_10_bits_st_dep_mask <= _GEN_2166;
      ldq_10_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2080) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_10_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_10_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_10_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_10_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_10_bits_st_dep_mask <= _GEN_2069;
      ldq_10_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1791) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_10_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_10_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_10_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_10_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_10_bits_st_dep_mask <= _GEN_1685;
      ldq_10_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1599) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_10_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_10_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_10_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_10_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_10_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_10_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_10_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_10_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_10_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_10_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_10_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_10_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_10_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_10_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_10_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_10_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_10_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_10_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_10_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_10_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_10_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_10_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_10_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_10_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_10_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_10_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_10_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_10_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_10_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_10_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_10_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_10_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_10_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_10_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_10_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_10_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_10_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_10_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_10_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_10_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_10_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_10_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_10_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_10_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_10_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_10_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_10_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_10_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_10_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_10_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_10_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_10_bits_st_dep_mask <= next_live_store_mask;
      ldq_10_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_10_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_10_bits_st_dep_mask;
    if (ldq_10_valid)
      ldq_10_bits_uop_br_mask <= ldq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2282)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2080)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1791)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1599)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2762) begin
      if (_exe_tlb_uop_T_9)
        ldq_10_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_10_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_10_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_10_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_10_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_10_bits_addr_bits <= casez_tmp_202;
        else
          ldq_10_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_10_bits_addr_bits <= _GEN_280;
      ldq_10_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_10_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2656) begin
      if (_exe_tlb_uop_T_2)
        ldq_10_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_10_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_10_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_10_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_10_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_10_bits_addr_bits <= casez_tmp_202;
        else
          ldq_10_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_10_bits_addr_bits <= _GEN_274;
      ldq_10_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_10_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2282)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2080)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1791)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1599)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_10_bits_addr_valid <= ~_GEN_5749 & _GEN_5631 & _GEN_5568 & _GEN_5473 & (_GEN_5336 ? ~_GEN_5250 & _GEN_2763 : ~_GEN_5346 & _GEN_2763);
    ldq_10_bits_executed <= ~_GEN_5749 & _GEN_5631 & _GEN_5568 & _GEN_5473 & _GEN_5378 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1484) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1445)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_345 & _GEN_5055 : ~(_GEN_1425 & _GEN_345) & _GEN_5055) : _GEN_5055) | (dis_ld_val_3 ? ~_GEN_2198 & _GEN_1855 : ~_GEN_2080 & _GEN_1855));
    ldq_10_bits_succeeded <= _GEN_5631 & _GEN_5568 & _GEN_5473 & _GEN_5378 & (_GEN_5165 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hA ? _ldq_bits_succeeded_T_1 : _GEN_5100 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hA ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2198 & _GEN_1887 : ~_GEN_2080 & _GEN_1887) : casez_tmp_490) : casez_tmp_524);
    ldq_10_bits_order_fail <= _GEN_5631 & _GEN_5568 & _GEN_5473 & _GEN_5378 & (_GEN_587 ? _GEN_2942 : _GEN_589 ? _GEN_590 | _GEN_2942 : _GEN_592 | _GEN_2942);
    ldq_10_bits_observed <= _GEN_587 | _GEN_574 | (dis_ld_val_3 ? ~_GEN_2198 & _GEN_1951 : ~_GEN_2080 & _GEN_1951);
    ldq_10_bits_forward_std_val <= _GEN_5631 & _GEN_5568 & _GEN_5473 & _GEN_5378 & (~_GEN_1508 & _GEN_5164 | ~_GEN_1468 & _GEN_5099 | (dis_ld_val_3 ? ~_GEN_2198 & _GEN_1983 : ~_GEN_2080 & _GEN_1983));
    if (_GEN_5165) begin
      if (_GEN_5100) begin
      end
      else
        ldq_10_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_10_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_11_valid <= ~_GEN_5749 & _GEN_5632 & _GEN_5569 & _GEN_5474 & (_GEN_5336 ? ~_GEN_5251 & _GEN_2202 : ~_GEN_5347 & _GEN_2202);
    if (_GEN_2284) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_11_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_11_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_11_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_11_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_11_bits_st_dep_mask <= _GEN_2166;
      ldq_11_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2081) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_11_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_11_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_11_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_11_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_11_bits_st_dep_mask <= _GEN_2069;
      ldq_11_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1792) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_11_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_11_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_11_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_11_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_11_bits_st_dep_mask <= _GEN_1685;
      ldq_11_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1600) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_11_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_11_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_11_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_11_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_11_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_11_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_11_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_11_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_11_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_11_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_11_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_11_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_11_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_11_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_11_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_11_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_11_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_11_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_11_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_11_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_11_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_11_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_11_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_11_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_11_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_11_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_11_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_11_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_11_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_11_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_11_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_11_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_11_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_11_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_11_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_11_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_11_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_11_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_11_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_11_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_11_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_11_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_11_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_11_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_11_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_11_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_11_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_11_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_11_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_11_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_11_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_11_bits_st_dep_mask <= next_live_store_mask;
      ldq_11_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_11_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_11_bits_st_dep_mask;
    if (ldq_11_valid)
      ldq_11_bits_uop_br_mask <= ldq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2284)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2081)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1792)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1600)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2764) begin
      if (_exe_tlb_uop_T_9)
        ldq_11_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_11_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_11_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_11_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_11_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_11_bits_addr_bits <= casez_tmp_202;
        else
          ldq_11_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_11_bits_addr_bits <= _GEN_280;
      ldq_11_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_11_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2657) begin
      if (_exe_tlb_uop_T_2)
        ldq_11_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_11_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_11_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_11_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_11_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_11_bits_addr_bits <= casez_tmp_202;
        else
          ldq_11_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_11_bits_addr_bits <= _GEN_274;
      ldq_11_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_11_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2284)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2081)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1792)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1600)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_11_bits_addr_valid <= ~_GEN_5749 & _GEN_5632 & _GEN_5569 & _GEN_5474 & (_GEN_5336 ? ~_GEN_5251 & _GEN_2765 : ~_GEN_5347 & _GEN_2765);
    ldq_11_bits_executed <= ~_GEN_5749 & _GEN_5632 & _GEN_5569 & _GEN_5474 & _GEN_5379 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1485) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1446)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_346 & _GEN_5056 : ~(_GEN_1425 & _GEN_346) & _GEN_5056) : _GEN_5056) | (dis_ld_val_3 ? ~_GEN_2201 & _GEN_1856 : ~_GEN_2081 & _GEN_1856));
    ldq_11_bits_succeeded <= _GEN_5632 & _GEN_5569 & _GEN_5474 & _GEN_5379 & (_GEN_5167 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hB ? _ldq_bits_succeeded_T_1 : _GEN_5102 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hB ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2201 & _GEN_1888 : ~_GEN_2081 & _GEN_1888) : casez_tmp_490) : casez_tmp_524);
    ldq_11_bits_order_fail <= _GEN_5632 & _GEN_5569 & _GEN_5474 & _GEN_5379 & (_GEN_610 ? _GEN_2943 : _GEN_612 ? _GEN_613 | _GEN_2943 : _GEN_615 | _GEN_2943);
    ldq_11_bits_observed <= _GEN_610 | _GEN_597 | (dis_ld_val_3 ? ~_GEN_2201 & _GEN_1952 : ~_GEN_2081 & _GEN_1952);
    ldq_11_bits_forward_std_val <= _GEN_5632 & _GEN_5569 & _GEN_5474 & _GEN_5379 & (~_GEN_1508 & _GEN_5166 | ~_GEN_1468 & _GEN_5101 | (dis_ld_val_3 ? ~_GEN_2201 & _GEN_1984 : ~_GEN_2081 & _GEN_1984));
    if (_GEN_5167) begin
      if (_GEN_5102) begin
      end
      else
        ldq_11_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_11_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_12_valid <= ~_GEN_5749 & _GEN_5633 & _GEN_5570 & _GEN_5475 & (_GEN_5336 ? ~_GEN_5252 & _GEN_2205 : ~_GEN_5348 & _GEN_2205);
    if (_GEN_2286) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_12_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_12_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_12_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_12_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_12_bits_st_dep_mask <= _GEN_2166;
      ldq_12_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2082) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_12_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_12_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_12_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_12_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_12_bits_st_dep_mask <= _GEN_2069;
      ldq_12_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1793) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_12_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_12_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_12_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_12_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_12_bits_st_dep_mask <= _GEN_1685;
      ldq_12_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1601) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_12_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_12_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_12_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_12_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_12_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_12_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_12_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_12_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_12_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_12_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_12_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_12_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_12_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_12_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_12_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_12_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_12_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_12_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_12_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_12_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_12_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_12_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_12_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_12_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_12_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_12_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_12_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_12_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_12_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_12_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_12_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_12_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_12_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_12_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_12_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_12_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_12_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_12_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_12_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_12_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_12_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_12_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_12_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_12_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_12_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_12_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_12_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_12_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_12_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_12_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_12_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_12_bits_st_dep_mask <= next_live_store_mask;
      ldq_12_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_12_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_12_bits_st_dep_mask;
    if (ldq_12_valid)
      ldq_12_bits_uop_br_mask <= ldq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2286)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2082)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1793)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1601)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2766) begin
      if (_exe_tlb_uop_T_9)
        ldq_12_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_12_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_12_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_12_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_12_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_12_bits_addr_bits <= casez_tmp_202;
        else
          ldq_12_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_12_bits_addr_bits <= _GEN_280;
      ldq_12_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_12_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2658) begin
      if (_exe_tlb_uop_T_2)
        ldq_12_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_12_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_12_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_12_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_12_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_12_bits_addr_bits <= casez_tmp_202;
        else
          ldq_12_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_12_bits_addr_bits <= _GEN_274;
      ldq_12_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_12_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2286)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2082)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1793)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1601)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_12_bits_addr_valid <= ~_GEN_5749 & _GEN_5633 & _GEN_5570 & _GEN_5475 & (_GEN_5336 ? ~_GEN_5252 & _GEN_2767 : ~_GEN_5348 & _GEN_2767);
    ldq_12_bits_executed <= ~_GEN_5749 & _GEN_5633 & _GEN_5570 & _GEN_5475 & _GEN_5380 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1486) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1447)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_347 & _GEN_5057 : ~(_GEN_1425 & _GEN_347) & _GEN_5057) : _GEN_5057) | (dis_ld_val_3 ? ~_GEN_2204 & _GEN_1857 : ~_GEN_2082 & _GEN_1857));
    ldq_12_bits_succeeded <= _GEN_5633 & _GEN_5570 & _GEN_5475 & _GEN_5380 & (_GEN_5169 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hC ? _ldq_bits_succeeded_T_1 : _GEN_5104 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hC ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2204 & _GEN_1889 : ~_GEN_2082 & _GEN_1889) : casez_tmp_490) : casez_tmp_524);
    ldq_12_bits_order_fail <= _GEN_5633 & _GEN_5570 & _GEN_5475 & _GEN_5380 & (_GEN_633 ? _GEN_2944 : _GEN_635 ? _GEN_636 | _GEN_2944 : _GEN_638 | _GEN_2944);
    ldq_12_bits_observed <= _GEN_633 | _GEN_620 | (dis_ld_val_3 ? ~_GEN_2204 & _GEN_1953 : ~_GEN_2082 & _GEN_1953);
    ldq_12_bits_forward_std_val <= _GEN_5633 & _GEN_5570 & _GEN_5475 & _GEN_5380 & (~_GEN_1508 & _GEN_5168 | ~_GEN_1468 & _GEN_5103 | (dis_ld_val_3 ? ~_GEN_2204 & _GEN_1985 : ~_GEN_2082 & _GEN_1985));
    if (_GEN_5169) begin
      if (_GEN_5104) begin
      end
      else
        ldq_12_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_12_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_13_valid <= ~_GEN_5749 & _GEN_5634 & _GEN_5571 & _GEN_5476 & (_GEN_5336 ? ~_GEN_5253 & _GEN_2208 : ~_GEN_5349 & _GEN_2208);
    if (_GEN_2288) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_13_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_13_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_13_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_13_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_13_bits_st_dep_mask <= _GEN_2166;
      ldq_13_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2083) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_13_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_13_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_13_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_13_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_13_bits_st_dep_mask <= _GEN_2069;
      ldq_13_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1794) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_13_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_13_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_13_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_13_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_13_bits_st_dep_mask <= _GEN_1685;
      ldq_13_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1602) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_13_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_13_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_13_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_13_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_13_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_13_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_13_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_13_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_13_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_13_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_13_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_13_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_13_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_13_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_13_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_13_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_13_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_13_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_13_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_13_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_13_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_13_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_13_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_13_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_13_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_13_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_13_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_13_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_13_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_13_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_13_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_13_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_13_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_13_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_13_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_13_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_13_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_13_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_13_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_13_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_13_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_13_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_13_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_13_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_13_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_13_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_13_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_13_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_13_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_13_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_13_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_13_bits_st_dep_mask <= next_live_store_mask;
      ldq_13_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_13_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_13_bits_st_dep_mask;
    if (ldq_13_valid)
      ldq_13_bits_uop_br_mask <= ldq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2288)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2083)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1794)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1602)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2768) begin
      if (_exe_tlb_uop_T_9)
        ldq_13_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_13_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_13_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_13_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_13_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_13_bits_addr_bits <= casez_tmp_202;
        else
          ldq_13_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_13_bits_addr_bits <= _GEN_280;
      ldq_13_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_13_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2659) begin
      if (_exe_tlb_uop_T_2)
        ldq_13_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_13_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_13_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_13_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_13_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_13_bits_addr_bits <= casez_tmp_202;
        else
          ldq_13_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_13_bits_addr_bits <= _GEN_274;
      ldq_13_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_13_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2288)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2083)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1794)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1602)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_13_bits_addr_valid <= ~_GEN_5749 & _GEN_5634 & _GEN_5571 & _GEN_5476 & (_GEN_5336 ? ~_GEN_5253 & _GEN_2769 : ~_GEN_5349 & _GEN_2769);
    ldq_13_bits_executed <= ~_GEN_5749 & _GEN_5634 & _GEN_5571 & _GEN_5476 & _GEN_5381 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1487) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1448)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_348 & _GEN_5058 : ~(_GEN_1425 & _GEN_348) & _GEN_5058) : _GEN_5058) | (dis_ld_val_3 ? ~_GEN_2207 & _GEN_1858 : ~_GEN_2083 & _GEN_1858));
    ldq_13_bits_succeeded <= _GEN_5634 & _GEN_5571 & _GEN_5476 & _GEN_5381 & (_GEN_5171 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hD ? _ldq_bits_succeeded_T_1 : _GEN_5106 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hD ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2207 & _GEN_1890 : ~_GEN_2083 & _GEN_1890) : casez_tmp_490) : casez_tmp_524);
    ldq_13_bits_order_fail <= _GEN_5634 & _GEN_5571 & _GEN_5476 & _GEN_5381 & (_GEN_656 ? _GEN_2945 : _GEN_658 ? _GEN_659 | _GEN_2945 : _GEN_661 | _GEN_2945);
    ldq_13_bits_observed <= _GEN_656 | _GEN_643 | (dis_ld_val_3 ? ~_GEN_2207 & _GEN_1954 : ~_GEN_2083 & _GEN_1954);
    ldq_13_bits_forward_std_val <= _GEN_5634 & _GEN_5571 & _GEN_5476 & _GEN_5381 & (~_GEN_1508 & _GEN_5170 | ~_GEN_1468 & _GEN_5105 | (dis_ld_val_3 ? ~_GEN_2207 & _GEN_1986 : ~_GEN_2083 & _GEN_1986));
    if (_GEN_5171) begin
      if (_GEN_5106) begin
      end
      else
        ldq_13_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_13_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_14_valid <= ~_GEN_5749 & _GEN_5635 & _GEN_5572 & _GEN_5477 & (_GEN_5336 ? ~_GEN_5254 & _GEN_2211 : ~_GEN_5350 & _GEN_2211);
    if (_GEN_2290) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_14_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_14_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_14_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_14_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_14_bits_st_dep_mask <= _GEN_2166;
      ldq_14_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2084) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_14_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_14_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_14_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_14_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_14_bits_st_dep_mask <= _GEN_2069;
      ldq_14_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1795) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_14_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_14_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_14_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_14_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_14_bits_st_dep_mask <= _GEN_1685;
      ldq_14_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1603) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_14_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_14_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_14_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_14_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_14_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_14_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_14_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_14_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_14_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_14_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_14_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_14_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_14_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_14_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_14_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_14_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_14_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_14_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_14_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_14_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_14_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_14_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_14_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_14_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_14_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_14_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_14_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_14_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_14_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_14_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_14_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_14_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_14_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_14_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_14_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_14_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_14_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_14_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_14_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_14_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_14_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_14_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_14_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_14_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_14_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_14_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_14_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_14_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_14_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_14_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_14_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_14_bits_st_dep_mask <= next_live_store_mask;
      ldq_14_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_14_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_14_bits_st_dep_mask;
    if (ldq_14_valid)
      ldq_14_bits_uop_br_mask <= ldq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2290)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2084)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1795)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1603)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2770) begin
      if (_exe_tlb_uop_T_9)
        ldq_14_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_14_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_14_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_14_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_14_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_14_bits_addr_bits <= casez_tmp_202;
        else
          ldq_14_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_14_bits_addr_bits <= _GEN_280;
      ldq_14_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_14_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2660) begin
      if (_exe_tlb_uop_T_2)
        ldq_14_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_14_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_14_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_14_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_14_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_14_bits_addr_bits <= casez_tmp_202;
        else
          ldq_14_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_14_bits_addr_bits <= _GEN_274;
      ldq_14_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_14_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2290)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2084)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1795)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1603)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_14_bits_addr_valid <= ~_GEN_5749 & _GEN_5635 & _GEN_5572 & _GEN_5477 & (_GEN_5336 ? ~_GEN_5254 & _GEN_2771 : ~_GEN_5350 & _GEN_2771);
    ldq_14_bits_executed <= ~_GEN_5749 & _GEN_5635 & _GEN_5572 & _GEN_5477 & _GEN_5382 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1488) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1449)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_349 & _GEN_5059 : ~(_GEN_1425 & _GEN_349) & _GEN_5059) : _GEN_5059) | (dis_ld_val_3 ? ~_GEN_2210 & _GEN_1859 : ~_GEN_2084 & _GEN_1859));
    ldq_14_bits_succeeded <= _GEN_5635 & _GEN_5572 & _GEN_5477 & _GEN_5382 & (_GEN_5173 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hE ? _ldq_bits_succeeded_T_1 : _GEN_5108 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hE ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2210 & _GEN_1891 : ~_GEN_2084 & _GEN_1891) : casez_tmp_490) : casez_tmp_524);
    ldq_14_bits_order_fail <= _GEN_5635 & _GEN_5572 & _GEN_5477 & _GEN_5382 & (_GEN_679 ? _GEN_2946 : _GEN_681 ? _GEN_682 | _GEN_2946 : _GEN_684 | _GEN_2946);
    ldq_14_bits_observed <= _GEN_679 | _GEN_666 | (dis_ld_val_3 ? ~_GEN_2210 & _GEN_1955 : ~_GEN_2084 & _GEN_1955);
    ldq_14_bits_forward_std_val <= _GEN_5635 & _GEN_5572 & _GEN_5477 & _GEN_5382 & (~_GEN_1508 & _GEN_5172 | ~_GEN_1468 & _GEN_5107 | (dis_ld_val_3 ? ~_GEN_2210 & _GEN_1987 : ~_GEN_2084 & _GEN_1987));
    if (_GEN_5173) begin
      if (_GEN_5108) begin
      end
      else
        ldq_14_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_14_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_15_valid <= ~_GEN_5749 & _GEN_5636 & _GEN_5573 & _GEN_5478 & (_GEN_5336 ? ~_GEN_5255 & _GEN_2214 : ~_GEN_5351 & _GEN_2214);
    if (_GEN_2292) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_15_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_15_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_15_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_15_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_15_bits_st_dep_mask <= _GEN_2166;
      ldq_15_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2085) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_15_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_15_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_15_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_15_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_15_bits_st_dep_mask <= _GEN_2069;
      ldq_15_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1796) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_15_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_15_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_15_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_15_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_15_bits_st_dep_mask <= _GEN_1685;
      ldq_15_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1604) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_15_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_15_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_15_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_15_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_15_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_15_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_15_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_15_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_15_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_15_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_15_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_15_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_15_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_15_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_15_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_15_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_15_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_15_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_15_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_15_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_15_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_15_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_15_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_15_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_15_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_15_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_15_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_15_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_15_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_15_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_15_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_15_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_15_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_15_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_15_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_15_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_15_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_15_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_15_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_15_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_15_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_15_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_15_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_15_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_15_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_15_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_15_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_15_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_15_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_15_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_15_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_15_bits_st_dep_mask <= next_live_store_mask;
      ldq_15_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_15_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_15_bits_st_dep_mask;
    if (ldq_15_valid)
      ldq_15_bits_uop_br_mask <= ldq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2292)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2085)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1796)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1604)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2772) begin
      if (_exe_tlb_uop_T_9)
        ldq_15_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_15_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_15_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_15_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_15_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_15_bits_addr_bits <= casez_tmp_202;
        else
          ldq_15_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_15_bits_addr_bits <= _GEN_280;
      ldq_15_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_15_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2661) begin
      if (_exe_tlb_uop_T_2)
        ldq_15_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_15_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_15_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_15_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_15_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_15_bits_addr_bits <= casez_tmp_202;
        else
          ldq_15_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_15_bits_addr_bits <= _GEN_274;
      ldq_15_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_15_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2292)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2085)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1796)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1604)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_15_bits_addr_valid <= ~_GEN_5749 & _GEN_5636 & _GEN_5573 & _GEN_5478 & (_GEN_5336 ? ~_GEN_5255 & _GEN_2773 : ~_GEN_5351 & _GEN_2773);
    ldq_15_bits_executed <= ~_GEN_5749 & _GEN_5636 & _GEN_5573 & _GEN_5478 & _GEN_5383 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1489) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1450)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_350 & _GEN_5060 : ~(_GEN_1425 & _GEN_350) & _GEN_5060) : _GEN_5060) | (dis_ld_val_3 ? ~_GEN_2213 & _GEN_1860 : ~_GEN_2085 & _GEN_1860));
    ldq_15_bits_succeeded <= _GEN_5636 & _GEN_5573 & _GEN_5478 & _GEN_5383 & (_GEN_5175 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hF ? _ldq_bits_succeeded_T_1 : _GEN_5110 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hF ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2213 & _GEN_1892 : ~_GEN_2085 & _GEN_1892) : casez_tmp_490) : casez_tmp_524);
    ldq_15_bits_order_fail <= _GEN_5636 & _GEN_5573 & _GEN_5478 & _GEN_5383 & (_GEN_702 ? _GEN_2947 : _GEN_704 ? _GEN_705 | _GEN_2947 : _GEN_707 | _GEN_2947);
    ldq_15_bits_observed <= _GEN_702 | _GEN_689 | (dis_ld_val_3 ? ~_GEN_2213 & _GEN_1956 : ~_GEN_2085 & _GEN_1956);
    ldq_15_bits_forward_std_val <= _GEN_5636 & _GEN_5573 & _GEN_5478 & _GEN_5383 & (~_GEN_1508 & _GEN_5174 | ~_GEN_1468 & _GEN_5109 | (dis_ld_val_3 ? ~_GEN_2213 & _GEN_1988 : ~_GEN_2085 & _GEN_1988));
    if (_GEN_5175) begin
      if (_GEN_5110) begin
      end
      else
        ldq_15_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_15_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_16_valid <= ~_GEN_5749 & _GEN_5637 & _GEN_5574 & _GEN_5479 & (_GEN_5336 ? ~_GEN_5256 & _GEN_2217 : ~_GEN_5352 & _GEN_2217);
    if (_GEN_2294) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_16_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_16_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_16_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_16_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_16_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_16_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_16_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_16_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_16_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_16_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_16_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_16_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_16_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_16_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_16_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_16_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_16_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_16_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_16_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_16_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_16_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_16_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_16_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_16_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_16_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_16_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_16_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_16_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_16_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_16_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_16_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_16_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_16_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_16_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_16_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_16_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_16_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_16_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_16_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_16_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_16_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_16_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_16_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_16_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_16_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_16_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_16_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_16_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_16_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_16_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_16_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_16_bits_st_dep_mask <= _GEN_2166;
      ldq_16_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2086) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_16_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_16_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_16_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_16_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_16_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_16_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_16_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_16_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_16_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_16_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_16_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_16_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_16_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_16_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_16_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_16_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_16_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_16_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_16_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_16_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_16_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_16_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_16_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_16_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_16_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_16_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_16_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_16_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_16_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_16_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_16_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_16_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_16_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_16_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_16_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_16_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_16_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_16_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_16_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_16_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_16_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_16_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_16_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_16_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_16_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_16_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_16_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_16_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_16_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_16_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_16_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_16_bits_st_dep_mask <= _GEN_2069;
      ldq_16_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1797) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_16_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_16_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_16_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_16_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_16_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_16_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_16_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_16_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_16_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_16_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_16_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_16_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_16_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_16_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_16_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_16_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_16_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_16_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_16_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_16_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_16_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_16_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_16_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_16_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_16_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_16_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_16_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_16_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_16_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_16_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_16_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_16_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_16_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_16_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_16_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_16_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_16_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_16_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_16_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_16_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_16_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_16_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_16_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_16_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_16_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_16_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_16_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_16_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_16_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_16_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_16_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_16_bits_st_dep_mask <= _GEN_1685;
      ldq_16_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1605) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_16_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_16_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_16_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_16_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_16_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_16_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_16_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_16_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_16_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_16_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_16_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_16_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_16_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_16_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_16_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_16_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_16_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_16_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_16_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_16_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_16_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_16_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_16_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_16_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_16_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_16_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_16_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_16_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_16_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_16_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_16_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_16_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_16_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_16_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_16_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_16_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_16_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_16_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_16_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_16_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_16_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_16_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_16_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_16_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_16_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_16_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_16_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_16_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_16_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_16_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_16_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_16_bits_st_dep_mask <= next_live_store_mask;
      ldq_16_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_16_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_16_bits_st_dep_mask;
    if (ldq_16_valid)
      ldq_16_bits_uop_br_mask <= ldq_16_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2294)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2086)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1797)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1605)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2774) begin
      if (_exe_tlb_uop_T_9)
        ldq_16_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_16_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_16_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_16_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_16_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_16_bits_addr_bits <= casez_tmp_202;
        else
          ldq_16_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_16_bits_addr_bits <= _GEN_280;
      ldq_16_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_16_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2662) begin
      if (_exe_tlb_uop_T_2)
        ldq_16_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_16_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_16_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_16_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_16_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_16_bits_addr_bits <= casez_tmp_202;
        else
          ldq_16_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_16_bits_addr_bits <= _GEN_274;
      ldq_16_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_16_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2294)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2086)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1797)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1605)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_16_bits_addr_valid <= ~_GEN_5749 & _GEN_5637 & _GEN_5574 & _GEN_5479 & (_GEN_5336 ? ~_GEN_5256 & _GEN_2775 : ~_GEN_5352 & _GEN_2775);
    ldq_16_bits_executed <= ~_GEN_5749 & _GEN_5637 & _GEN_5574 & _GEN_5479 & _GEN_5384 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1490) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1451)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_351 & _GEN_5061 : ~(_GEN_1425 & _GEN_351) & _GEN_5061) : _GEN_5061) | (dis_ld_val_3 ? ~_GEN_2216 & _GEN_1861 : ~_GEN_2086 & _GEN_1861));
    ldq_16_bits_succeeded <= _GEN_5637 & _GEN_5574 & _GEN_5479 & _GEN_5384 & (_GEN_5177 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h10 ? _ldq_bits_succeeded_T_1 : _GEN_5112 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h10 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2216 & _GEN_1893 : ~_GEN_2086 & _GEN_1893) : casez_tmp_490) : casez_tmp_524);
    ldq_16_bits_order_fail <= _GEN_5637 & _GEN_5574 & _GEN_5479 & _GEN_5384 & (_GEN_725 ? _GEN_2948 : _GEN_727 ? _GEN_728 | _GEN_2948 : _GEN_730 | _GEN_2948);
    ldq_16_bits_observed <= _GEN_725 | _GEN_712 | (dis_ld_val_3 ? ~_GEN_2216 & _GEN_1957 : ~_GEN_2086 & _GEN_1957);
    ldq_16_bits_forward_std_val <= _GEN_5637 & _GEN_5574 & _GEN_5479 & _GEN_5384 & (~_GEN_1508 & _GEN_5176 | ~_GEN_1468 & _GEN_5111 | (dis_ld_val_3 ? ~_GEN_2216 & _GEN_1989 : ~_GEN_2086 & _GEN_1989));
    if (_GEN_5177) begin
      if (_GEN_5112) begin
      end
      else
        ldq_16_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_16_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_17_valid <= ~_GEN_5749 & _GEN_5638 & _GEN_5575 & _GEN_5480 & (_GEN_5336 ? ~_GEN_5257 & _GEN_2220 : ~_GEN_5353 & _GEN_2220);
    if (_GEN_2296) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_17_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_17_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_17_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_17_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_17_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_17_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_17_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_17_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_17_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_17_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_17_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_17_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_17_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_17_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_17_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_17_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_17_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_17_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_17_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_17_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_17_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_17_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_17_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_17_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_17_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_17_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_17_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_17_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_17_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_17_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_17_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_17_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_17_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_17_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_17_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_17_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_17_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_17_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_17_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_17_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_17_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_17_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_17_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_17_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_17_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_17_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_17_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_17_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_17_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_17_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_17_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_17_bits_st_dep_mask <= _GEN_2166;
      ldq_17_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2087) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_17_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_17_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_17_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_17_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_17_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_17_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_17_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_17_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_17_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_17_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_17_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_17_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_17_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_17_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_17_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_17_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_17_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_17_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_17_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_17_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_17_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_17_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_17_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_17_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_17_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_17_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_17_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_17_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_17_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_17_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_17_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_17_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_17_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_17_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_17_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_17_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_17_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_17_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_17_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_17_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_17_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_17_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_17_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_17_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_17_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_17_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_17_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_17_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_17_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_17_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_17_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_17_bits_st_dep_mask <= _GEN_2069;
      ldq_17_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1798) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_17_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_17_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_17_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_17_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_17_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_17_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_17_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_17_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_17_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_17_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_17_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_17_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_17_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_17_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_17_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_17_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_17_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_17_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_17_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_17_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_17_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_17_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_17_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_17_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_17_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_17_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_17_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_17_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_17_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_17_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_17_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_17_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_17_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_17_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_17_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_17_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_17_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_17_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_17_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_17_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_17_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_17_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_17_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_17_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_17_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_17_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_17_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_17_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_17_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_17_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_17_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_17_bits_st_dep_mask <= _GEN_1685;
      ldq_17_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1606) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_17_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_17_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_17_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_17_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_17_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_17_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_17_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_17_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_17_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_17_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_17_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_17_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_17_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_17_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_17_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_17_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_17_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_17_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_17_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_17_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_17_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_17_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_17_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_17_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_17_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_17_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_17_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_17_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_17_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_17_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_17_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_17_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_17_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_17_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_17_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_17_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_17_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_17_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_17_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_17_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_17_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_17_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_17_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_17_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_17_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_17_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_17_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_17_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_17_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_17_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_17_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_17_bits_st_dep_mask <= next_live_store_mask;
      ldq_17_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_17_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_17_bits_st_dep_mask;
    if (ldq_17_valid)
      ldq_17_bits_uop_br_mask <= ldq_17_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2296)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2087)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1798)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1606)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2776) begin
      if (_exe_tlb_uop_T_9)
        ldq_17_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_17_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_17_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_17_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_17_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_17_bits_addr_bits <= casez_tmp_202;
        else
          ldq_17_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_17_bits_addr_bits <= _GEN_280;
      ldq_17_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_17_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2663) begin
      if (_exe_tlb_uop_T_2)
        ldq_17_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_17_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_17_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_17_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_17_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_17_bits_addr_bits <= casez_tmp_202;
        else
          ldq_17_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_17_bits_addr_bits <= _GEN_274;
      ldq_17_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_17_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2296)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2087)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1798)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1606)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_17_bits_addr_valid <= ~_GEN_5749 & _GEN_5638 & _GEN_5575 & _GEN_5480 & (_GEN_5336 ? ~_GEN_5257 & _GEN_2777 : ~_GEN_5353 & _GEN_2777);
    ldq_17_bits_executed <= ~_GEN_5749 & _GEN_5638 & _GEN_5575 & _GEN_5480 & _GEN_5385 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1491) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1452)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_352 & _GEN_5062 : ~(_GEN_1425 & _GEN_352) & _GEN_5062) : _GEN_5062) | (dis_ld_val_3 ? ~_GEN_2219 & _GEN_1862 : ~_GEN_2087 & _GEN_1862));
    ldq_17_bits_succeeded <= _GEN_5638 & _GEN_5575 & _GEN_5480 & _GEN_5385 & (_GEN_5179 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h11 ? _ldq_bits_succeeded_T_1 : _GEN_5114 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h11 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2219 & _GEN_1894 : ~_GEN_2087 & _GEN_1894) : casez_tmp_490) : casez_tmp_524);
    ldq_17_bits_order_fail <= _GEN_5638 & _GEN_5575 & _GEN_5480 & _GEN_5385 & (_GEN_748 ? _GEN_2949 : _GEN_750 ? _GEN_751 | _GEN_2949 : _GEN_753 | _GEN_2949);
    ldq_17_bits_observed <= _GEN_748 | _GEN_735 | (dis_ld_val_3 ? ~_GEN_2219 & _GEN_1958 : ~_GEN_2087 & _GEN_1958);
    ldq_17_bits_forward_std_val <= _GEN_5638 & _GEN_5575 & _GEN_5480 & _GEN_5385 & (~_GEN_1508 & _GEN_5178 | ~_GEN_1468 & _GEN_5113 | (dis_ld_val_3 ? ~_GEN_2219 & _GEN_1990 : ~_GEN_2087 & _GEN_1990));
    if (_GEN_5179) begin
      if (_GEN_5114) begin
      end
      else
        ldq_17_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_17_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_18_valid <= ~_GEN_5749 & _GEN_5639 & _GEN_5576 & _GEN_5481 & (_GEN_5336 ? ~_GEN_5258 & _GEN_2223 : ~_GEN_5354 & _GEN_2223);
    if (_GEN_2298) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_18_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_18_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_18_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_18_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_18_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_18_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_18_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_18_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_18_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_18_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_18_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_18_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_18_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_18_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_18_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_18_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_18_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_18_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_18_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_18_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_18_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_18_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_18_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_18_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_18_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_18_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_18_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_18_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_18_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_18_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_18_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_18_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_18_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_18_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_18_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_18_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_18_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_18_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_18_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_18_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_18_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_18_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_18_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_18_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_18_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_18_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_18_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_18_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_18_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_18_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_18_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_18_bits_st_dep_mask <= _GEN_2166;
      ldq_18_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2088) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_18_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_18_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_18_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_18_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_18_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_18_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_18_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_18_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_18_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_18_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_18_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_18_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_18_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_18_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_18_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_18_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_18_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_18_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_18_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_18_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_18_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_18_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_18_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_18_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_18_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_18_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_18_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_18_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_18_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_18_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_18_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_18_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_18_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_18_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_18_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_18_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_18_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_18_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_18_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_18_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_18_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_18_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_18_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_18_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_18_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_18_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_18_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_18_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_18_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_18_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_18_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_18_bits_st_dep_mask <= _GEN_2069;
      ldq_18_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1799) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_18_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_18_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_18_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_18_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_18_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_18_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_18_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_18_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_18_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_18_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_18_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_18_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_18_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_18_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_18_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_18_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_18_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_18_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_18_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_18_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_18_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_18_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_18_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_18_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_18_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_18_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_18_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_18_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_18_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_18_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_18_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_18_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_18_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_18_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_18_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_18_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_18_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_18_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_18_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_18_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_18_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_18_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_18_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_18_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_18_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_18_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_18_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_18_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_18_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_18_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_18_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_18_bits_st_dep_mask <= _GEN_1685;
      ldq_18_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1607) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_18_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_18_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_18_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_18_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_18_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_18_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_18_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_18_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_18_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_18_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_18_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_18_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_18_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_18_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_18_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_18_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_18_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_18_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_18_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_18_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_18_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_18_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_18_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_18_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_18_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_18_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_18_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_18_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_18_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_18_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_18_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_18_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_18_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_18_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_18_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_18_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_18_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_18_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_18_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_18_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_18_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_18_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_18_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_18_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_18_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_18_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_18_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_18_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_18_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_18_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_18_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_18_bits_st_dep_mask <= next_live_store_mask;
      ldq_18_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_18_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_18_bits_st_dep_mask;
    if (ldq_18_valid)
      ldq_18_bits_uop_br_mask <= ldq_18_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2298)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2088)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1799)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1607)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2778) begin
      if (_exe_tlb_uop_T_9)
        ldq_18_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_18_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_18_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_18_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_18_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_18_bits_addr_bits <= casez_tmp_202;
        else
          ldq_18_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_18_bits_addr_bits <= _GEN_280;
      ldq_18_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_18_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2664) begin
      if (_exe_tlb_uop_T_2)
        ldq_18_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_18_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_18_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_18_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_18_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_18_bits_addr_bits <= casez_tmp_202;
        else
          ldq_18_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_18_bits_addr_bits <= _GEN_274;
      ldq_18_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_18_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2298)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2088)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1799)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1607)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_18_bits_addr_valid <= ~_GEN_5749 & _GEN_5639 & _GEN_5576 & _GEN_5481 & (_GEN_5336 ? ~_GEN_5258 & _GEN_2779 : ~_GEN_5354 & _GEN_2779);
    ldq_18_bits_executed <= ~_GEN_5749 & _GEN_5639 & _GEN_5576 & _GEN_5481 & _GEN_5386 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1492) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1453)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_353 & _GEN_5063 : ~(_GEN_1425 & _GEN_353) & _GEN_5063) : _GEN_5063) | (dis_ld_val_3 ? ~_GEN_2222 & _GEN_1863 : ~_GEN_2088 & _GEN_1863));
    ldq_18_bits_succeeded <= _GEN_5639 & _GEN_5576 & _GEN_5481 & _GEN_5386 & (_GEN_5181 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h12 ? _ldq_bits_succeeded_T_1 : _GEN_5116 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h12 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2222 & _GEN_1895 : ~_GEN_2088 & _GEN_1895) : casez_tmp_490) : casez_tmp_524);
    ldq_18_bits_order_fail <= _GEN_5639 & _GEN_5576 & _GEN_5481 & _GEN_5386 & (_GEN_771 ? _GEN_2950 : _GEN_773 ? _GEN_774 | _GEN_2950 : _GEN_776 | _GEN_2950);
    ldq_18_bits_observed <= _GEN_771 | _GEN_758 | (dis_ld_val_3 ? ~_GEN_2222 & _GEN_1959 : ~_GEN_2088 & _GEN_1959);
    ldq_18_bits_forward_std_val <= _GEN_5639 & _GEN_5576 & _GEN_5481 & _GEN_5386 & (~_GEN_1508 & _GEN_5180 | ~_GEN_1468 & _GEN_5115 | (dis_ld_val_3 ? ~_GEN_2222 & _GEN_1991 : ~_GEN_2088 & _GEN_1991));
    if (_GEN_5181) begin
      if (_GEN_5116) begin
      end
      else
        ldq_18_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_18_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_19_valid <= ~_GEN_5749 & _GEN_5640 & _GEN_5577 & _GEN_5482 & (_GEN_5336 ? ~_GEN_5259 & _GEN_2226 : ~_GEN_5355 & _GEN_2226);
    if (_GEN_2300) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_19_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_19_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_19_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_19_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_19_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_19_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_19_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_19_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_19_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_19_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_19_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_19_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_19_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_19_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_19_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_19_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_19_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_19_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_19_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_19_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_19_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_19_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_19_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_19_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_19_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_19_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_19_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_19_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_19_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_19_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_19_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_19_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_19_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_19_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_19_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_19_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_19_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_19_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_19_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_19_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_19_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_19_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_19_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_19_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_19_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_19_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_19_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_19_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_19_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_19_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_19_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_19_bits_st_dep_mask <= _GEN_2166;
      ldq_19_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2089) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_19_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_19_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_19_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_19_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_19_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_19_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_19_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_19_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_19_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_19_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_19_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_19_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_19_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_19_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_19_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_19_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_19_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_19_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_19_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_19_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_19_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_19_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_19_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_19_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_19_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_19_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_19_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_19_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_19_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_19_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_19_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_19_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_19_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_19_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_19_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_19_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_19_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_19_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_19_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_19_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_19_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_19_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_19_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_19_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_19_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_19_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_19_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_19_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_19_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_19_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_19_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_19_bits_st_dep_mask <= _GEN_2069;
      ldq_19_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1800) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_19_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_19_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_19_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_19_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_19_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_19_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_19_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_19_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_19_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_19_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_19_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_19_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_19_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_19_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_19_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_19_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_19_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_19_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_19_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_19_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_19_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_19_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_19_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_19_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_19_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_19_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_19_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_19_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_19_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_19_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_19_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_19_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_19_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_19_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_19_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_19_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_19_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_19_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_19_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_19_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_19_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_19_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_19_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_19_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_19_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_19_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_19_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_19_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_19_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_19_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_19_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_19_bits_st_dep_mask <= _GEN_1685;
      ldq_19_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1608) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_19_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_19_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_19_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_19_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_19_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_19_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_19_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_19_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_19_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_19_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_19_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_19_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_19_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_19_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_19_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_19_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_19_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_19_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_19_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_19_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_19_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_19_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_19_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_19_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_19_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_19_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_19_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_19_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_19_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_19_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_19_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_19_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_19_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_19_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_19_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_19_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_19_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_19_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_19_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_19_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_19_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_19_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_19_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_19_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_19_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_19_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_19_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_19_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_19_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_19_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_19_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_19_bits_st_dep_mask <= next_live_store_mask;
      ldq_19_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_19_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_19_bits_st_dep_mask;
    if (ldq_19_valid)
      ldq_19_bits_uop_br_mask <= ldq_19_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2300)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2089)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1800)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1608)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2780) begin
      if (_exe_tlb_uop_T_9)
        ldq_19_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_19_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_19_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_19_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_19_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_19_bits_addr_bits <= casez_tmp_202;
        else
          ldq_19_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_19_bits_addr_bits <= _GEN_280;
      ldq_19_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_19_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2665) begin
      if (_exe_tlb_uop_T_2)
        ldq_19_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_19_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_19_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_19_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_19_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_19_bits_addr_bits <= casez_tmp_202;
        else
          ldq_19_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_19_bits_addr_bits <= _GEN_274;
      ldq_19_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_19_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2300)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2089)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1800)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1608)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_19_bits_addr_valid <= ~_GEN_5749 & _GEN_5640 & _GEN_5577 & _GEN_5482 & (_GEN_5336 ? ~_GEN_5259 & _GEN_2781 : ~_GEN_5355 & _GEN_2781);
    ldq_19_bits_executed <= ~_GEN_5749 & _GEN_5640 & _GEN_5577 & _GEN_5482 & _GEN_5387 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1493) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1454)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_354 & _GEN_5064 : ~(_GEN_1425 & _GEN_354) & _GEN_5064) : _GEN_5064) | (dis_ld_val_3 ? ~_GEN_2225 & _GEN_1864 : ~_GEN_2089 & _GEN_1864));
    ldq_19_bits_succeeded <= _GEN_5640 & _GEN_5577 & _GEN_5482 & _GEN_5387 & (_GEN_5183 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h13 ? _ldq_bits_succeeded_T_1 : _GEN_5118 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h13 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2225 & _GEN_1896 : ~_GEN_2089 & _GEN_1896) : casez_tmp_490) : casez_tmp_524);
    ldq_19_bits_order_fail <= _GEN_5640 & _GEN_5577 & _GEN_5482 & _GEN_5387 & (_GEN_794 ? _GEN_2951 : _GEN_796 ? _GEN_797 | _GEN_2951 : _GEN_799 | _GEN_2951);
    ldq_19_bits_observed <= _GEN_794 | _GEN_781 | (dis_ld_val_3 ? ~_GEN_2225 & _GEN_1960 : ~_GEN_2089 & _GEN_1960);
    ldq_19_bits_forward_std_val <= _GEN_5640 & _GEN_5577 & _GEN_5482 & _GEN_5387 & (~_GEN_1508 & _GEN_5182 | ~_GEN_1468 & _GEN_5117 | (dis_ld_val_3 ? ~_GEN_2225 & _GEN_1992 : ~_GEN_2089 & _GEN_1992));
    if (_GEN_5183) begin
      if (_GEN_5118) begin
      end
      else
        ldq_19_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_19_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_20_valid <= ~_GEN_5749 & _GEN_5641 & _GEN_5578 & _GEN_5483 & (_GEN_5336 ? ~_GEN_5260 & _GEN_2229 : ~_GEN_5356 & _GEN_2229);
    if (_GEN_2302) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_20_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_20_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_20_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_20_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_20_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_20_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_20_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_20_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_20_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_20_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_20_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_20_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_20_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_20_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_20_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_20_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_20_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_20_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_20_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_20_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_20_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_20_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_20_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_20_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_20_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_20_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_20_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_20_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_20_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_20_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_20_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_20_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_20_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_20_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_20_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_20_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_20_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_20_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_20_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_20_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_20_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_20_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_20_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_20_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_20_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_20_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_20_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_20_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_20_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_20_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_20_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_20_bits_st_dep_mask <= _GEN_2166;
      ldq_20_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2090) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_20_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_20_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_20_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_20_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_20_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_20_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_20_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_20_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_20_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_20_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_20_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_20_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_20_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_20_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_20_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_20_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_20_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_20_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_20_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_20_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_20_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_20_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_20_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_20_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_20_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_20_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_20_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_20_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_20_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_20_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_20_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_20_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_20_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_20_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_20_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_20_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_20_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_20_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_20_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_20_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_20_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_20_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_20_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_20_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_20_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_20_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_20_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_20_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_20_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_20_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_20_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_20_bits_st_dep_mask <= _GEN_2069;
      ldq_20_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1801) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_20_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_20_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_20_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_20_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_20_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_20_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_20_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_20_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_20_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_20_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_20_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_20_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_20_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_20_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_20_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_20_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_20_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_20_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_20_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_20_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_20_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_20_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_20_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_20_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_20_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_20_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_20_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_20_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_20_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_20_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_20_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_20_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_20_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_20_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_20_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_20_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_20_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_20_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_20_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_20_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_20_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_20_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_20_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_20_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_20_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_20_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_20_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_20_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_20_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_20_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_20_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_20_bits_st_dep_mask <= _GEN_1685;
      ldq_20_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1609) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_20_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_20_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_20_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_20_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_20_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_20_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_20_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_20_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_20_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_20_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_20_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_20_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_20_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_20_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_20_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_20_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_20_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_20_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_20_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_20_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_20_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_20_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_20_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_20_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_20_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_20_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_20_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_20_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_20_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_20_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_20_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_20_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_20_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_20_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_20_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_20_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_20_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_20_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_20_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_20_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_20_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_20_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_20_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_20_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_20_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_20_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_20_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_20_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_20_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_20_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_20_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_20_bits_st_dep_mask <= next_live_store_mask;
      ldq_20_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_20_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_20_bits_st_dep_mask;
    if (ldq_20_valid)
      ldq_20_bits_uop_br_mask <= ldq_20_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2302)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2090)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1801)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1609)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2782) begin
      if (_exe_tlb_uop_T_9)
        ldq_20_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_20_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_20_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_20_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_20_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_20_bits_addr_bits <= casez_tmp_202;
        else
          ldq_20_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_20_bits_addr_bits <= _GEN_280;
      ldq_20_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_20_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2666) begin
      if (_exe_tlb_uop_T_2)
        ldq_20_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_20_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_20_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_20_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_20_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_20_bits_addr_bits <= casez_tmp_202;
        else
          ldq_20_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_20_bits_addr_bits <= _GEN_274;
      ldq_20_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_20_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2302)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2090)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1801)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1609)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_20_bits_addr_valid <= ~_GEN_5749 & _GEN_5641 & _GEN_5578 & _GEN_5483 & (_GEN_5336 ? ~_GEN_5260 & _GEN_2783 : ~_GEN_5356 & _GEN_2783);
    ldq_20_bits_executed <= ~_GEN_5749 & _GEN_5641 & _GEN_5578 & _GEN_5483 & _GEN_5388 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1494) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1455)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_355 & _GEN_5065 : ~(_GEN_1425 & _GEN_355) & _GEN_5065) : _GEN_5065) | (dis_ld_val_3 ? ~_GEN_2228 & _GEN_1865 : ~_GEN_2090 & _GEN_1865));
    ldq_20_bits_succeeded <= _GEN_5641 & _GEN_5578 & _GEN_5483 & _GEN_5388 & (_GEN_5185 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h14 ? _ldq_bits_succeeded_T_1 : _GEN_5120 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h14 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2228 & _GEN_1897 : ~_GEN_2090 & _GEN_1897) : casez_tmp_490) : casez_tmp_524);
    ldq_20_bits_order_fail <= _GEN_5641 & _GEN_5578 & _GEN_5483 & _GEN_5388 & (_GEN_817 ? _GEN_2952 : _GEN_819 ? _GEN_820 | _GEN_2952 : _GEN_822 | _GEN_2952);
    ldq_20_bits_observed <= _GEN_817 | _GEN_804 | (dis_ld_val_3 ? ~_GEN_2228 & _GEN_1961 : ~_GEN_2090 & _GEN_1961);
    ldq_20_bits_forward_std_val <= _GEN_5641 & _GEN_5578 & _GEN_5483 & _GEN_5388 & (~_GEN_1508 & _GEN_5184 | ~_GEN_1468 & _GEN_5119 | (dis_ld_val_3 ? ~_GEN_2228 & _GEN_1993 : ~_GEN_2090 & _GEN_1993));
    if (_GEN_5185) begin
      if (_GEN_5120) begin
      end
      else
        ldq_20_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_20_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_21_valid <= ~_GEN_5749 & _GEN_5642 & _GEN_5579 & _GEN_5484 & (_GEN_5336 ? ~_GEN_5261 & _GEN_2232 : ~_GEN_5357 & _GEN_2232);
    if (_GEN_2304) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_21_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_21_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_21_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_21_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_21_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_21_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_21_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_21_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_21_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_21_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_21_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_21_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_21_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_21_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_21_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_21_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_21_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_21_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_21_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_21_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_21_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_21_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_21_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_21_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_21_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_21_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_21_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_21_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_21_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_21_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_21_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_21_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_21_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_21_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_21_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_21_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_21_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_21_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_21_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_21_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_21_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_21_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_21_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_21_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_21_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_21_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_21_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_21_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_21_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_21_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_21_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_21_bits_st_dep_mask <= _GEN_2166;
      ldq_21_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2091) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_21_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_21_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_21_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_21_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_21_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_21_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_21_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_21_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_21_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_21_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_21_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_21_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_21_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_21_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_21_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_21_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_21_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_21_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_21_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_21_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_21_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_21_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_21_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_21_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_21_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_21_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_21_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_21_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_21_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_21_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_21_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_21_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_21_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_21_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_21_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_21_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_21_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_21_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_21_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_21_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_21_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_21_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_21_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_21_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_21_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_21_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_21_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_21_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_21_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_21_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_21_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_21_bits_st_dep_mask <= _GEN_2069;
      ldq_21_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1802) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_21_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_21_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_21_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_21_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_21_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_21_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_21_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_21_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_21_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_21_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_21_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_21_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_21_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_21_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_21_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_21_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_21_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_21_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_21_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_21_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_21_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_21_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_21_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_21_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_21_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_21_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_21_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_21_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_21_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_21_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_21_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_21_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_21_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_21_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_21_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_21_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_21_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_21_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_21_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_21_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_21_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_21_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_21_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_21_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_21_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_21_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_21_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_21_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_21_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_21_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_21_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_21_bits_st_dep_mask <= _GEN_1685;
      ldq_21_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1610) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_21_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_21_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_21_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_21_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_21_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_21_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_21_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_21_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_21_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_21_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_21_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_21_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_21_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_21_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_21_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_21_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_21_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_21_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_21_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_21_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_21_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_21_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_21_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_21_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_21_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_21_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_21_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_21_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_21_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_21_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_21_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_21_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_21_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_21_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_21_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_21_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_21_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_21_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_21_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_21_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_21_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_21_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_21_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_21_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_21_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_21_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_21_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_21_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_21_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_21_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_21_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_21_bits_st_dep_mask <= next_live_store_mask;
      ldq_21_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_21_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_21_bits_st_dep_mask;
    if (ldq_21_valid)
      ldq_21_bits_uop_br_mask <= ldq_21_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2304)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2091)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1802)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1610)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2784) begin
      if (_exe_tlb_uop_T_9)
        ldq_21_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_21_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_21_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_21_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_21_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_21_bits_addr_bits <= casez_tmp_202;
        else
          ldq_21_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_21_bits_addr_bits <= _GEN_280;
      ldq_21_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_21_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2667) begin
      if (_exe_tlb_uop_T_2)
        ldq_21_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_21_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_21_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_21_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_21_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_21_bits_addr_bits <= casez_tmp_202;
        else
          ldq_21_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_21_bits_addr_bits <= _GEN_274;
      ldq_21_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_21_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2304)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2091)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1802)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1610)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_21_bits_addr_valid <= ~_GEN_5749 & _GEN_5642 & _GEN_5579 & _GEN_5484 & (_GEN_5336 ? ~_GEN_5261 & _GEN_2785 : ~_GEN_5357 & _GEN_2785);
    ldq_21_bits_executed <= ~_GEN_5749 & _GEN_5642 & _GEN_5579 & _GEN_5484 & _GEN_5389 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1495) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1456)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_356 & _GEN_5066 : ~(_GEN_1425 & _GEN_356) & _GEN_5066) : _GEN_5066) | (dis_ld_val_3 ? ~_GEN_2231 & _GEN_1866 : ~_GEN_2091 & _GEN_1866));
    ldq_21_bits_succeeded <= _GEN_5642 & _GEN_5579 & _GEN_5484 & _GEN_5389 & (_GEN_5187 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h15 ? _ldq_bits_succeeded_T_1 : _GEN_5122 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h15 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2231 & _GEN_1898 : ~_GEN_2091 & _GEN_1898) : casez_tmp_490) : casez_tmp_524);
    ldq_21_bits_order_fail <= _GEN_5642 & _GEN_5579 & _GEN_5484 & _GEN_5389 & (_GEN_840 ? _GEN_2953 : _GEN_842 ? _GEN_843 | _GEN_2953 : _GEN_845 | _GEN_2953);
    ldq_21_bits_observed <= _GEN_840 | _GEN_827 | (dis_ld_val_3 ? ~_GEN_2231 & _GEN_1962 : ~_GEN_2091 & _GEN_1962);
    ldq_21_bits_forward_std_val <= _GEN_5642 & _GEN_5579 & _GEN_5484 & _GEN_5389 & (~_GEN_1508 & _GEN_5186 | ~_GEN_1468 & _GEN_5121 | (dis_ld_val_3 ? ~_GEN_2231 & _GEN_1994 : ~_GEN_2091 & _GEN_1994));
    if (_GEN_5187) begin
      if (_GEN_5122) begin
      end
      else
        ldq_21_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_21_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_22_valid <= ~_GEN_5749 & _GEN_5643 & _GEN_5580 & _GEN_5485 & (_GEN_5336 ? ~_GEN_5262 & _GEN_2235 : ~_GEN_5358 & _GEN_2235);
    if (_GEN_2306) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_22_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_22_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_22_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_22_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_22_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_22_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_22_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_22_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_22_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_22_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_22_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_22_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_22_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_22_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_22_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_22_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_22_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_22_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_22_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_22_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_22_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_22_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_22_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_22_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_22_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_22_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_22_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_22_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_22_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_22_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_22_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_22_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_22_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_22_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_22_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_22_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_22_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_22_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_22_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_22_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_22_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_22_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_22_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_22_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_22_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_22_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_22_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_22_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_22_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_22_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_22_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_22_bits_st_dep_mask <= _GEN_2166;
      ldq_22_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2092) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_22_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_22_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_22_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_22_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_22_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_22_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_22_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_22_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_22_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_22_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_22_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_22_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_22_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_22_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_22_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_22_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_22_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_22_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_22_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_22_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_22_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_22_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_22_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_22_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_22_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_22_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_22_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_22_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_22_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_22_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_22_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_22_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_22_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_22_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_22_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_22_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_22_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_22_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_22_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_22_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_22_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_22_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_22_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_22_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_22_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_22_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_22_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_22_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_22_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_22_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_22_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_22_bits_st_dep_mask <= _GEN_2069;
      ldq_22_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1803) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_22_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_22_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_22_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_22_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_22_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_22_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_22_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_22_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_22_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_22_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_22_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_22_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_22_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_22_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_22_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_22_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_22_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_22_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_22_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_22_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_22_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_22_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_22_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_22_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_22_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_22_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_22_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_22_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_22_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_22_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_22_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_22_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_22_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_22_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_22_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_22_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_22_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_22_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_22_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_22_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_22_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_22_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_22_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_22_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_22_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_22_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_22_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_22_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_22_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_22_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_22_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_22_bits_st_dep_mask <= _GEN_1685;
      ldq_22_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1611) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_22_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_22_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_22_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_22_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_22_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_22_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_22_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_22_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_22_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_22_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_22_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_22_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_22_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_22_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_22_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_22_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_22_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_22_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_22_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_22_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_22_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_22_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_22_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_22_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_22_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_22_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_22_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_22_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_22_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_22_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_22_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_22_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_22_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_22_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_22_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_22_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_22_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_22_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_22_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_22_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_22_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_22_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_22_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_22_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_22_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_22_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_22_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_22_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_22_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_22_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_22_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_22_bits_st_dep_mask <= next_live_store_mask;
      ldq_22_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_22_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_22_bits_st_dep_mask;
    if (ldq_22_valid)
      ldq_22_bits_uop_br_mask <= ldq_22_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2306)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2092)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1803)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1611)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2786) begin
      if (_exe_tlb_uop_T_9)
        ldq_22_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_22_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_22_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_22_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_22_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_22_bits_addr_bits <= casez_tmp_202;
        else
          ldq_22_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_22_bits_addr_bits <= _GEN_280;
      ldq_22_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_22_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2668) begin
      if (_exe_tlb_uop_T_2)
        ldq_22_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_22_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_22_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_22_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_22_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_22_bits_addr_bits <= casez_tmp_202;
        else
          ldq_22_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_22_bits_addr_bits <= _GEN_274;
      ldq_22_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_22_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2306)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2092)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1803)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1611)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_22_bits_addr_valid <= ~_GEN_5749 & _GEN_5643 & _GEN_5580 & _GEN_5485 & (_GEN_5336 ? ~_GEN_5262 & _GEN_2787 : ~_GEN_5358 & _GEN_2787);
    ldq_22_bits_executed <= ~_GEN_5749 & _GEN_5643 & _GEN_5580 & _GEN_5485 & _GEN_5390 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1496) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1457)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_357 & _GEN_5067 : ~(_GEN_1425 & _GEN_357) & _GEN_5067) : _GEN_5067) | (dis_ld_val_3 ? ~_GEN_2234 & _GEN_1867 : ~_GEN_2092 & _GEN_1867));
    ldq_22_bits_succeeded <= _GEN_5643 & _GEN_5580 & _GEN_5485 & _GEN_5390 & (_GEN_5189 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h16 ? _ldq_bits_succeeded_T_1 : _GEN_5124 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h16 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2234 & _GEN_1899 : ~_GEN_2092 & _GEN_1899) : casez_tmp_490) : casez_tmp_524);
    ldq_22_bits_order_fail <= _GEN_5643 & _GEN_5580 & _GEN_5485 & _GEN_5390 & (_GEN_863 ? _GEN_2954 : _GEN_865 ? _GEN_866 | _GEN_2954 : _GEN_868 | _GEN_2954);
    ldq_22_bits_observed <= _GEN_863 | _GEN_850 | (dis_ld_val_3 ? ~_GEN_2234 & _GEN_1963 : ~_GEN_2092 & _GEN_1963);
    ldq_22_bits_forward_std_val <= _GEN_5643 & _GEN_5580 & _GEN_5485 & _GEN_5390 & (~_GEN_1508 & _GEN_5188 | ~_GEN_1468 & _GEN_5123 | (dis_ld_val_3 ? ~_GEN_2234 & _GEN_1995 : ~_GEN_2092 & _GEN_1995));
    if (_GEN_5189) begin
      if (_GEN_5124) begin
      end
      else
        ldq_22_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_22_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_23_valid <= ~_GEN_5749 & _GEN_5644 & _GEN_5581 & _GEN_5486 & (_GEN_5336 ? ~_GEN_5263 & _GEN_2238 : ~_GEN_5359 & _GEN_2238);
    if (_GEN_2308) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_23_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_23_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_23_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_23_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_23_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_23_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_23_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_23_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_23_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_23_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_23_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_23_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_23_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_23_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_23_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_23_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_23_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_23_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_23_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_23_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_23_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_23_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_23_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_23_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_23_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_23_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_23_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_23_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_23_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_23_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_23_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_23_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_23_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_23_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_23_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_23_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_23_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_23_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_23_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_23_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_23_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_23_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_23_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_23_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_23_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_23_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_23_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_23_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_23_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_23_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_23_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_23_bits_st_dep_mask <= _GEN_2166;
      ldq_23_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2093) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_23_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_23_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_23_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_23_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_23_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_23_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_23_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_23_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_23_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_23_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_23_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_23_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_23_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_23_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_23_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_23_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_23_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_23_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_23_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_23_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_23_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_23_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_23_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_23_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_23_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_23_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_23_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_23_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_23_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_23_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_23_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_23_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_23_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_23_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_23_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_23_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_23_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_23_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_23_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_23_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_23_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_23_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_23_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_23_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_23_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_23_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_23_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_23_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_23_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_23_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_23_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_23_bits_st_dep_mask <= _GEN_2069;
      ldq_23_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1804) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_23_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_23_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_23_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_23_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_23_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_23_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_23_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_23_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_23_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_23_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_23_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_23_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_23_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_23_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_23_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_23_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_23_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_23_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_23_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_23_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_23_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_23_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_23_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_23_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_23_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_23_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_23_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_23_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_23_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_23_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_23_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_23_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_23_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_23_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_23_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_23_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_23_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_23_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_23_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_23_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_23_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_23_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_23_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_23_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_23_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_23_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_23_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_23_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_23_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_23_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_23_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_23_bits_st_dep_mask <= _GEN_1685;
      ldq_23_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1612) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_23_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_23_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_23_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_23_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_23_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_23_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_23_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_23_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_23_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_23_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_23_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_23_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_23_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_23_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_23_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_23_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_23_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_23_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_23_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_23_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_23_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_23_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_23_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_23_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_23_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_23_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_23_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_23_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_23_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_23_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_23_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_23_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_23_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_23_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_23_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_23_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_23_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_23_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_23_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_23_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_23_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_23_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_23_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_23_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_23_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_23_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_23_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_23_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_23_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_23_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_23_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_23_bits_st_dep_mask <= next_live_store_mask;
      ldq_23_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_23_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_23_bits_st_dep_mask;
    if (ldq_23_valid)
      ldq_23_bits_uop_br_mask <= ldq_23_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2308)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2093)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1804)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1612)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2788) begin
      if (_exe_tlb_uop_T_9)
        ldq_23_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_23_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_23_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_23_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_23_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_23_bits_addr_bits <= casez_tmp_202;
        else
          ldq_23_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_23_bits_addr_bits <= _GEN_280;
      ldq_23_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_23_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2669) begin
      if (_exe_tlb_uop_T_2)
        ldq_23_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_23_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_23_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_23_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_23_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_23_bits_addr_bits <= casez_tmp_202;
        else
          ldq_23_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_23_bits_addr_bits <= _GEN_274;
      ldq_23_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_23_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2308)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2093)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1804)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1612)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_23_bits_addr_valid <= ~_GEN_5749 & _GEN_5644 & _GEN_5581 & _GEN_5486 & (_GEN_5336 ? ~_GEN_5263 & _GEN_2789 : ~_GEN_5359 & _GEN_2789);
    ldq_23_bits_executed <= ~_GEN_5749 & _GEN_5644 & _GEN_5581 & _GEN_5486 & _GEN_5391 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1497) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1458)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_358 & _GEN_5068 : ~(_GEN_1425 & _GEN_358) & _GEN_5068) : _GEN_5068) | (dis_ld_val_3 ? ~_GEN_2237 & _GEN_1868 : ~_GEN_2093 & _GEN_1868));
    ldq_23_bits_succeeded <= _GEN_5644 & _GEN_5581 & _GEN_5486 & _GEN_5391 & (_GEN_5191 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h17 ? _ldq_bits_succeeded_T_1 : _GEN_5126 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h17 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2237 & _GEN_1900 : ~_GEN_2093 & _GEN_1900) : casez_tmp_490) : casez_tmp_524);
    ldq_23_bits_order_fail <= _GEN_5644 & _GEN_5581 & _GEN_5486 & _GEN_5391 & (_GEN_886 ? _GEN_2955 : _GEN_888 ? _GEN_889 | _GEN_2955 : _GEN_891 | _GEN_2955);
    ldq_23_bits_observed <= _GEN_886 | _GEN_873 | (dis_ld_val_3 ? ~_GEN_2237 & _GEN_1964 : ~_GEN_2093 & _GEN_1964);
    ldq_23_bits_forward_std_val <= _GEN_5644 & _GEN_5581 & _GEN_5486 & _GEN_5391 & (~_GEN_1508 & _GEN_5190 | ~_GEN_1468 & _GEN_5125 | (dis_ld_val_3 ? ~_GEN_2237 & _GEN_1996 : ~_GEN_2093 & _GEN_1996));
    if (_GEN_5191) begin
      if (_GEN_5126) begin
      end
      else
        ldq_23_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_23_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_24_valid <= ~_GEN_5749 & _GEN_5645 & _GEN_5582 & _GEN_5487 & (_GEN_5336 ? ~_GEN_5264 & _GEN_2241 : ~_GEN_5360 & _GEN_2241);
    if (_GEN_2310) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_24_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_24_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_24_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_24_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_24_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_24_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_24_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_24_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_24_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_24_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_24_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_24_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_24_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_24_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_24_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_24_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_24_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_24_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_24_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_24_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_24_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_24_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_24_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_24_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_24_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_24_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_24_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_24_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_24_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_24_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_24_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_24_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_24_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_24_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_24_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_24_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_24_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_24_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_24_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_24_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_24_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_24_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_24_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_24_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_24_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_24_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_24_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_24_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_24_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_24_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_24_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_24_bits_st_dep_mask <= _GEN_2166;
      ldq_24_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2094) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_24_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_24_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_24_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_24_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_24_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_24_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_24_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_24_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_24_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_24_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_24_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_24_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_24_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_24_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_24_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_24_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_24_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_24_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_24_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_24_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_24_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_24_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_24_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_24_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_24_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_24_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_24_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_24_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_24_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_24_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_24_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_24_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_24_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_24_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_24_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_24_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_24_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_24_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_24_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_24_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_24_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_24_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_24_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_24_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_24_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_24_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_24_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_24_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_24_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_24_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_24_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_24_bits_st_dep_mask <= _GEN_2069;
      ldq_24_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1805) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_24_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_24_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_24_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_24_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_24_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_24_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_24_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_24_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_24_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_24_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_24_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_24_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_24_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_24_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_24_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_24_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_24_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_24_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_24_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_24_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_24_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_24_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_24_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_24_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_24_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_24_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_24_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_24_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_24_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_24_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_24_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_24_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_24_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_24_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_24_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_24_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_24_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_24_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_24_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_24_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_24_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_24_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_24_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_24_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_24_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_24_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_24_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_24_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_24_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_24_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_24_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_24_bits_st_dep_mask <= _GEN_1685;
      ldq_24_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1613) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_24_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_24_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_24_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_24_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_24_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_24_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_24_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_24_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_24_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_24_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_24_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_24_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_24_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_24_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_24_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_24_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_24_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_24_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_24_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_24_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_24_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_24_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_24_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_24_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_24_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_24_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_24_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_24_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_24_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_24_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_24_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_24_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_24_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_24_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_24_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_24_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_24_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_24_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_24_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_24_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_24_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_24_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_24_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_24_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_24_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_24_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_24_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_24_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_24_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_24_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_24_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_24_bits_st_dep_mask <= next_live_store_mask;
      ldq_24_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_24_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_24_bits_st_dep_mask;
    if (ldq_24_valid)
      ldq_24_bits_uop_br_mask <= ldq_24_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2310)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2094)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1805)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1613)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2790) begin
      if (_exe_tlb_uop_T_9)
        ldq_24_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_24_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_24_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_24_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_24_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_24_bits_addr_bits <= casez_tmp_202;
        else
          ldq_24_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_24_bits_addr_bits <= _GEN_280;
      ldq_24_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_24_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2670) begin
      if (_exe_tlb_uop_T_2)
        ldq_24_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_24_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_24_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_24_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_24_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_24_bits_addr_bits <= casez_tmp_202;
        else
          ldq_24_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_24_bits_addr_bits <= _GEN_274;
      ldq_24_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_24_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2310)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2094)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1805)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1613)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_24_bits_addr_valid <= ~_GEN_5749 & _GEN_5645 & _GEN_5582 & _GEN_5487 & (_GEN_5336 ? ~_GEN_5264 & _GEN_2791 : ~_GEN_5360 & _GEN_2791);
    ldq_24_bits_executed <= ~_GEN_5749 & _GEN_5645 & _GEN_5582 & _GEN_5487 & _GEN_5392 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1498) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1459)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_359 & _GEN_5069 : ~(_GEN_1425 & _GEN_359) & _GEN_5069) : _GEN_5069) | (dis_ld_val_3 ? ~_GEN_2240 & _GEN_1869 : ~_GEN_2094 & _GEN_1869));
    ldq_24_bits_succeeded <= _GEN_5645 & _GEN_5582 & _GEN_5487 & _GEN_5392 & (_GEN_5193 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h18 ? _ldq_bits_succeeded_T_1 : _GEN_5128 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h18 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2240 & _GEN_1901 : ~_GEN_2094 & _GEN_1901) : casez_tmp_490) : casez_tmp_524);
    ldq_24_bits_order_fail <= _GEN_5645 & _GEN_5582 & _GEN_5487 & _GEN_5392 & (_GEN_909 ? _GEN_2956 : _GEN_911 ? _GEN_912 | _GEN_2956 : _GEN_914 | _GEN_2956);
    ldq_24_bits_observed <= _GEN_909 | _GEN_896 | (dis_ld_val_3 ? ~_GEN_2240 & _GEN_1965 : ~_GEN_2094 & _GEN_1965);
    ldq_24_bits_forward_std_val <= _GEN_5645 & _GEN_5582 & _GEN_5487 & _GEN_5392 & (~_GEN_1508 & _GEN_5192 | ~_GEN_1468 & _GEN_5127 | (dis_ld_val_3 ? ~_GEN_2240 & _GEN_1997 : ~_GEN_2094 & _GEN_1997));
    if (_GEN_5193) begin
      if (_GEN_5128) begin
      end
      else
        ldq_24_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_24_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_25_valid <= ~_GEN_5749 & _GEN_5646 & _GEN_5583 & _GEN_5488 & (_GEN_5336 ? ~_GEN_5265 & _GEN_2244 : ~_GEN_5361 & _GEN_2244);
    if (_GEN_2312) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_25_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_25_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_25_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_25_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_25_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_25_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_25_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_25_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_25_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_25_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_25_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_25_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_25_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_25_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_25_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_25_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_25_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_25_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_25_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_25_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_25_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_25_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_25_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_25_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_25_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_25_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_25_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_25_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_25_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_25_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_25_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_25_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_25_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_25_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_25_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_25_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_25_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_25_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_25_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_25_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_25_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_25_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_25_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_25_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_25_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_25_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_25_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_25_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_25_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_25_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_25_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_25_bits_st_dep_mask <= _GEN_2166;
      ldq_25_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2095) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_25_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_25_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_25_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_25_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_25_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_25_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_25_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_25_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_25_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_25_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_25_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_25_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_25_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_25_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_25_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_25_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_25_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_25_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_25_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_25_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_25_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_25_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_25_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_25_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_25_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_25_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_25_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_25_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_25_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_25_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_25_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_25_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_25_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_25_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_25_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_25_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_25_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_25_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_25_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_25_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_25_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_25_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_25_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_25_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_25_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_25_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_25_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_25_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_25_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_25_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_25_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_25_bits_st_dep_mask <= _GEN_2069;
      ldq_25_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1806) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_25_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_25_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_25_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_25_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_25_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_25_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_25_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_25_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_25_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_25_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_25_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_25_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_25_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_25_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_25_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_25_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_25_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_25_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_25_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_25_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_25_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_25_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_25_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_25_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_25_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_25_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_25_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_25_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_25_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_25_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_25_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_25_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_25_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_25_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_25_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_25_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_25_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_25_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_25_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_25_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_25_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_25_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_25_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_25_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_25_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_25_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_25_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_25_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_25_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_25_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_25_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_25_bits_st_dep_mask <= _GEN_1685;
      ldq_25_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1614) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_25_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_25_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_25_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_25_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_25_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_25_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_25_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_25_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_25_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_25_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_25_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_25_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_25_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_25_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_25_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_25_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_25_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_25_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_25_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_25_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_25_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_25_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_25_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_25_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_25_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_25_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_25_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_25_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_25_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_25_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_25_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_25_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_25_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_25_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_25_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_25_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_25_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_25_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_25_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_25_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_25_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_25_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_25_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_25_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_25_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_25_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_25_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_25_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_25_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_25_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_25_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_25_bits_st_dep_mask <= next_live_store_mask;
      ldq_25_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_25_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_25_bits_st_dep_mask;
    if (ldq_25_valid)
      ldq_25_bits_uop_br_mask <= ldq_25_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2312)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2095)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1806)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1614)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2792) begin
      if (_exe_tlb_uop_T_9)
        ldq_25_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_25_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_25_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_25_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_25_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_25_bits_addr_bits <= casez_tmp_202;
        else
          ldq_25_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_25_bits_addr_bits <= _GEN_280;
      ldq_25_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_25_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2671) begin
      if (_exe_tlb_uop_T_2)
        ldq_25_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_25_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_25_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_25_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_25_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_25_bits_addr_bits <= casez_tmp_202;
        else
          ldq_25_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_25_bits_addr_bits <= _GEN_274;
      ldq_25_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_25_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2312)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2095)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1806)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1614)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_25_bits_addr_valid <= ~_GEN_5749 & _GEN_5646 & _GEN_5583 & _GEN_5488 & (_GEN_5336 ? ~_GEN_5265 & _GEN_2793 : ~_GEN_5361 & _GEN_2793);
    ldq_25_bits_executed <= ~_GEN_5749 & _GEN_5646 & _GEN_5583 & _GEN_5488 & _GEN_5393 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1499) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1460)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_360 & _GEN_5070 : ~(_GEN_1425 & _GEN_360) & _GEN_5070) : _GEN_5070) | (dis_ld_val_3 ? ~_GEN_2243 & _GEN_1870 : ~_GEN_2095 & _GEN_1870));
    ldq_25_bits_succeeded <= _GEN_5646 & _GEN_5583 & _GEN_5488 & _GEN_5393 & (_GEN_5195 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h19 ? _ldq_bits_succeeded_T_1 : _GEN_5130 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h19 ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2243 & _GEN_1902 : ~_GEN_2095 & _GEN_1902) : casez_tmp_490) : casez_tmp_524);
    ldq_25_bits_order_fail <= _GEN_5646 & _GEN_5583 & _GEN_5488 & _GEN_5393 & (_GEN_932 ? _GEN_2957 : _GEN_934 ? _GEN_935 | _GEN_2957 : _GEN_937 | _GEN_2957);
    ldq_25_bits_observed <= _GEN_932 | _GEN_919 | (dis_ld_val_3 ? ~_GEN_2243 & _GEN_1966 : ~_GEN_2095 & _GEN_1966);
    ldq_25_bits_forward_std_val <= _GEN_5646 & _GEN_5583 & _GEN_5488 & _GEN_5393 & (~_GEN_1508 & _GEN_5194 | ~_GEN_1468 & _GEN_5129 | (dis_ld_val_3 ? ~_GEN_2243 & _GEN_1998 : ~_GEN_2095 & _GEN_1998));
    if (_GEN_5195) begin
      if (_GEN_5130) begin
      end
      else
        ldq_25_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_25_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_26_valid <= ~_GEN_5749 & _GEN_5647 & _GEN_5584 & _GEN_5489 & (_GEN_5336 ? ~_GEN_5266 & _GEN_2247 : ~_GEN_5362 & _GEN_2247);
    if (_GEN_2314) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_26_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_26_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_26_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_26_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_26_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_26_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_26_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_26_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_26_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_26_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_26_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_26_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_26_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_26_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_26_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_26_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_26_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_26_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_26_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_26_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_26_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_26_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_26_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_26_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_26_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_26_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_26_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_26_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_26_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_26_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_26_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_26_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_26_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_26_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_26_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_26_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_26_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_26_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_26_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_26_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_26_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_26_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_26_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_26_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_26_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_26_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_26_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_26_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_26_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_26_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_26_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_26_bits_st_dep_mask <= _GEN_2166;
      ldq_26_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2096) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_26_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_26_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_26_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_26_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_26_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_26_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_26_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_26_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_26_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_26_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_26_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_26_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_26_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_26_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_26_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_26_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_26_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_26_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_26_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_26_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_26_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_26_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_26_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_26_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_26_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_26_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_26_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_26_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_26_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_26_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_26_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_26_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_26_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_26_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_26_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_26_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_26_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_26_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_26_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_26_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_26_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_26_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_26_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_26_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_26_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_26_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_26_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_26_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_26_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_26_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_26_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_26_bits_st_dep_mask <= _GEN_2069;
      ldq_26_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1807) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_26_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_26_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_26_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_26_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_26_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_26_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_26_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_26_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_26_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_26_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_26_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_26_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_26_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_26_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_26_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_26_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_26_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_26_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_26_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_26_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_26_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_26_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_26_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_26_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_26_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_26_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_26_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_26_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_26_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_26_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_26_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_26_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_26_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_26_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_26_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_26_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_26_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_26_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_26_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_26_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_26_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_26_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_26_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_26_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_26_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_26_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_26_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_26_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_26_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_26_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_26_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_26_bits_st_dep_mask <= _GEN_1685;
      ldq_26_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1615) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_26_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_26_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_26_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_26_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_26_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_26_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_26_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_26_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_26_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_26_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_26_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_26_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_26_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_26_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_26_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_26_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_26_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_26_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_26_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_26_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_26_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_26_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_26_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_26_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_26_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_26_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_26_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_26_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_26_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_26_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_26_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_26_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_26_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_26_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_26_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_26_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_26_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_26_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_26_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_26_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_26_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_26_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_26_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_26_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_26_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_26_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_26_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_26_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_26_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_26_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_26_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_26_bits_st_dep_mask <= next_live_store_mask;
      ldq_26_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_26_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_26_bits_st_dep_mask;
    if (ldq_26_valid)
      ldq_26_bits_uop_br_mask <= ldq_26_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2314)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2096)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1807)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1615)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2794) begin
      if (_exe_tlb_uop_T_9)
        ldq_26_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_26_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_26_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_26_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_26_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_26_bits_addr_bits <= casez_tmp_202;
        else
          ldq_26_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_26_bits_addr_bits <= _GEN_280;
      ldq_26_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_26_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2672) begin
      if (_exe_tlb_uop_T_2)
        ldq_26_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_26_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_26_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_26_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_26_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_26_bits_addr_bits <= casez_tmp_202;
        else
          ldq_26_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_26_bits_addr_bits <= _GEN_274;
      ldq_26_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_26_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2314)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2096)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1807)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1615)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_26_bits_addr_valid <= ~_GEN_5749 & _GEN_5647 & _GEN_5584 & _GEN_5489 & (_GEN_5336 ? ~_GEN_5266 & _GEN_2795 : ~_GEN_5362 & _GEN_2795);
    ldq_26_bits_executed <= ~_GEN_5749 & _GEN_5647 & _GEN_5584 & _GEN_5489 & _GEN_5394 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1500) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1461)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_361 & _GEN_5071 : ~(_GEN_1425 & _GEN_361) & _GEN_5071) : _GEN_5071) | (dis_ld_val_3 ? ~_GEN_2246 & _GEN_1871 : ~_GEN_2096 & _GEN_1871));
    ldq_26_bits_succeeded <= _GEN_5647 & _GEN_5584 & _GEN_5489 & _GEN_5394 & (_GEN_5197 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1A ? _ldq_bits_succeeded_T_1 : _GEN_5132 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1A ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2246 & _GEN_1903 : ~_GEN_2096 & _GEN_1903) : casez_tmp_490) : casez_tmp_524);
    ldq_26_bits_order_fail <= _GEN_5647 & _GEN_5584 & _GEN_5489 & _GEN_5394 & (_GEN_955 ? _GEN_2958 : _GEN_957 ? _GEN_958 | _GEN_2958 : _GEN_960 | _GEN_2958);
    ldq_26_bits_observed <= _GEN_955 | _GEN_942 | (dis_ld_val_3 ? ~_GEN_2246 & _GEN_1967 : ~_GEN_2096 & _GEN_1967);
    ldq_26_bits_forward_std_val <= _GEN_5647 & _GEN_5584 & _GEN_5489 & _GEN_5394 & (~_GEN_1508 & _GEN_5196 | ~_GEN_1468 & _GEN_5131 | (dis_ld_val_3 ? ~_GEN_2246 & _GEN_1999 : ~_GEN_2096 & _GEN_1999));
    if (_GEN_5197) begin
      if (_GEN_5132) begin
      end
      else
        ldq_26_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_26_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_27_valid <= ~_GEN_5749 & _GEN_5648 & _GEN_5585 & _GEN_5490 & (_GEN_5336 ? ~_GEN_5267 & _GEN_2250 : ~_GEN_5363 & _GEN_2250);
    if (_GEN_2316) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_27_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_27_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_27_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_27_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_27_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_27_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_27_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_27_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_27_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_27_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_27_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_27_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_27_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_27_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_27_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_27_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_27_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_27_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_27_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_27_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_27_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_27_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_27_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_27_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_27_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_27_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_27_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_27_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_27_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_27_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_27_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_27_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_27_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_27_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_27_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_27_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_27_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_27_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_27_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_27_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_27_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_27_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_27_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_27_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_27_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_27_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_27_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_27_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_27_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_27_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_27_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_27_bits_st_dep_mask <= _GEN_2166;
      ldq_27_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2097) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_27_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_27_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_27_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_27_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_27_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_27_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_27_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_27_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_27_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_27_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_27_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_27_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_27_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_27_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_27_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_27_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_27_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_27_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_27_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_27_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_27_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_27_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_27_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_27_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_27_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_27_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_27_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_27_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_27_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_27_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_27_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_27_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_27_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_27_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_27_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_27_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_27_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_27_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_27_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_27_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_27_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_27_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_27_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_27_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_27_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_27_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_27_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_27_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_27_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_27_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_27_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_27_bits_st_dep_mask <= _GEN_2069;
      ldq_27_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1808) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_27_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_27_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_27_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_27_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_27_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_27_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_27_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_27_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_27_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_27_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_27_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_27_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_27_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_27_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_27_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_27_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_27_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_27_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_27_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_27_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_27_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_27_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_27_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_27_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_27_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_27_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_27_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_27_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_27_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_27_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_27_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_27_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_27_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_27_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_27_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_27_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_27_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_27_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_27_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_27_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_27_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_27_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_27_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_27_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_27_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_27_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_27_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_27_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_27_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_27_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_27_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_27_bits_st_dep_mask <= _GEN_1685;
      ldq_27_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1616) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_27_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_27_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_27_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_27_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_27_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_27_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_27_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_27_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_27_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_27_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_27_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_27_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_27_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_27_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_27_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_27_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_27_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_27_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_27_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_27_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_27_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_27_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_27_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_27_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_27_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_27_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_27_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_27_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_27_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_27_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_27_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_27_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_27_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_27_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_27_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_27_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_27_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_27_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_27_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_27_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_27_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_27_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_27_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_27_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_27_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_27_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_27_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_27_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_27_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_27_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_27_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_27_bits_st_dep_mask <= next_live_store_mask;
      ldq_27_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_27_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_27_bits_st_dep_mask;
    if (ldq_27_valid)
      ldq_27_bits_uop_br_mask <= ldq_27_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2316)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2097)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1808)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1616)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2796) begin
      if (_exe_tlb_uop_T_9)
        ldq_27_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_27_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_27_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_27_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_27_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_27_bits_addr_bits <= casez_tmp_202;
        else
          ldq_27_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_27_bits_addr_bits <= _GEN_280;
      ldq_27_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_27_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2673) begin
      if (_exe_tlb_uop_T_2)
        ldq_27_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_27_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_27_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_27_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_27_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_27_bits_addr_bits <= casez_tmp_202;
        else
          ldq_27_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_27_bits_addr_bits <= _GEN_274;
      ldq_27_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_27_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2316)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2097)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1808)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1616)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_27_bits_addr_valid <= ~_GEN_5749 & _GEN_5648 & _GEN_5585 & _GEN_5490 & (_GEN_5336 ? ~_GEN_5267 & _GEN_2797 : ~_GEN_5363 & _GEN_2797);
    ldq_27_bits_executed <= ~_GEN_5749 & _GEN_5648 & _GEN_5585 & _GEN_5490 & _GEN_5395 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1501) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1462)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_362 & _GEN_5072 : ~(_GEN_1425 & _GEN_362) & _GEN_5072) : _GEN_5072) | (dis_ld_val_3 ? ~_GEN_2249 & _GEN_1872 : ~_GEN_2097 & _GEN_1872));
    ldq_27_bits_succeeded <= _GEN_5648 & _GEN_5585 & _GEN_5490 & _GEN_5395 & (_GEN_5199 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1B ? _ldq_bits_succeeded_T_1 : _GEN_5134 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1B ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2249 & _GEN_1904 : ~_GEN_2097 & _GEN_1904) : casez_tmp_490) : casez_tmp_524);
    ldq_27_bits_order_fail <= _GEN_5648 & _GEN_5585 & _GEN_5490 & _GEN_5395 & (_GEN_978 ? _GEN_2959 : _GEN_980 ? _GEN_981 | _GEN_2959 : _GEN_983 | _GEN_2959);
    ldq_27_bits_observed <= _GEN_978 | _GEN_965 | (dis_ld_val_3 ? ~_GEN_2249 & _GEN_1968 : ~_GEN_2097 & _GEN_1968);
    ldq_27_bits_forward_std_val <= _GEN_5648 & _GEN_5585 & _GEN_5490 & _GEN_5395 & (~_GEN_1508 & _GEN_5198 | ~_GEN_1468 & _GEN_5133 | (dis_ld_val_3 ? ~_GEN_2249 & _GEN_2000 : ~_GEN_2097 & _GEN_2000));
    if (_GEN_5199) begin
      if (_GEN_5134) begin
      end
      else
        ldq_27_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_27_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_28_valid <= ~_GEN_5749 & _GEN_5649 & _GEN_5586 & _GEN_5491 & (_GEN_5336 ? ~_GEN_5268 & _GEN_2253 : ~_GEN_5364 & _GEN_2253);
    if (_GEN_2318) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_28_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_28_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_28_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_28_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_28_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_28_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_28_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_28_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_28_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_28_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_28_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_28_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_28_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_28_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_28_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_28_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_28_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_28_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_28_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_28_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_28_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_28_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_28_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_28_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_28_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_28_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_28_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_28_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_28_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_28_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_28_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_28_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_28_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_28_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_28_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_28_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_28_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_28_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_28_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_28_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_28_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_28_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_28_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_28_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_28_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_28_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_28_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_28_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_28_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_28_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_28_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_28_bits_st_dep_mask <= _GEN_2166;
      ldq_28_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2098) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_28_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_28_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_28_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_28_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_28_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_28_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_28_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_28_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_28_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_28_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_28_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_28_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_28_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_28_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_28_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_28_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_28_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_28_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_28_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_28_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_28_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_28_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_28_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_28_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_28_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_28_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_28_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_28_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_28_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_28_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_28_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_28_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_28_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_28_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_28_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_28_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_28_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_28_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_28_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_28_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_28_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_28_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_28_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_28_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_28_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_28_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_28_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_28_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_28_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_28_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_28_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_28_bits_st_dep_mask <= _GEN_2069;
      ldq_28_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1809) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_28_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_28_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_28_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_28_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_28_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_28_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_28_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_28_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_28_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_28_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_28_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_28_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_28_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_28_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_28_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_28_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_28_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_28_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_28_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_28_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_28_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_28_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_28_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_28_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_28_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_28_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_28_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_28_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_28_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_28_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_28_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_28_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_28_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_28_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_28_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_28_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_28_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_28_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_28_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_28_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_28_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_28_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_28_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_28_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_28_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_28_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_28_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_28_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_28_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_28_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_28_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_28_bits_st_dep_mask <= _GEN_1685;
      ldq_28_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1617) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_28_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_28_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_28_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_28_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_28_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_28_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_28_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_28_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_28_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_28_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_28_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_28_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_28_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_28_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_28_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_28_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_28_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_28_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_28_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_28_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_28_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_28_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_28_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_28_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_28_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_28_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_28_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_28_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_28_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_28_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_28_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_28_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_28_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_28_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_28_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_28_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_28_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_28_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_28_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_28_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_28_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_28_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_28_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_28_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_28_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_28_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_28_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_28_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_28_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_28_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_28_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_28_bits_st_dep_mask <= next_live_store_mask;
      ldq_28_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_28_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_28_bits_st_dep_mask;
    if (ldq_28_valid)
      ldq_28_bits_uop_br_mask <= ldq_28_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2318)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2098)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1809)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1617)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2798) begin
      if (_exe_tlb_uop_T_9)
        ldq_28_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_28_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_28_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_28_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_28_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_28_bits_addr_bits <= casez_tmp_202;
        else
          ldq_28_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_28_bits_addr_bits <= _GEN_280;
      ldq_28_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_28_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2674) begin
      if (_exe_tlb_uop_T_2)
        ldq_28_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_28_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_28_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_28_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_28_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_28_bits_addr_bits <= casez_tmp_202;
        else
          ldq_28_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_28_bits_addr_bits <= _GEN_274;
      ldq_28_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_28_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2318)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2098)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1809)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1617)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_28_bits_addr_valid <= ~_GEN_5749 & _GEN_5649 & _GEN_5586 & _GEN_5491 & (_GEN_5336 ? ~_GEN_5268 & _GEN_2799 : ~_GEN_5364 & _GEN_2799);
    ldq_28_bits_executed <= ~_GEN_5749 & _GEN_5649 & _GEN_5586 & _GEN_5491 & _GEN_5396 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1502) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1463)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_363 & _GEN_5073 : ~(_GEN_1425 & _GEN_363) & _GEN_5073) : _GEN_5073) | (dis_ld_val_3 ? ~_GEN_2252 & _GEN_1873 : ~_GEN_2098 & _GEN_1873));
    ldq_28_bits_succeeded <= _GEN_5649 & _GEN_5586 & _GEN_5491 & _GEN_5396 & (_GEN_5201 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1C ? _ldq_bits_succeeded_T_1 : _GEN_5136 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1C ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2252 & _GEN_1905 : ~_GEN_2098 & _GEN_1905) : casez_tmp_490) : casez_tmp_524);
    ldq_28_bits_order_fail <= _GEN_5649 & _GEN_5586 & _GEN_5491 & _GEN_5396 & (_GEN_1001 ? _GEN_2960 : _GEN_1003 ? _GEN_1004 | _GEN_2960 : _GEN_1006 | _GEN_2960);
    ldq_28_bits_observed <= _GEN_1001 | _GEN_988 | (dis_ld_val_3 ? ~_GEN_2252 & _GEN_1969 : ~_GEN_2098 & _GEN_1969);
    ldq_28_bits_forward_std_val <= _GEN_5649 & _GEN_5586 & _GEN_5491 & _GEN_5396 & (~_GEN_1508 & _GEN_5200 | ~_GEN_1468 & _GEN_5135 | (dis_ld_val_3 ? ~_GEN_2252 & _GEN_2001 : ~_GEN_2098 & _GEN_2001));
    if (_GEN_5201) begin
      if (_GEN_5136) begin
      end
      else
        ldq_28_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_28_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_29_valid <= ~_GEN_5749 & _GEN_5650 & _GEN_5587 & _GEN_5492 & (_GEN_5336 ? ~_GEN_5269 & _GEN_2256 : ~_GEN_5365 & _GEN_2256);
    if (_GEN_2320) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_29_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_29_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_29_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_29_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_29_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_29_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_29_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_29_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_29_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_29_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_29_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_29_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_29_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_29_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_29_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_29_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_29_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_29_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_29_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_29_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_29_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_29_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_29_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_29_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_29_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_29_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_29_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_29_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_29_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_29_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_29_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_29_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_29_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_29_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_29_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_29_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_29_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_29_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_29_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_29_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_29_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_29_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_29_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_29_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_29_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_29_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_29_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_29_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_29_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_29_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_29_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_29_bits_st_dep_mask <= _GEN_2166;
      ldq_29_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2099) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_29_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_29_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_29_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_29_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_29_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_29_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_29_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_29_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_29_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_29_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_29_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_29_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_29_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_29_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_29_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_29_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_29_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_29_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_29_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_29_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_29_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_29_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_29_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_29_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_29_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_29_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_29_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_29_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_29_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_29_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_29_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_29_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_29_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_29_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_29_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_29_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_29_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_29_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_29_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_29_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_29_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_29_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_29_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_29_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_29_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_29_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_29_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_29_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_29_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_29_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_29_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_29_bits_st_dep_mask <= _GEN_2069;
      ldq_29_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1810) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_29_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_29_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_29_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_29_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_29_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_29_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_29_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_29_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_29_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_29_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_29_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_29_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_29_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_29_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_29_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_29_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_29_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_29_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_29_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_29_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_29_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_29_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_29_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_29_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_29_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_29_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_29_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_29_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_29_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_29_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_29_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_29_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_29_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_29_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_29_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_29_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_29_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_29_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_29_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_29_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_29_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_29_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_29_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_29_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_29_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_29_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_29_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_29_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_29_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_29_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_29_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_29_bits_st_dep_mask <= _GEN_1685;
      ldq_29_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1618) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_29_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_29_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_29_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_29_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_29_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_29_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_29_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_29_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_29_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_29_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_29_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_29_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_29_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_29_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_29_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_29_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_29_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_29_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_29_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_29_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_29_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_29_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_29_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_29_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_29_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_29_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_29_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_29_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_29_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_29_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_29_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_29_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_29_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_29_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_29_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_29_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_29_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_29_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_29_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_29_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_29_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_29_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_29_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_29_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_29_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_29_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_29_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_29_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_29_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_29_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_29_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_29_bits_st_dep_mask <= next_live_store_mask;
      ldq_29_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_29_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_29_bits_st_dep_mask;
    if (ldq_29_valid)
      ldq_29_bits_uop_br_mask <= ldq_29_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2320)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2099)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1810)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1618)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2800) begin
      if (_exe_tlb_uop_T_9)
        ldq_29_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_29_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_29_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_29_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_29_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_29_bits_addr_bits <= casez_tmp_202;
        else
          ldq_29_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_29_bits_addr_bits <= _GEN_280;
      ldq_29_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_29_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2675) begin
      if (_exe_tlb_uop_T_2)
        ldq_29_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_29_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_29_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_29_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_29_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_29_bits_addr_bits <= casez_tmp_202;
        else
          ldq_29_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_29_bits_addr_bits <= _GEN_274;
      ldq_29_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_29_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2320)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2099)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1810)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1618)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_29_bits_addr_valid <= ~_GEN_5749 & _GEN_5650 & _GEN_5587 & _GEN_5492 & (_GEN_5336 ? ~_GEN_5269 & _GEN_2801 : ~_GEN_5365 & _GEN_2801);
    ldq_29_bits_executed <= ~_GEN_5749 & _GEN_5650 & _GEN_5587 & _GEN_5492 & _GEN_5397 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1503) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1464)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_364 & _GEN_5074 : ~(_GEN_1425 & _GEN_364) & _GEN_5074) : _GEN_5074) | (dis_ld_val_3 ? ~_GEN_2255 & _GEN_1874 : ~_GEN_2099 & _GEN_1874));
    ldq_29_bits_succeeded <= _GEN_5650 & _GEN_5587 & _GEN_5492 & _GEN_5397 & (_GEN_5203 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1D ? _ldq_bits_succeeded_T_1 : _GEN_5138 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1D ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2255 & _GEN_1906 : ~_GEN_2099 & _GEN_1906) : casez_tmp_490) : casez_tmp_524);
    ldq_29_bits_order_fail <= _GEN_5650 & _GEN_5587 & _GEN_5492 & _GEN_5397 & (_GEN_1024 ? _GEN_2961 : _GEN_1026 ? _GEN_1027 | _GEN_2961 : _GEN_1029 | _GEN_2961);
    ldq_29_bits_observed <= _GEN_1024 | _GEN_1011 | (dis_ld_val_3 ? ~_GEN_2255 & _GEN_1970 : ~_GEN_2099 & _GEN_1970);
    ldq_29_bits_forward_std_val <= _GEN_5650 & _GEN_5587 & _GEN_5492 & _GEN_5397 & (~_GEN_1508 & _GEN_5202 | ~_GEN_1468 & _GEN_5137 | (dis_ld_val_3 ? ~_GEN_2255 & _GEN_2002 : ~_GEN_2099 & _GEN_2002));
    if (_GEN_5203) begin
      if (_GEN_5138) begin
      end
      else
        ldq_29_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_29_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_30_valid <= ~_GEN_5749 & _GEN_5651 & _GEN_5588 & _GEN_5493 & (_GEN_5336 ? ~_GEN_5270 & _GEN_2259 : ~_GEN_5366 & _GEN_2259);
    if (_GEN_2322) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_30_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_30_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_30_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_30_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_30_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_30_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_30_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_30_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_30_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_30_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_30_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_30_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_30_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_30_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_30_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_30_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_30_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_30_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_30_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_30_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_30_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_30_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_30_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_30_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_30_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_30_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_30_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_30_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_30_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_30_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_30_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_30_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_30_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_30_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_30_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_30_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_30_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_30_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_30_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_30_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_30_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_30_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_30_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_30_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_30_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_30_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_30_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_30_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_30_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_30_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_30_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_30_bits_st_dep_mask <= _GEN_2166;
      ldq_30_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2100) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_30_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_30_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_30_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_30_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_30_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_30_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_30_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_30_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_30_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_30_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_30_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_30_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_30_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_30_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_30_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_30_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_30_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_30_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_30_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_30_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_30_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_30_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_30_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_30_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_30_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_30_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_30_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_30_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_30_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_30_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_30_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_30_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_30_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_30_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_30_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_30_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_30_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_30_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_30_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_30_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_30_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_30_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_30_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_30_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_30_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_30_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_30_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_30_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_30_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_30_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_30_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_30_bits_st_dep_mask <= _GEN_2069;
      ldq_30_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1811) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_30_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_30_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_30_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_30_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_30_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_30_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_30_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_30_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_30_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_30_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_30_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_30_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_30_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_30_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_30_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_30_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_30_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_30_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_30_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_30_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_30_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_30_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_30_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_30_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_30_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_30_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_30_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_30_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_30_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_30_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_30_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_30_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_30_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_30_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_30_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_30_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_30_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_30_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_30_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_30_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_30_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_30_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_30_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_30_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_30_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_30_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_30_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_30_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_30_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_30_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_30_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_30_bits_st_dep_mask <= _GEN_1685;
      ldq_30_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1619) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_30_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_30_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_30_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_30_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_30_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_30_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_30_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_30_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_30_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_30_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_30_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_30_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_30_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_30_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_30_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_30_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_30_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_30_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_30_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_30_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_30_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_30_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_30_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_30_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_30_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_30_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_30_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_30_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_30_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_30_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_30_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_30_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_30_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_30_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_30_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_30_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_30_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_30_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_30_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_30_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_30_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_30_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_30_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_30_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_30_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_30_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_30_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_30_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_30_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_30_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_30_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_30_bits_st_dep_mask <= next_live_store_mask;
      ldq_30_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_30_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_30_bits_st_dep_mask;
    if (ldq_30_valid)
      ldq_30_bits_uop_br_mask <= ldq_30_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2322)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2100)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1811)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1619)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & _GEN_2802) begin
      if (_exe_tlb_uop_T_9)
        ldq_30_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_30_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_30_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_30_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_30_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_30_bits_addr_bits <= casez_tmp_202;
        else
          ldq_30_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_30_bits_addr_bits <= _GEN_280;
      ldq_30_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_30_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2676) begin
      if (_exe_tlb_uop_T_2)
        ldq_30_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_30_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_30_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_30_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_30_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_30_bits_addr_bits <= casez_tmp_202;
        else
          ldq_30_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_30_bits_addr_bits <= _GEN_274;
      ldq_30_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_30_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2322)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2100)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1811)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1619)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_30_bits_addr_valid <= ~_GEN_5749 & _GEN_5651 & _GEN_5588 & _GEN_5493 & (_GEN_5336 ? ~_GEN_5270 & _GEN_2803 : ~_GEN_5366 & _GEN_2803);
    ldq_30_bits_executed <= ~_GEN_5749 & _GEN_5651 & _GEN_5588 & _GEN_5493 & _GEN_5398 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1504) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_1465)) & ((_GEN_1426 ? (_GEN_5077 ? ~_GEN_365 & _GEN_5075 : ~(_GEN_1425 & _GEN_365) & _GEN_5075) : _GEN_5075) | (dis_ld_val_3 ? ~_GEN_2258 & _GEN_1875 : ~_GEN_2100 & _GEN_1875));
    ldq_30_bits_succeeded <= _GEN_5651 & _GEN_5588 & _GEN_5493 & _GEN_5398 & (_GEN_5205 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1E ? _ldq_bits_succeeded_T_1 : _GEN_5140 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1E ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2258 & _GEN_1907 : ~_GEN_2100 & _GEN_1907) : casez_tmp_490) : casez_tmp_524);
    ldq_30_bits_order_fail <= _GEN_5651 & _GEN_5588 & _GEN_5493 & _GEN_5398 & (_GEN_1047 ? _GEN_2962 : _GEN_1049 ? _GEN_1050 | _GEN_2962 : _GEN_1052 | _GEN_2962);
    ldq_30_bits_observed <= _GEN_1047 | _GEN_1034 | (dis_ld_val_3 ? ~_GEN_2258 & _GEN_1971 : ~_GEN_2100 & _GEN_1971);
    ldq_30_bits_forward_std_val <= _GEN_5651 & _GEN_5588 & _GEN_5493 & _GEN_5398 & (~_GEN_1508 & _GEN_5204 | ~_GEN_1468 & _GEN_5139 | (dis_ld_val_3 ? ~_GEN_2258 & _GEN_2003 : ~_GEN_2100 & _GEN_2003));
    if (_GEN_5205) begin
      if (_GEN_5140) begin
      end
      else
        ldq_30_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_30_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_31_valid <= ~_GEN_5749 & _GEN_5652 & _GEN_5589 & _GEN_5494 & (_GEN_5336 ? ~_GEN_5271 & _GEN_2261 : ~_GEN_5367 & _GEN_2261);
    if (_GEN_2324) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_31_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
      ldq_31_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
      ldq_31_bits_uop_is_rvc <= io_core_dis_uops_3_bits_is_rvc;
      ldq_31_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
      ldq_31_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
      ldq_31_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
      ldq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
      ldq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
      ldq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
      ldq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
      ldq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
      ldq_31_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_3_bits_ctrl_fcn_dw;
      ldq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_31_bits_uop_ctrl_is_std <= io_core_dis_uops_3_bits_ctrl_is_std;
      ldq_31_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      ldq_31_bits_uop_iw_p1_poisoned <= io_core_dis_uops_3_bits_iw_p1_poisoned;
      ldq_31_bits_uop_iw_p2_poisoned <= io_core_dis_uops_3_bits_iw_p2_poisoned;
      ldq_31_bits_uop_is_br <= io_core_dis_uops_3_bits_is_br;
      ldq_31_bits_uop_is_jalr <= io_core_dis_uops_3_bits_is_jalr;
      ldq_31_bits_uop_is_jal <= io_core_dis_uops_3_bits_is_jal;
      ldq_31_bits_uop_is_sfb <= io_core_dis_uops_3_bits_is_sfb;
      ldq_31_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
      ldq_31_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
      ldq_31_bits_uop_edge_inst <= io_core_dis_uops_3_bits_edge_inst;
      ldq_31_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
      ldq_31_bits_uop_taken <= io_core_dis_uops_3_bits_taken;
      ldq_31_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
      ldq_31_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_31_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      ldq_31_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
      ldq_31_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
      ldq_31_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      ldq_31_bits_uop_prs1_busy <= io_core_dis_uops_3_bits_prs1_busy;
      ldq_31_bits_uop_prs2_busy <= io_core_dis_uops_3_bits_prs2_busy;
      ldq_31_bits_uop_prs3_busy <= io_core_dis_uops_3_bits_prs3_busy;
      ldq_31_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
      ldq_31_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
      ldq_31_bits_uop_bypassable <= io_core_dis_uops_3_bits_bypassable;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
      ldq_31_bits_uop_is_fencei <= io_core_dis_uops_3_bits_is_fencei;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_31_bits_uop_is_sys_pc2epc <= io_core_dis_uops_3_bits_is_sys_pc2epc;
      ldq_31_bits_uop_is_unique <= io_core_dis_uops_3_bits_is_unique;
      ldq_31_bits_uop_flush_on_commit <= io_core_dis_uops_3_bits_flush_on_commit;
      ldq_31_bits_uop_ldst_is_rs1 <= io_core_dis_uops_3_bits_ldst_is_rs1;
      ldq_31_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
      ldq_31_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
      ldq_31_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
      ldq_31_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
      ldq_31_bits_uop_ldst_val <= io_core_dis_uops_3_bits_ldst_val;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
      ldq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
      ldq_31_bits_uop_frs3_en <= io_core_dis_uops_3_bits_frs3_en;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_31_bits_uop_fp_single <= io_core_dis_uops_3_bits_fp_single;
      ldq_31_bits_uop_xcpt_pf_if <= io_core_dis_uops_3_bits_xcpt_pf_if;
      ldq_31_bits_uop_xcpt_ae_if <= io_core_dis_uops_3_bits_xcpt_ae_if;
      ldq_31_bits_uop_xcpt_ma_if <= io_core_dis_uops_3_bits_xcpt_ma_if;
      ldq_31_bits_uop_bp_debug_if <= io_core_dis_uops_3_bits_bp_debug_if;
      ldq_31_bits_uop_bp_xcpt_if <= io_core_dis_uops_3_bits_bp_xcpt_if;
      ldq_31_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
      ldq_31_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      ldq_31_bits_st_dep_mask <= _GEN_2166;
      ldq_31_bits_youngest_stq_idx <= _GEN_14;
    end
    else if (_GEN_2101) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_31_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
      ldq_31_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
      ldq_31_bits_uop_is_rvc <= io_core_dis_uops_2_bits_is_rvc;
      ldq_31_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
      ldq_31_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
      ldq_31_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
      ldq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
      ldq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
      ldq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
      ldq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
      ldq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
      ldq_31_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_2_bits_ctrl_fcn_dw;
      ldq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_31_bits_uop_ctrl_is_std <= io_core_dis_uops_2_bits_ctrl_is_std;
      ldq_31_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
      ldq_31_bits_uop_iw_p1_poisoned <= io_core_dis_uops_2_bits_iw_p1_poisoned;
      ldq_31_bits_uop_iw_p2_poisoned <= io_core_dis_uops_2_bits_iw_p2_poisoned;
      ldq_31_bits_uop_is_br <= io_core_dis_uops_2_bits_is_br;
      ldq_31_bits_uop_is_jalr <= io_core_dis_uops_2_bits_is_jalr;
      ldq_31_bits_uop_is_jal <= io_core_dis_uops_2_bits_is_jal;
      ldq_31_bits_uop_is_sfb <= io_core_dis_uops_2_bits_is_sfb;
      ldq_31_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
      ldq_31_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
      ldq_31_bits_uop_edge_inst <= io_core_dis_uops_2_bits_edge_inst;
      ldq_31_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
      ldq_31_bits_uop_taken <= io_core_dis_uops_2_bits_taken;
      ldq_31_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
      ldq_31_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_31_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
      ldq_31_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
      ldq_31_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
      ldq_31_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
      ldq_31_bits_uop_prs1_busy <= io_core_dis_uops_2_bits_prs1_busy;
      ldq_31_bits_uop_prs2_busy <= io_core_dis_uops_2_bits_prs2_busy;
      ldq_31_bits_uop_prs3_busy <= io_core_dis_uops_2_bits_prs3_busy;
      ldq_31_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
      ldq_31_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
      ldq_31_bits_uop_bypassable <= io_core_dis_uops_2_bits_bypassable;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
      ldq_31_bits_uop_is_fencei <= io_core_dis_uops_2_bits_is_fencei;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_31_bits_uop_is_sys_pc2epc <= io_core_dis_uops_2_bits_is_sys_pc2epc;
      ldq_31_bits_uop_is_unique <= io_core_dis_uops_2_bits_is_unique;
      ldq_31_bits_uop_flush_on_commit <= io_core_dis_uops_2_bits_flush_on_commit;
      ldq_31_bits_uop_ldst_is_rs1 <= io_core_dis_uops_2_bits_ldst_is_rs1;
      ldq_31_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
      ldq_31_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
      ldq_31_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
      ldq_31_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
      ldq_31_bits_uop_ldst_val <= io_core_dis_uops_2_bits_ldst_val;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
      ldq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
      ldq_31_bits_uop_frs3_en <= io_core_dis_uops_2_bits_frs3_en;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_31_bits_uop_fp_single <= io_core_dis_uops_2_bits_fp_single;
      ldq_31_bits_uop_xcpt_pf_if <= io_core_dis_uops_2_bits_xcpt_pf_if;
      ldq_31_bits_uop_xcpt_ae_if <= io_core_dis_uops_2_bits_xcpt_ae_if;
      ldq_31_bits_uop_xcpt_ma_if <= io_core_dis_uops_2_bits_xcpt_ma_if;
      ldq_31_bits_uop_bp_debug_if <= io_core_dis_uops_2_bits_bp_debug_if;
      ldq_31_bits_uop_bp_xcpt_if <= io_core_dis_uops_2_bits_bp_xcpt_if;
      ldq_31_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
      ldq_31_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
      ldq_31_bits_st_dep_mask <= _GEN_2069;
      ldq_31_bits_youngest_stq_idx <= _GEN_10;
    end
    else if (_GEN_1812) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_31_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
      ldq_31_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
      ldq_31_bits_uop_is_rvc <= io_core_dis_uops_1_bits_is_rvc;
      ldq_31_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
      ldq_31_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
      ldq_31_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
      ldq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
      ldq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
      ldq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
      ldq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
      ldq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
      ldq_31_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_1_bits_ctrl_fcn_dw;
      ldq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_31_bits_uop_ctrl_is_std <= io_core_dis_uops_1_bits_ctrl_is_std;
      ldq_31_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
      ldq_31_bits_uop_iw_p1_poisoned <= io_core_dis_uops_1_bits_iw_p1_poisoned;
      ldq_31_bits_uop_iw_p2_poisoned <= io_core_dis_uops_1_bits_iw_p2_poisoned;
      ldq_31_bits_uop_is_br <= io_core_dis_uops_1_bits_is_br;
      ldq_31_bits_uop_is_jalr <= io_core_dis_uops_1_bits_is_jalr;
      ldq_31_bits_uop_is_jal <= io_core_dis_uops_1_bits_is_jal;
      ldq_31_bits_uop_is_sfb <= io_core_dis_uops_1_bits_is_sfb;
      ldq_31_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
      ldq_31_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
      ldq_31_bits_uop_edge_inst <= io_core_dis_uops_1_bits_edge_inst;
      ldq_31_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
      ldq_31_bits_uop_taken <= io_core_dis_uops_1_bits_taken;
      ldq_31_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
      ldq_31_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_31_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
      ldq_31_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
      ldq_31_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
      ldq_31_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
      ldq_31_bits_uop_prs1_busy <= io_core_dis_uops_1_bits_prs1_busy;
      ldq_31_bits_uop_prs2_busy <= io_core_dis_uops_1_bits_prs2_busy;
      ldq_31_bits_uop_prs3_busy <= io_core_dis_uops_1_bits_prs3_busy;
      ldq_31_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
      ldq_31_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
      ldq_31_bits_uop_bypassable <= io_core_dis_uops_1_bits_bypassable;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
      ldq_31_bits_uop_is_fencei <= io_core_dis_uops_1_bits_is_fencei;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_31_bits_uop_is_sys_pc2epc <= io_core_dis_uops_1_bits_is_sys_pc2epc;
      ldq_31_bits_uop_is_unique <= io_core_dis_uops_1_bits_is_unique;
      ldq_31_bits_uop_flush_on_commit <= io_core_dis_uops_1_bits_flush_on_commit;
      ldq_31_bits_uop_ldst_is_rs1 <= io_core_dis_uops_1_bits_ldst_is_rs1;
      ldq_31_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
      ldq_31_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
      ldq_31_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
      ldq_31_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
      ldq_31_bits_uop_ldst_val <= io_core_dis_uops_1_bits_ldst_val;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
      ldq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
      ldq_31_bits_uop_frs3_en <= io_core_dis_uops_1_bits_frs3_en;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_31_bits_uop_fp_single <= io_core_dis_uops_1_bits_fp_single;
      ldq_31_bits_uop_xcpt_pf_if <= io_core_dis_uops_1_bits_xcpt_pf_if;
      ldq_31_bits_uop_xcpt_ae_if <= io_core_dis_uops_1_bits_xcpt_ae_if;
      ldq_31_bits_uop_xcpt_ma_if <= io_core_dis_uops_1_bits_xcpt_ma_if;
      ldq_31_bits_uop_bp_debug_if <= io_core_dis_uops_1_bits_bp_debug_if;
      ldq_31_bits_uop_bp_xcpt_if <= io_core_dis_uops_1_bits_bp_xcpt_if;
      ldq_31_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
      ldq_31_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
      ldq_31_bits_st_dep_mask <= _GEN_1685;
      ldq_31_bits_youngest_stq_idx <= _GEN_6;
    end
    else if (_GEN_1620) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_31_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
      ldq_31_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
      ldq_31_bits_uop_is_rvc <= io_core_dis_uops_0_bits_is_rvc;
      ldq_31_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
      ldq_31_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
      ldq_31_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
      ldq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
      ldq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
      ldq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
      ldq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
      ldq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
      ldq_31_bits_uop_ctrl_fcn_dw <= io_core_dis_uops_0_bits_ctrl_fcn_dw;
      ldq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_31_bits_uop_ctrl_is_std <= io_core_dis_uops_0_bits_ctrl_is_std;
      ldq_31_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
      ldq_31_bits_uop_iw_p1_poisoned <= io_core_dis_uops_0_bits_iw_p1_poisoned;
      ldq_31_bits_uop_iw_p2_poisoned <= io_core_dis_uops_0_bits_iw_p2_poisoned;
      ldq_31_bits_uop_is_br <= io_core_dis_uops_0_bits_is_br;
      ldq_31_bits_uop_is_jalr <= io_core_dis_uops_0_bits_is_jalr;
      ldq_31_bits_uop_is_jal <= io_core_dis_uops_0_bits_is_jal;
      ldq_31_bits_uop_is_sfb <= io_core_dis_uops_0_bits_is_sfb;
      ldq_31_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
      ldq_31_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
      ldq_31_bits_uop_edge_inst <= io_core_dis_uops_0_bits_edge_inst;
      ldq_31_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
      ldq_31_bits_uop_taken <= io_core_dis_uops_0_bits_taken;
      ldq_31_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
      ldq_31_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_31_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
      ldq_31_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
      ldq_31_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
      ldq_31_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
      ldq_31_bits_uop_prs1_busy <= io_core_dis_uops_0_bits_prs1_busy;
      ldq_31_bits_uop_prs2_busy <= io_core_dis_uops_0_bits_prs2_busy;
      ldq_31_bits_uop_prs3_busy <= io_core_dis_uops_0_bits_prs3_busy;
      ldq_31_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
      ldq_31_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
      ldq_31_bits_uop_bypassable <= io_core_dis_uops_0_bits_bypassable;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
      ldq_31_bits_uop_is_fencei <= io_core_dis_uops_0_bits_is_fencei;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_31_bits_uop_is_sys_pc2epc <= io_core_dis_uops_0_bits_is_sys_pc2epc;
      ldq_31_bits_uop_is_unique <= io_core_dis_uops_0_bits_is_unique;
      ldq_31_bits_uop_flush_on_commit <= io_core_dis_uops_0_bits_flush_on_commit;
      ldq_31_bits_uop_ldst_is_rs1 <= io_core_dis_uops_0_bits_ldst_is_rs1;
      ldq_31_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
      ldq_31_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
      ldq_31_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
      ldq_31_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
      ldq_31_bits_uop_ldst_val <= io_core_dis_uops_0_bits_ldst_val;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
      ldq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
      ldq_31_bits_uop_frs3_en <= io_core_dis_uops_0_bits_frs3_en;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_31_bits_uop_fp_single <= io_core_dis_uops_0_bits_fp_single;
      ldq_31_bits_uop_xcpt_pf_if <= io_core_dis_uops_0_bits_xcpt_pf_if;
      ldq_31_bits_uop_xcpt_ae_if <= io_core_dis_uops_0_bits_xcpt_ae_if;
      ldq_31_bits_uop_xcpt_ma_if <= io_core_dis_uops_0_bits_xcpt_ma_if;
      ldq_31_bits_uop_bp_debug_if <= io_core_dis_uops_0_bits_bp_debug_if;
      ldq_31_bits_uop_bp_xcpt_if <= io_core_dis_uops_0_bits_bp_xcpt_if;
      ldq_31_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
      ldq_31_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
      ldq_31_bits_st_dep_mask <= next_live_store_mask;
      ldq_31_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_31_bits_st_dep_mask <= (_GEN_1588 | ~_ldq_31_bits_st_dep_mask_T) & ldq_31_bits_st_dep_mask;
    if (ldq_31_valid)
      ldq_31_bits_uop_br_mask <= ldq_31_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_2324)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_2101)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_1812)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_1620)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_281 & (&ldq_idx_1)) begin
      if (_exe_tlb_uop_T_9)
        ldq_31_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
      else if (will_fire_load_retry_1_will_fire)
        ldq_31_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_31_bits_uop_pdst <= _exe_tlb_uop_T_11_pdst;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          ldq_31_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          ldq_31_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          ldq_31_bits_addr_bits <= casez_tmp_202;
        else
          ldq_31_bits_addr_bits <= _exe_tlb_vaddr_T_10;
      end
      else
        ldq_31_bits_addr_bits <= _GEN_280;
      ldq_31_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_31_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_3;
    end
    else if (_GEN_2677) begin
      if (_exe_tlb_uop_T_2)
        ldq_31_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
      else if (will_fire_load_retry_0_will_fire)
        ldq_31_bits_uop_pdst <= casez_tmp_160;
      else
        ldq_31_bits_uop_pdst <= _exe_tlb_uop_T_4_pdst;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          ldq_31_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          ldq_31_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          ldq_31_bits_addr_bits <= casez_tmp_202;
        else
          ldq_31_bits_addr_bits <= _exe_tlb_vaddr_T_3;
      end
      else
        ldq_31_bits_addr_bits <= _GEN_274;
      ldq_31_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_31_bits_addr_is_uncacheable <= _ldq_bits_addr_is_uncacheable_T_1;
    end
    else if (_GEN_2324)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_2101)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_1812)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_1620)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_31_bits_addr_valid <= ~_GEN_5749 & _GEN_5652 & _GEN_5589 & _GEN_5494 & (_GEN_5336 ? ~_GEN_5271 & _GEN_2804 : ~_GEN_5367 & _GEN_2804);
    ldq_31_bits_executed <= ~_GEN_5749 & _GEN_5652 & _GEN_5589 & _GEN_5494 & _GEN_5399 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_1505) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & (&io_dmem_nack_0_bits_uop_ldq_idx))) & ((_GEN_1426 ? (_GEN_5077 ? ~(&lcam_ldq_idx_1) & _GEN_5076 : ~(_GEN_1425 & (&lcam_ldq_idx_1)) & _GEN_5076) : _GEN_5076) | (dis_ld_val_3 ? ~_GEN_2260 & _GEN_1876 : ~_GEN_2101 & _GEN_1876));
    ldq_31_bits_succeeded <= _GEN_5652 & _GEN_5589 & _GEN_5494 & _GEN_5399 & (_GEN_5207 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & (&io_dmem_resp_1_bits_uop_ldq_idx) ? _ldq_bits_succeeded_T_1 : _GEN_5142 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & (&io_dmem_resp_0_bits_uop_ldq_idx) ? _ldq_bits_succeeded_T : dis_ld_val_3 ? ~_GEN_2260 & _GEN_1908 : ~_GEN_2101 & _GEN_1908) : casez_tmp_490) : casez_tmp_524);
    ldq_31_bits_order_fail <= _GEN_5652 & _GEN_5589 & _GEN_5494 & _GEN_5399 & (_GEN_1070 ? _GEN_2964 : _GEN_1072 ? _GEN_1073 | _GEN_2964 : _GEN_1075 | _GEN_2964);
    ldq_31_bits_observed <= _GEN_1070 | _GEN_1057 | (dis_ld_val_3 ? ~_GEN_2260 & _GEN_1972 : ~_GEN_2101 & _GEN_1972);
    ldq_31_bits_forward_std_val <= _GEN_5652 & _GEN_5589 & _GEN_5494 & _GEN_5399 & (~_GEN_1508 & _GEN_5206 | ~_GEN_1468 & _GEN_5141 | (dis_ld_val_3 ? ~_GEN_2260 & _GEN_2004 : ~_GEN_2101 & _GEN_2004));
    if (_GEN_5207) begin
      if (_GEN_5142) begin
      end
      else
        ldq_31_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_31_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    stq_0_valid <= ~_GEN_5752 & (clear_store ? ~_GEN_5654 & _GEN_2391 : ~_GEN_5208 & _GEN_2391);
    if (_GEN_5750) begin
      stq_0_bits_uop_uopc <= 7'h0;
      stq_0_bits_uop_inst <= 32'h0;
      stq_0_bits_uop_debug_inst <= 32'h0;
      stq_0_bits_uop_debug_pc <= 40'h0;
      stq_0_bits_uop_iq_type <= 3'h0;
      stq_0_bits_uop_fu_code <= 10'h0;
      stq_0_bits_uop_ctrl_br_type <= 4'h0;
      stq_0_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_0_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_0_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_0_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_0_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_0_bits_uop_iw_state <= 2'h0;
      stq_0_bits_uop_br_mask <= 20'h0;
      stq_0_bits_uop_br_tag <= 5'h0;
      stq_0_bits_uop_ftq_idx <= 6'h0;
      stq_0_bits_uop_pc_lob <= 6'h0;
      stq_0_bits_uop_imm_packed <= 20'h0;
      stq_0_bits_uop_csr_addr <= 12'h0;
      stq_0_bits_uop_rob_idx <= 7'h0;
      stq_0_bits_uop_ldq_idx <= 5'h0;
      stq_0_bits_uop_stq_idx <= 5'h0;
      stq_0_bits_uop_rxq_idx <= 2'h0;
      stq_0_bits_uop_pdst <= 7'h0;
      stq_0_bits_uop_prs1 <= 7'h0;
      stq_0_bits_uop_prs2 <= 7'h0;
      stq_0_bits_uop_prs3 <= 7'h0;
      stq_0_bits_uop_ppred <= 6'h0;
      stq_0_bits_uop_stale_pdst <= 7'h0;
      stq_0_bits_uop_exc_cause <= 64'h0;
      stq_0_bits_uop_mem_cmd <= 5'h0;
      stq_0_bits_uop_mem_size <= 2'h0;
      stq_0_bits_uop_ldst <= 6'h0;
      stq_0_bits_uop_lrs1 <= 6'h0;
      stq_0_bits_uop_lrs2 <= 6'h0;
      stq_0_bits_uop_lrs3 <= 6'h0;
      stq_0_bits_uop_dst_rtype <= 2'h2;
      stq_0_bits_uop_lrs1_rtype <= 2'h0;
      stq_0_bits_uop_lrs2_rtype <= 2'h0;
      stq_0_bits_uop_debug_fsrc <= 2'h0;
      stq_0_bits_uop_debug_tsrc <= 2'h0;
      stq_1_bits_uop_uopc <= 7'h0;
      stq_1_bits_uop_inst <= 32'h0;
      stq_1_bits_uop_debug_inst <= 32'h0;
      stq_1_bits_uop_debug_pc <= 40'h0;
      stq_1_bits_uop_iq_type <= 3'h0;
      stq_1_bits_uop_fu_code <= 10'h0;
      stq_1_bits_uop_ctrl_br_type <= 4'h0;
      stq_1_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_1_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_1_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_1_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_1_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_1_bits_uop_iw_state <= 2'h0;
      stq_1_bits_uop_br_mask <= 20'h0;
      stq_1_bits_uop_br_tag <= 5'h0;
      stq_1_bits_uop_ftq_idx <= 6'h0;
      stq_1_bits_uop_pc_lob <= 6'h0;
      stq_1_bits_uop_imm_packed <= 20'h0;
      stq_1_bits_uop_csr_addr <= 12'h0;
      stq_1_bits_uop_rob_idx <= 7'h0;
      stq_1_bits_uop_ldq_idx <= 5'h0;
      stq_1_bits_uop_stq_idx <= 5'h0;
      stq_1_bits_uop_rxq_idx <= 2'h0;
      stq_1_bits_uop_pdst <= 7'h0;
      stq_1_bits_uop_prs1 <= 7'h0;
      stq_1_bits_uop_prs2 <= 7'h0;
      stq_1_bits_uop_prs3 <= 7'h0;
      stq_1_bits_uop_ppred <= 6'h0;
      stq_1_bits_uop_stale_pdst <= 7'h0;
      stq_1_bits_uop_exc_cause <= 64'h0;
      stq_1_bits_uop_mem_cmd <= 5'h0;
      stq_1_bits_uop_mem_size <= 2'h0;
      stq_1_bits_uop_ldst <= 6'h0;
      stq_1_bits_uop_lrs1 <= 6'h0;
      stq_1_bits_uop_lrs2 <= 6'h0;
      stq_1_bits_uop_lrs3 <= 6'h0;
      stq_1_bits_uop_dst_rtype <= 2'h2;
      stq_1_bits_uop_lrs1_rtype <= 2'h0;
      stq_1_bits_uop_lrs2_rtype <= 2'h0;
      stq_1_bits_uop_debug_fsrc <= 2'h0;
      stq_1_bits_uop_debug_tsrc <= 2'h0;
      stq_2_bits_uop_uopc <= 7'h0;
      stq_2_bits_uop_inst <= 32'h0;
      stq_2_bits_uop_debug_inst <= 32'h0;
      stq_2_bits_uop_debug_pc <= 40'h0;
      stq_2_bits_uop_iq_type <= 3'h0;
      stq_2_bits_uop_fu_code <= 10'h0;
      stq_2_bits_uop_ctrl_br_type <= 4'h0;
      stq_2_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_2_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_2_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_2_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_2_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_2_bits_uop_iw_state <= 2'h0;
      stq_2_bits_uop_br_mask <= 20'h0;
      stq_2_bits_uop_br_tag <= 5'h0;
      stq_2_bits_uop_ftq_idx <= 6'h0;
      stq_2_bits_uop_pc_lob <= 6'h0;
      stq_2_bits_uop_imm_packed <= 20'h0;
      stq_2_bits_uop_csr_addr <= 12'h0;
      stq_2_bits_uop_rob_idx <= 7'h0;
      stq_2_bits_uop_ldq_idx <= 5'h0;
      stq_2_bits_uop_stq_idx <= 5'h0;
      stq_2_bits_uop_rxq_idx <= 2'h0;
      stq_2_bits_uop_pdst <= 7'h0;
      stq_2_bits_uop_prs1 <= 7'h0;
      stq_2_bits_uop_prs2 <= 7'h0;
      stq_2_bits_uop_prs3 <= 7'h0;
      stq_2_bits_uop_ppred <= 6'h0;
      stq_2_bits_uop_stale_pdst <= 7'h0;
      stq_2_bits_uop_exc_cause <= 64'h0;
      stq_2_bits_uop_mem_cmd <= 5'h0;
      stq_2_bits_uop_mem_size <= 2'h0;
      stq_2_bits_uop_ldst <= 6'h0;
      stq_2_bits_uop_lrs1 <= 6'h0;
      stq_2_bits_uop_lrs2 <= 6'h0;
      stq_2_bits_uop_lrs3 <= 6'h0;
      stq_2_bits_uop_dst_rtype <= 2'h2;
      stq_2_bits_uop_lrs1_rtype <= 2'h0;
      stq_2_bits_uop_lrs2_rtype <= 2'h0;
      stq_2_bits_uop_debug_fsrc <= 2'h0;
      stq_2_bits_uop_debug_tsrc <= 2'h0;
      stq_3_bits_uop_uopc <= 7'h0;
      stq_3_bits_uop_inst <= 32'h0;
      stq_3_bits_uop_debug_inst <= 32'h0;
      stq_3_bits_uop_debug_pc <= 40'h0;
      stq_3_bits_uop_iq_type <= 3'h0;
      stq_3_bits_uop_fu_code <= 10'h0;
      stq_3_bits_uop_ctrl_br_type <= 4'h0;
      stq_3_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_3_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_3_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_3_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_3_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_3_bits_uop_iw_state <= 2'h0;
      stq_3_bits_uop_br_mask <= 20'h0;
      stq_3_bits_uop_br_tag <= 5'h0;
      stq_3_bits_uop_ftq_idx <= 6'h0;
      stq_3_bits_uop_pc_lob <= 6'h0;
      stq_3_bits_uop_imm_packed <= 20'h0;
      stq_3_bits_uop_csr_addr <= 12'h0;
      stq_3_bits_uop_rob_idx <= 7'h0;
      stq_3_bits_uop_ldq_idx <= 5'h0;
      stq_3_bits_uop_stq_idx <= 5'h0;
      stq_3_bits_uop_rxq_idx <= 2'h0;
      stq_3_bits_uop_pdst <= 7'h0;
      stq_3_bits_uop_prs1 <= 7'h0;
      stq_3_bits_uop_prs2 <= 7'h0;
      stq_3_bits_uop_prs3 <= 7'h0;
      stq_3_bits_uop_ppred <= 6'h0;
      stq_3_bits_uop_stale_pdst <= 7'h0;
      stq_3_bits_uop_exc_cause <= 64'h0;
      stq_3_bits_uop_mem_cmd <= 5'h0;
      stq_3_bits_uop_mem_size <= 2'h0;
      stq_3_bits_uop_ldst <= 6'h0;
      stq_3_bits_uop_lrs1 <= 6'h0;
      stq_3_bits_uop_lrs2 <= 6'h0;
      stq_3_bits_uop_lrs3 <= 6'h0;
      stq_3_bits_uop_dst_rtype <= 2'h2;
      stq_3_bits_uop_lrs1_rtype <= 2'h0;
      stq_3_bits_uop_lrs2_rtype <= 2'h0;
      stq_3_bits_uop_debug_fsrc <= 2'h0;
      stq_3_bits_uop_debug_tsrc <= 2'h0;
      stq_4_bits_uop_uopc <= 7'h0;
      stq_4_bits_uop_inst <= 32'h0;
      stq_4_bits_uop_debug_inst <= 32'h0;
      stq_4_bits_uop_debug_pc <= 40'h0;
      stq_4_bits_uop_iq_type <= 3'h0;
      stq_4_bits_uop_fu_code <= 10'h0;
      stq_4_bits_uop_ctrl_br_type <= 4'h0;
      stq_4_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_4_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_4_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_4_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_4_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_4_bits_uop_iw_state <= 2'h0;
      stq_4_bits_uop_br_mask <= 20'h0;
      stq_4_bits_uop_br_tag <= 5'h0;
      stq_4_bits_uop_ftq_idx <= 6'h0;
      stq_4_bits_uop_pc_lob <= 6'h0;
      stq_4_bits_uop_imm_packed <= 20'h0;
      stq_4_bits_uop_csr_addr <= 12'h0;
      stq_4_bits_uop_rob_idx <= 7'h0;
      stq_4_bits_uop_ldq_idx <= 5'h0;
      stq_4_bits_uop_stq_idx <= 5'h0;
      stq_4_bits_uop_rxq_idx <= 2'h0;
      stq_4_bits_uop_pdst <= 7'h0;
      stq_4_bits_uop_prs1 <= 7'h0;
      stq_4_bits_uop_prs2 <= 7'h0;
      stq_4_bits_uop_prs3 <= 7'h0;
      stq_4_bits_uop_ppred <= 6'h0;
      stq_4_bits_uop_stale_pdst <= 7'h0;
      stq_4_bits_uop_exc_cause <= 64'h0;
      stq_4_bits_uop_mem_cmd <= 5'h0;
      stq_4_bits_uop_mem_size <= 2'h0;
      stq_4_bits_uop_ldst <= 6'h0;
      stq_4_bits_uop_lrs1 <= 6'h0;
      stq_4_bits_uop_lrs2 <= 6'h0;
      stq_4_bits_uop_lrs3 <= 6'h0;
      stq_4_bits_uop_dst_rtype <= 2'h2;
      stq_4_bits_uop_lrs1_rtype <= 2'h0;
      stq_4_bits_uop_lrs2_rtype <= 2'h0;
      stq_4_bits_uop_debug_fsrc <= 2'h0;
      stq_4_bits_uop_debug_tsrc <= 2'h0;
      stq_5_bits_uop_uopc <= 7'h0;
      stq_5_bits_uop_inst <= 32'h0;
      stq_5_bits_uop_debug_inst <= 32'h0;
      stq_5_bits_uop_debug_pc <= 40'h0;
      stq_5_bits_uop_iq_type <= 3'h0;
      stq_5_bits_uop_fu_code <= 10'h0;
      stq_5_bits_uop_ctrl_br_type <= 4'h0;
      stq_5_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_5_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_5_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_5_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_5_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_5_bits_uop_iw_state <= 2'h0;
      stq_5_bits_uop_br_mask <= 20'h0;
      stq_5_bits_uop_br_tag <= 5'h0;
      stq_5_bits_uop_ftq_idx <= 6'h0;
      stq_5_bits_uop_pc_lob <= 6'h0;
      stq_5_bits_uop_imm_packed <= 20'h0;
      stq_5_bits_uop_csr_addr <= 12'h0;
      stq_5_bits_uop_rob_idx <= 7'h0;
      stq_5_bits_uop_ldq_idx <= 5'h0;
      stq_5_bits_uop_stq_idx <= 5'h0;
      stq_5_bits_uop_rxq_idx <= 2'h0;
      stq_5_bits_uop_pdst <= 7'h0;
      stq_5_bits_uop_prs1 <= 7'h0;
      stq_5_bits_uop_prs2 <= 7'h0;
      stq_5_bits_uop_prs3 <= 7'h0;
      stq_5_bits_uop_ppred <= 6'h0;
      stq_5_bits_uop_stale_pdst <= 7'h0;
      stq_5_bits_uop_exc_cause <= 64'h0;
      stq_5_bits_uop_mem_cmd <= 5'h0;
      stq_5_bits_uop_mem_size <= 2'h0;
      stq_5_bits_uop_ldst <= 6'h0;
      stq_5_bits_uop_lrs1 <= 6'h0;
      stq_5_bits_uop_lrs2 <= 6'h0;
      stq_5_bits_uop_lrs3 <= 6'h0;
      stq_5_bits_uop_dst_rtype <= 2'h2;
      stq_5_bits_uop_lrs1_rtype <= 2'h0;
      stq_5_bits_uop_lrs2_rtype <= 2'h0;
      stq_5_bits_uop_debug_fsrc <= 2'h0;
      stq_5_bits_uop_debug_tsrc <= 2'h0;
      stq_6_bits_uop_uopc <= 7'h0;
      stq_6_bits_uop_inst <= 32'h0;
      stq_6_bits_uop_debug_inst <= 32'h0;
      stq_6_bits_uop_debug_pc <= 40'h0;
      stq_6_bits_uop_iq_type <= 3'h0;
      stq_6_bits_uop_fu_code <= 10'h0;
      stq_6_bits_uop_ctrl_br_type <= 4'h0;
      stq_6_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_6_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_6_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_6_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_6_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_6_bits_uop_iw_state <= 2'h0;
      stq_6_bits_uop_br_mask <= 20'h0;
      stq_6_bits_uop_br_tag <= 5'h0;
      stq_6_bits_uop_ftq_idx <= 6'h0;
      stq_6_bits_uop_pc_lob <= 6'h0;
      stq_6_bits_uop_imm_packed <= 20'h0;
      stq_6_bits_uop_csr_addr <= 12'h0;
      stq_6_bits_uop_rob_idx <= 7'h0;
      stq_6_bits_uop_ldq_idx <= 5'h0;
      stq_6_bits_uop_stq_idx <= 5'h0;
      stq_6_bits_uop_rxq_idx <= 2'h0;
      stq_6_bits_uop_pdst <= 7'h0;
      stq_6_bits_uop_prs1 <= 7'h0;
      stq_6_bits_uop_prs2 <= 7'h0;
      stq_6_bits_uop_prs3 <= 7'h0;
      stq_6_bits_uop_ppred <= 6'h0;
      stq_6_bits_uop_stale_pdst <= 7'h0;
      stq_6_bits_uop_exc_cause <= 64'h0;
      stq_6_bits_uop_mem_cmd <= 5'h0;
      stq_6_bits_uop_mem_size <= 2'h0;
      stq_6_bits_uop_ldst <= 6'h0;
      stq_6_bits_uop_lrs1 <= 6'h0;
      stq_6_bits_uop_lrs2 <= 6'h0;
      stq_6_bits_uop_lrs3 <= 6'h0;
      stq_6_bits_uop_dst_rtype <= 2'h2;
      stq_6_bits_uop_lrs1_rtype <= 2'h0;
      stq_6_bits_uop_lrs2_rtype <= 2'h0;
      stq_6_bits_uop_debug_fsrc <= 2'h0;
      stq_6_bits_uop_debug_tsrc <= 2'h0;
      stq_7_bits_uop_uopc <= 7'h0;
      stq_7_bits_uop_inst <= 32'h0;
      stq_7_bits_uop_debug_inst <= 32'h0;
      stq_7_bits_uop_debug_pc <= 40'h0;
      stq_7_bits_uop_iq_type <= 3'h0;
      stq_7_bits_uop_fu_code <= 10'h0;
      stq_7_bits_uop_ctrl_br_type <= 4'h0;
      stq_7_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_7_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_7_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_7_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_7_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_7_bits_uop_iw_state <= 2'h0;
      stq_7_bits_uop_br_mask <= 20'h0;
      stq_7_bits_uop_br_tag <= 5'h0;
      stq_7_bits_uop_ftq_idx <= 6'h0;
      stq_7_bits_uop_pc_lob <= 6'h0;
      stq_7_bits_uop_imm_packed <= 20'h0;
      stq_7_bits_uop_csr_addr <= 12'h0;
      stq_7_bits_uop_rob_idx <= 7'h0;
      stq_7_bits_uop_ldq_idx <= 5'h0;
      stq_7_bits_uop_stq_idx <= 5'h0;
      stq_7_bits_uop_rxq_idx <= 2'h0;
      stq_7_bits_uop_pdst <= 7'h0;
      stq_7_bits_uop_prs1 <= 7'h0;
      stq_7_bits_uop_prs2 <= 7'h0;
      stq_7_bits_uop_prs3 <= 7'h0;
      stq_7_bits_uop_ppred <= 6'h0;
      stq_7_bits_uop_stale_pdst <= 7'h0;
      stq_7_bits_uop_exc_cause <= 64'h0;
      stq_7_bits_uop_mem_cmd <= 5'h0;
      stq_7_bits_uop_mem_size <= 2'h0;
      stq_7_bits_uop_ldst <= 6'h0;
      stq_7_bits_uop_lrs1 <= 6'h0;
      stq_7_bits_uop_lrs2 <= 6'h0;
      stq_7_bits_uop_lrs3 <= 6'h0;
      stq_7_bits_uop_dst_rtype <= 2'h2;
      stq_7_bits_uop_lrs1_rtype <= 2'h0;
      stq_7_bits_uop_lrs2_rtype <= 2'h0;
      stq_7_bits_uop_debug_fsrc <= 2'h0;
      stq_7_bits_uop_debug_tsrc <= 2'h0;
      stq_8_bits_uop_uopc <= 7'h0;
      stq_8_bits_uop_inst <= 32'h0;
      stq_8_bits_uop_debug_inst <= 32'h0;
      stq_8_bits_uop_debug_pc <= 40'h0;
      stq_8_bits_uop_iq_type <= 3'h0;
      stq_8_bits_uop_fu_code <= 10'h0;
      stq_8_bits_uop_ctrl_br_type <= 4'h0;
      stq_8_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_8_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_8_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_8_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_8_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_8_bits_uop_iw_state <= 2'h0;
      stq_8_bits_uop_br_mask <= 20'h0;
      stq_8_bits_uop_br_tag <= 5'h0;
      stq_8_bits_uop_ftq_idx <= 6'h0;
      stq_8_bits_uop_pc_lob <= 6'h0;
      stq_8_bits_uop_imm_packed <= 20'h0;
      stq_8_bits_uop_csr_addr <= 12'h0;
      stq_8_bits_uop_rob_idx <= 7'h0;
      stq_8_bits_uop_ldq_idx <= 5'h0;
      stq_8_bits_uop_stq_idx <= 5'h0;
      stq_8_bits_uop_rxq_idx <= 2'h0;
      stq_8_bits_uop_pdst <= 7'h0;
      stq_8_bits_uop_prs1 <= 7'h0;
      stq_8_bits_uop_prs2 <= 7'h0;
      stq_8_bits_uop_prs3 <= 7'h0;
      stq_8_bits_uop_ppred <= 6'h0;
      stq_8_bits_uop_stale_pdst <= 7'h0;
      stq_8_bits_uop_exc_cause <= 64'h0;
      stq_8_bits_uop_mem_cmd <= 5'h0;
      stq_8_bits_uop_mem_size <= 2'h0;
      stq_8_bits_uop_ldst <= 6'h0;
      stq_8_bits_uop_lrs1 <= 6'h0;
      stq_8_bits_uop_lrs2 <= 6'h0;
      stq_8_bits_uop_lrs3 <= 6'h0;
      stq_8_bits_uop_dst_rtype <= 2'h2;
      stq_8_bits_uop_lrs1_rtype <= 2'h0;
      stq_8_bits_uop_lrs2_rtype <= 2'h0;
      stq_8_bits_uop_debug_fsrc <= 2'h0;
      stq_8_bits_uop_debug_tsrc <= 2'h0;
      stq_9_bits_uop_uopc <= 7'h0;
      stq_9_bits_uop_inst <= 32'h0;
      stq_9_bits_uop_debug_inst <= 32'h0;
      stq_9_bits_uop_debug_pc <= 40'h0;
      stq_9_bits_uop_iq_type <= 3'h0;
      stq_9_bits_uop_fu_code <= 10'h0;
      stq_9_bits_uop_ctrl_br_type <= 4'h0;
      stq_9_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_9_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_9_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_9_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_9_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_9_bits_uop_iw_state <= 2'h0;
      stq_9_bits_uop_br_mask <= 20'h0;
      stq_9_bits_uop_br_tag <= 5'h0;
      stq_9_bits_uop_ftq_idx <= 6'h0;
      stq_9_bits_uop_pc_lob <= 6'h0;
      stq_9_bits_uop_imm_packed <= 20'h0;
      stq_9_bits_uop_csr_addr <= 12'h0;
      stq_9_bits_uop_rob_idx <= 7'h0;
      stq_9_bits_uop_ldq_idx <= 5'h0;
      stq_9_bits_uop_stq_idx <= 5'h0;
      stq_9_bits_uop_rxq_idx <= 2'h0;
      stq_9_bits_uop_pdst <= 7'h0;
      stq_9_bits_uop_prs1 <= 7'h0;
      stq_9_bits_uop_prs2 <= 7'h0;
      stq_9_bits_uop_prs3 <= 7'h0;
      stq_9_bits_uop_ppred <= 6'h0;
      stq_9_bits_uop_stale_pdst <= 7'h0;
      stq_9_bits_uop_exc_cause <= 64'h0;
      stq_9_bits_uop_mem_cmd <= 5'h0;
      stq_9_bits_uop_mem_size <= 2'h0;
      stq_9_bits_uop_ldst <= 6'h0;
      stq_9_bits_uop_lrs1 <= 6'h0;
      stq_9_bits_uop_lrs2 <= 6'h0;
      stq_9_bits_uop_lrs3 <= 6'h0;
      stq_9_bits_uop_dst_rtype <= 2'h2;
      stq_9_bits_uop_lrs1_rtype <= 2'h0;
      stq_9_bits_uop_lrs2_rtype <= 2'h0;
      stq_9_bits_uop_debug_fsrc <= 2'h0;
      stq_9_bits_uop_debug_tsrc <= 2'h0;
      stq_10_bits_uop_uopc <= 7'h0;
      stq_10_bits_uop_inst <= 32'h0;
      stq_10_bits_uop_debug_inst <= 32'h0;
      stq_10_bits_uop_debug_pc <= 40'h0;
      stq_10_bits_uop_iq_type <= 3'h0;
      stq_10_bits_uop_fu_code <= 10'h0;
      stq_10_bits_uop_ctrl_br_type <= 4'h0;
      stq_10_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_10_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_10_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_10_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_10_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_10_bits_uop_iw_state <= 2'h0;
      stq_10_bits_uop_br_mask <= 20'h0;
      stq_10_bits_uop_br_tag <= 5'h0;
      stq_10_bits_uop_ftq_idx <= 6'h0;
      stq_10_bits_uop_pc_lob <= 6'h0;
      stq_10_bits_uop_imm_packed <= 20'h0;
      stq_10_bits_uop_csr_addr <= 12'h0;
      stq_10_bits_uop_rob_idx <= 7'h0;
      stq_10_bits_uop_ldq_idx <= 5'h0;
      stq_10_bits_uop_stq_idx <= 5'h0;
      stq_10_bits_uop_rxq_idx <= 2'h0;
      stq_10_bits_uop_pdst <= 7'h0;
      stq_10_bits_uop_prs1 <= 7'h0;
      stq_10_bits_uop_prs2 <= 7'h0;
      stq_10_bits_uop_prs3 <= 7'h0;
      stq_10_bits_uop_ppred <= 6'h0;
      stq_10_bits_uop_stale_pdst <= 7'h0;
      stq_10_bits_uop_exc_cause <= 64'h0;
      stq_10_bits_uop_mem_cmd <= 5'h0;
      stq_10_bits_uop_mem_size <= 2'h0;
      stq_10_bits_uop_ldst <= 6'h0;
      stq_10_bits_uop_lrs1 <= 6'h0;
      stq_10_bits_uop_lrs2 <= 6'h0;
      stq_10_bits_uop_lrs3 <= 6'h0;
      stq_10_bits_uop_dst_rtype <= 2'h2;
      stq_10_bits_uop_lrs1_rtype <= 2'h0;
      stq_10_bits_uop_lrs2_rtype <= 2'h0;
      stq_10_bits_uop_debug_fsrc <= 2'h0;
      stq_10_bits_uop_debug_tsrc <= 2'h0;
      stq_11_bits_uop_uopc <= 7'h0;
      stq_11_bits_uop_inst <= 32'h0;
      stq_11_bits_uop_debug_inst <= 32'h0;
      stq_11_bits_uop_debug_pc <= 40'h0;
      stq_11_bits_uop_iq_type <= 3'h0;
      stq_11_bits_uop_fu_code <= 10'h0;
      stq_11_bits_uop_ctrl_br_type <= 4'h0;
      stq_11_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_11_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_11_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_11_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_11_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_11_bits_uop_iw_state <= 2'h0;
      stq_11_bits_uop_br_mask <= 20'h0;
      stq_11_bits_uop_br_tag <= 5'h0;
      stq_11_bits_uop_ftq_idx <= 6'h0;
      stq_11_bits_uop_pc_lob <= 6'h0;
      stq_11_bits_uop_imm_packed <= 20'h0;
      stq_11_bits_uop_csr_addr <= 12'h0;
      stq_11_bits_uop_rob_idx <= 7'h0;
      stq_11_bits_uop_ldq_idx <= 5'h0;
      stq_11_bits_uop_stq_idx <= 5'h0;
      stq_11_bits_uop_rxq_idx <= 2'h0;
      stq_11_bits_uop_pdst <= 7'h0;
      stq_11_bits_uop_prs1 <= 7'h0;
      stq_11_bits_uop_prs2 <= 7'h0;
      stq_11_bits_uop_prs3 <= 7'h0;
      stq_11_bits_uop_ppred <= 6'h0;
      stq_11_bits_uop_stale_pdst <= 7'h0;
      stq_11_bits_uop_exc_cause <= 64'h0;
      stq_11_bits_uop_mem_cmd <= 5'h0;
      stq_11_bits_uop_mem_size <= 2'h0;
      stq_11_bits_uop_ldst <= 6'h0;
      stq_11_bits_uop_lrs1 <= 6'h0;
      stq_11_bits_uop_lrs2 <= 6'h0;
      stq_11_bits_uop_lrs3 <= 6'h0;
      stq_11_bits_uop_dst_rtype <= 2'h2;
      stq_11_bits_uop_lrs1_rtype <= 2'h0;
      stq_11_bits_uop_lrs2_rtype <= 2'h0;
      stq_11_bits_uop_debug_fsrc <= 2'h0;
      stq_11_bits_uop_debug_tsrc <= 2'h0;
      stq_12_bits_uop_uopc <= 7'h0;
      stq_12_bits_uop_inst <= 32'h0;
      stq_12_bits_uop_debug_inst <= 32'h0;
      stq_12_bits_uop_debug_pc <= 40'h0;
      stq_12_bits_uop_iq_type <= 3'h0;
      stq_12_bits_uop_fu_code <= 10'h0;
      stq_12_bits_uop_ctrl_br_type <= 4'h0;
      stq_12_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_12_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_12_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_12_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_12_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_12_bits_uop_iw_state <= 2'h0;
      stq_12_bits_uop_br_mask <= 20'h0;
      stq_12_bits_uop_br_tag <= 5'h0;
      stq_12_bits_uop_ftq_idx <= 6'h0;
      stq_12_bits_uop_pc_lob <= 6'h0;
      stq_12_bits_uop_imm_packed <= 20'h0;
      stq_12_bits_uop_csr_addr <= 12'h0;
      stq_12_bits_uop_rob_idx <= 7'h0;
      stq_12_bits_uop_ldq_idx <= 5'h0;
      stq_12_bits_uop_stq_idx <= 5'h0;
      stq_12_bits_uop_rxq_idx <= 2'h0;
      stq_12_bits_uop_pdst <= 7'h0;
      stq_12_bits_uop_prs1 <= 7'h0;
      stq_12_bits_uop_prs2 <= 7'h0;
      stq_12_bits_uop_prs3 <= 7'h0;
      stq_12_bits_uop_ppred <= 6'h0;
      stq_12_bits_uop_stale_pdst <= 7'h0;
      stq_12_bits_uop_exc_cause <= 64'h0;
      stq_12_bits_uop_mem_cmd <= 5'h0;
      stq_12_bits_uop_mem_size <= 2'h0;
      stq_12_bits_uop_ldst <= 6'h0;
      stq_12_bits_uop_lrs1 <= 6'h0;
      stq_12_bits_uop_lrs2 <= 6'h0;
      stq_12_bits_uop_lrs3 <= 6'h0;
      stq_12_bits_uop_dst_rtype <= 2'h2;
      stq_12_bits_uop_lrs1_rtype <= 2'h0;
      stq_12_bits_uop_lrs2_rtype <= 2'h0;
      stq_12_bits_uop_debug_fsrc <= 2'h0;
      stq_12_bits_uop_debug_tsrc <= 2'h0;
      stq_13_bits_uop_uopc <= 7'h0;
      stq_13_bits_uop_inst <= 32'h0;
      stq_13_bits_uop_debug_inst <= 32'h0;
      stq_13_bits_uop_debug_pc <= 40'h0;
      stq_13_bits_uop_iq_type <= 3'h0;
      stq_13_bits_uop_fu_code <= 10'h0;
      stq_13_bits_uop_ctrl_br_type <= 4'h0;
      stq_13_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_13_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_13_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_13_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_13_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_13_bits_uop_iw_state <= 2'h0;
      stq_13_bits_uop_br_mask <= 20'h0;
      stq_13_bits_uop_br_tag <= 5'h0;
      stq_13_bits_uop_ftq_idx <= 6'h0;
      stq_13_bits_uop_pc_lob <= 6'h0;
      stq_13_bits_uop_imm_packed <= 20'h0;
      stq_13_bits_uop_csr_addr <= 12'h0;
      stq_13_bits_uop_rob_idx <= 7'h0;
      stq_13_bits_uop_ldq_idx <= 5'h0;
      stq_13_bits_uop_stq_idx <= 5'h0;
      stq_13_bits_uop_rxq_idx <= 2'h0;
      stq_13_bits_uop_pdst <= 7'h0;
      stq_13_bits_uop_prs1 <= 7'h0;
      stq_13_bits_uop_prs2 <= 7'h0;
      stq_13_bits_uop_prs3 <= 7'h0;
      stq_13_bits_uop_ppred <= 6'h0;
      stq_13_bits_uop_stale_pdst <= 7'h0;
      stq_13_bits_uop_exc_cause <= 64'h0;
      stq_13_bits_uop_mem_cmd <= 5'h0;
      stq_13_bits_uop_mem_size <= 2'h0;
      stq_13_bits_uop_ldst <= 6'h0;
      stq_13_bits_uop_lrs1 <= 6'h0;
      stq_13_bits_uop_lrs2 <= 6'h0;
      stq_13_bits_uop_lrs3 <= 6'h0;
      stq_13_bits_uop_dst_rtype <= 2'h2;
      stq_13_bits_uop_lrs1_rtype <= 2'h0;
      stq_13_bits_uop_lrs2_rtype <= 2'h0;
      stq_13_bits_uop_debug_fsrc <= 2'h0;
      stq_13_bits_uop_debug_tsrc <= 2'h0;
      stq_14_bits_uop_uopc <= 7'h0;
      stq_14_bits_uop_inst <= 32'h0;
      stq_14_bits_uop_debug_inst <= 32'h0;
      stq_14_bits_uop_debug_pc <= 40'h0;
      stq_14_bits_uop_iq_type <= 3'h0;
      stq_14_bits_uop_fu_code <= 10'h0;
      stq_14_bits_uop_ctrl_br_type <= 4'h0;
      stq_14_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_14_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_14_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_14_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_14_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_14_bits_uop_iw_state <= 2'h0;
      stq_14_bits_uop_br_mask <= 20'h0;
      stq_14_bits_uop_br_tag <= 5'h0;
      stq_14_bits_uop_ftq_idx <= 6'h0;
      stq_14_bits_uop_pc_lob <= 6'h0;
      stq_14_bits_uop_imm_packed <= 20'h0;
      stq_14_bits_uop_csr_addr <= 12'h0;
      stq_14_bits_uop_rob_idx <= 7'h0;
      stq_14_bits_uop_ldq_idx <= 5'h0;
      stq_14_bits_uop_stq_idx <= 5'h0;
      stq_14_bits_uop_rxq_idx <= 2'h0;
      stq_14_bits_uop_pdst <= 7'h0;
      stq_14_bits_uop_prs1 <= 7'h0;
      stq_14_bits_uop_prs2 <= 7'h0;
      stq_14_bits_uop_prs3 <= 7'h0;
      stq_14_bits_uop_ppred <= 6'h0;
      stq_14_bits_uop_stale_pdst <= 7'h0;
      stq_14_bits_uop_exc_cause <= 64'h0;
      stq_14_bits_uop_mem_cmd <= 5'h0;
      stq_14_bits_uop_mem_size <= 2'h0;
      stq_14_bits_uop_ldst <= 6'h0;
      stq_14_bits_uop_lrs1 <= 6'h0;
      stq_14_bits_uop_lrs2 <= 6'h0;
      stq_14_bits_uop_lrs3 <= 6'h0;
      stq_14_bits_uop_dst_rtype <= 2'h2;
      stq_14_bits_uop_lrs1_rtype <= 2'h0;
      stq_14_bits_uop_lrs2_rtype <= 2'h0;
      stq_14_bits_uop_debug_fsrc <= 2'h0;
      stq_14_bits_uop_debug_tsrc <= 2'h0;
      stq_15_bits_uop_uopc <= 7'h0;
      stq_15_bits_uop_inst <= 32'h0;
      stq_15_bits_uop_debug_inst <= 32'h0;
      stq_15_bits_uop_debug_pc <= 40'h0;
      stq_15_bits_uop_iq_type <= 3'h0;
      stq_15_bits_uop_fu_code <= 10'h0;
      stq_15_bits_uop_ctrl_br_type <= 4'h0;
      stq_15_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_15_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_15_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_15_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_15_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_15_bits_uop_iw_state <= 2'h0;
      stq_15_bits_uop_br_mask <= 20'h0;
      stq_15_bits_uop_br_tag <= 5'h0;
      stq_15_bits_uop_ftq_idx <= 6'h0;
      stq_15_bits_uop_pc_lob <= 6'h0;
      stq_15_bits_uop_imm_packed <= 20'h0;
      stq_15_bits_uop_csr_addr <= 12'h0;
      stq_15_bits_uop_rob_idx <= 7'h0;
      stq_15_bits_uop_ldq_idx <= 5'h0;
      stq_15_bits_uop_stq_idx <= 5'h0;
      stq_15_bits_uop_rxq_idx <= 2'h0;
      stq_15_bits_uop_pdst <= 7'h0;
      stq_15_bits_uop_prs1 <= 7'h0;
      stq_15_bits_uop_prs2 <= 7'h0;
      stq_15_bits_uop_prs3 <= 7'h0;
      stq_15_bits_uop_ppred <= 6'h0;
      stq_15_bits_uop_stale_pdst <= 7'h0;
      stq_15_bits_uop_exc_cause <= 64'h0;
      stq_15_bits_uop_mem_cmd <= 5'h0;
      stq_15_bits_uop_mem_size <= 2'h0;
      stq_15_bits_uop_ldst <= 6'h0;
      stq_15_bits_uop_lrs1 <= 6'h0;
      stq_15_bits_uop_lrs2 <= 6'h0;
      stq_15_bits_uop_lrs3 <= 6'h0;
      stq_15_bits_uop_dst_rtype <= 2'h2;
      stq_15_bits_uop_lrs1_rtype <= 2'h0;
      stq_15_bits_uop_lrs2_rtype <= 2'h0;
      stq_15_bits_uop_debug_fsrc <= 2'h0;
      stq_15_bits_uop_debug_tsrc <= 2'h0;
      stq_16_bits_uop_uopc <= 7'h0;
      stq_16_bits_uop_inst <= 32'h0;
      stq_16_bits_uop_debug_inst <= 32'h0;
      stq_16_bits_uop_debug_pc <= 40'h0;
      stq_16_bits_uop_iq_type <= 3'h0;
      stq_16_bits_uop_fu_code <= 10'h0;
      stq_16_bits_uop_ctrl_br_type <= 4'h0;
      stq_16_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_16_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_16_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_16_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_16_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_16_bits_uop_iw_state <= 2'h0;
      stq_16_bits_uop_br_mask <= 20'h0;
      stq_16_bits_uop_br_tag <= 5'h0;
      stq_16_bits_uop_ftq_idx <= 6'h0;
      stq_16_bits_uop_pc_lob <= 6'h0;
      stq_16_bits_uop_imm_packed <= 20'h0;
      stq_16_bits_uop_csr_addr <= 12'h0;
      stq_16_bits_uop_rob_idx <= 7'h0;
      stq_16_bits_uop_ldq_idx <= 5'h0;
      stq_16_bits_uop_stq_idx <= 5'h0;
      stq_16_bits_uop_rxq_idx <= 2'h0;
      stq_16_bits_uop_pdst <= 7'h0;
      stq_16_bits_uop_prs1 <= 7'h0;
      stq_16_bits_uop_prs2 <= 7'h0;
      stq_16_bits_uop_prs3 <= 7'h0;
      stq_16_bits_uop_ppred <= 6'h0;
      stq_16_bits_uop_stale_pdst <= 7'h0;
      stq_16_bits_uop_exc_cause <= 64'h0;
      stq_16_bits_uop_mem_cmd <= 5'h0;
      stq_16_bits_uop_mem_size <= 2'h0;
      stq_16_bits_uop_ldst <= 6'h0;
      stq_16_bits_uop_lrs1 <= 6'h0;
      stq_16_bits_uop_lrs2 <= 6'h0;
      stq_16_bits_uop_lrs3 <= 6'h0;
      stq_16_bits_uop_dst_rtype <= 2'h2;
      stq_16_bits_uop_lrs1_rtype <= 2'h0;
      stq_16_bits_uop_lrs2_rtype <= 2'h0;
      stq_16_bits_uop_debug_fsrc <= 2'h0;
      stq_16_bits_uop_debug_tsrc <= 2'h0;
      stq_17_bits_uop_uopc <= 7'h0;
      stq_17_bits_uop_inst <= 32'h0;
      stq_17_bits_uop_debug_inst <= 32'h0;
      stq_17_bits_uop_debug_pc <= 40'h0;
      stq_17_bits_uop_iq_type <= 3'h0;
      stq_17_bits_uop_fu_code <= 10'h0;
      stq_17_bits_uop_ctrl_br_type <= 4'h0;
      stq_17_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_17_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_17_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_17_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_17_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_17_bits_uop_iw_state <= 2'h0;
      stq_17_bits_uop_br_mask <= 20'h0;
      stq_17_bits_uop_br_tag <= 5'h0;
      stq_17_bits_uop_ftq_idx <= 6'h0;
      stq_17_bits_uop_pc_lob <= 6'h0;
      stq_17_bits_uop_imm_packed <= 20'h0;
      stq_17_bits_uop_csr_addr <= 12'h0;
      stq_17_bits_uop_rob_idx <= 7'h0;
      stq_17_bits_uop_ldq_idx <= 5'h0;
      stq_17_bits_uop_stq_idx <= 5'h0;
      stq_17_bits_uop_rxq_idx <= 2'h0;
      stq_17_bits_uop_pdst <= 7'h0;
      stq_17_bits_uop_prs1 <= 7'h0;
      stq_17_bits_uop_prs2 <= 7'h0;
      stq_17_bits_uop_prs3 <= 7'h0;
      stq_17_bits_uop_ppred <= 6'h0;
      stq_17_bits_uop_stale_pdst <= 7'h0;
      stq_17_bits_uop_exc_cause <= 64'h0;
      stq_17_bits_uop_mem_cmd <= 5'h0;
      stq_17_bits_uop_mem_size <= 2'h0;
      stq_17_bits_uop_ldst <= 6'h0;
      stq_17_bits_uop_lrs1 <= 6'h0;
      stq_17_bits_uop_lrs2 <= 6'h0;
      stq_17_bits_uop_lrs3 <= 6'h0;
      stq_17_bits_uop_dst_rtype <= 2'h2;
      stq_17_bits_uop_lrs1_rtype <= 2'h0;
      stq_17_bits_uop_lrs2_rtype <= 2'h0;
      stq_17_bits_uop_debug_fsrc <= 2'h0;
      stq_17_bits_uop_debug_tsrc <= 2'h0;
      stq_18_bits_uop_uopc <= 7'h0;
      stq_18_bits_uop_inst <= 32'h0;
      stq_18_bits_uop_debug_inst <= 32'h0;
      stq_18_bits_uop_debug_pc <= 40'h0;
      stq_18_bits_uop_iq_type <= 3'h0;
      stq_18_bits_uop_fu_code <= 10'h0;
      stq_18_bits_uop_ctrl_br_type <= 4'h0;
      stq_18_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_18_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_18_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_18_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_18_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_18_bits_uop_iw_state <= 2'h0;
      stq_18_bits_uop_br_mask <= 20'h0;
      stq_18_bits_uop_br_tag <= 5'h0;
      stq_18_bits_uop_ftq_idx <= 6'h0;
      stq_18_bits_uop_pc_lob <= 6'h0;
      stq_18_bits_uop_imm_packed <= 20'h0;
      stq_18_bits_uop_csr_addr <= 12'h0;
      stq_18_bits_uop_rob_idx <= 7'h0;
      stq_18_bits_uop_ldq_idx <= 5'h0;
      stq_18_bits_uop_stq_idx <= 5'h0;
      stq_18_bits_uop_rxq_idx <= 2'h0;
      stq_18_bits_uop_pdst <= 7'h0;
      stq_18_bits_uop_prs1 <= 7'h0;
      stq_18_bits_uop_prs2 <= 7'h0;
      stq_18_bits_uop_prs3 <= 7'h0;
      stq_18_bits_uop_ppred <= 6'h0;
      stq_18_bits_uop_stale_pdst <= 7'h0;
      stq_18_bits_uop_exc_cause <= 64'h0;
      stq_18_bits_uop_mem_cmd <= 5'h0;
      stq_18_bits_uop_mem_size <= 2'h0;
      stq_18_bits_uop_ldst <= 6'h0;
      stq_18_bits_uop_lrs1 <= 6'h0;
      stq_18_bits_uop_lrs2 <= 6'h0;
      stq_18_bits_uop_lrs3 <= 6'h0;
      stq_18_bits_uop_dst_rtype <= 2'h2;
      stq_18_bits_uop_lrs1_rtype <= 2'h0;
      stq_18_bits_uop_lrs2_rtype <= 2'h0;
      stq_18_bits_uop_debug_fsrc <= 2'h0;
      stq_18_bits_uop_debug_tsrc <= 2'h0;
      stq_19_bits_uop_uopc <= 7'h0;
      stq_19_bits_uop_inst <= 32'h0;
      stq_19_bits_uop_debug_inst <= 32'h0;
      stq_19_bits_uop_debug_pc <= 40'h0;
      stq_19_bits_uop_iq_type <= 3'h0;
      stq_19_bits_uop_fu_code <= 10'h0;
      stq_19_bits_uop_ctrl_br_type <= 4'h0;
      stq_19_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_19_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_19_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_19_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_19_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_19_bits_uop_iw_state <= 2'h0;
      stq_19_bits_uop_br_mask <= 20'h0;
      stq_19_bits_uop_br_tag <= 5'h0;
      stq_19_bits_uop_ftq_idx <= 6'h0;
      stq_19_bits_uop_pc_lob <= 6'h0;
      stq_19_bits_uop_imm_packed <= 20'h0;
      stq_19_bits_uop_csr_addr <= 12'h0;
      stq_19_bits_uop_rob_idx <= 7'h0;
      stq_19_bits_uop_ldq_idx <= 5'h0;
      stq_19_bits_uop_stq_idx <= 5'h0;
      stq_19_bits_uop_rxq_idx <= 2'h0;
      stq_19_bits_uop_pdst <= 7'h0;
      stq_19_bits_uop_prs1 <= 7'h0;
      stq_19_bits_uop_prs2 <= 7'h0;
      stq_19_bits_uop_prs3 <= 7'h0;
      stq_19_bits_uop_ppred <= 6'h0;
      stq_19_bits_uop_stale_pdst <= 7'h0;
      stq_19_bits_uop_exc_cause <= 64'h0;
      stq_19_bits_uop_mem_cmd <= 5'h0;
      stq_19_bits_uop_mem_size <= 2'h0;
      stq_19_bits_uop_ldst <= 6'h0;
      stq_19_bits_uop_lrs1 <= 6'h0;
      stq_19_bits_uop_lrs2 <= 6'h0;
      stq_19_bits_uop_lrs3 <= 6'h0;
      stq_19_bits_uop_dst_rtype <= 2'h2;
      stq_19_bits_uop_lrs1_rtype <= 2'h0;
      stq_19_bits_uop_lrs2_rtype <= 2'h0;
      stq_19_bits_uop_debug_fsrc <= 2'h0;
      stq_19_bits_uop_debug_tsrc <= 2'h0;
      stq_20_bits_uop_uopc <= 7'h0;
      stq_20_bits_uop_inst <= 32'h0;
      stq_20_bits_uop_debug_inst <= 32'h0;
      stq_20_bits_uop_debug_pc <= 40'h0;
      stq_20_bits_uop_iq_type <= 3'h0;
      stq_20_bits_uop_fu_code <= 10'h0;
      stq_20_bits_uop_ctrl_br_type <= 4'h0;
      stq_20_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_20_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_20_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_20_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_20_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_20_bits_uop_iw_state <= 2'h0;
      stq_20_bits_uop_br_mask <= 20'h0;
      stq_20_bits_uop_br_tag <= 5'h0;
      stq_20_bits_uop_ftq_idx <= 6'h0;
      stq_20_bits_uop_pc_lob <= 6'h0;
      stq_20_bits_uop_imm_packed <= 20'h0;
      stq_20_bits_uop_csr_addr <= 12'h0;
      stq_20_bits_uop_rob_idx <= 7'h0;
      stq_20_bits_uop_ldq_idx <= 5'h0;
      stq_20_bits_uop_stq_idx <= 5'h0;
      stq_20_bits_uop_rxq_idx <= 2'h0;
      stq_20_bits_uop_pdst <= 7'h0;
      stq_20_bits_uop_prs1 <= 7'h0;
      stq_20_bits_uop_prs2 <= 7'h0;
      stq_20_bits_uop_prs3 <= 7'h0;
      stq_20_bits_uop_ppred <= 6'h0;
      stq_20_bits_uop_stale_pdst <= 7'h0;
      stq_20_bits_uop_exc_cause <= 64'h0;
      stq_20_bits_uop_mem_cmd <= 5'h0;
      stq_20_bits_uop_mem_size <= 2'h0;
      stq_20_bits_uop_ldst <= 6'h0;
      stq_20_bits_uop_lrs1 <= 6'h0;
      stq_20_bits_uop_lrs2 <= 6'h0;
      stq_20_bits_uop_lrs3 <= 6'h0;
      stq_20_bits_uop_dst_rtype <= 2'h2;
      stq_20_bits_uop_lrs1_rtype <= 2'h0;
      stq_20_bits_uop_lrs2_rtype <= 2'h0;
      stq_20_bits_uop_debug_fsrc <= 2'h0;
      stq_20_bits_uop_debug_tsrc <= 2'h0;
      stq_21_bits_uop_uopc <= 7'h0;
      stq_21_bits_uop_inst <= 32'h0;
      stq_21_bits_uop_debug_inst <= 32'h0;
      stq_21_bits_uop_debug_pc <= 40'h0;
      stq_21_bits_uop_iq_type <= 3'h0;
      stq_21_bits_uop_fu_code <= 10'h0;
      stq_21_bits_uop_ctrl_br_type <= 4'h0;
      stq_21_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_21_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_21_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_21_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_21_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_21_bits_uop_iw_state <= 2'h0;
      stq_21_bits_uop_br_mask <= 20'h0;
      stq_21_bits_uop_br_tag <= 5'h0;
      stq_21_bits_uop_ftq_idx <= 6'h0;
      stq_21_bits_uop_pc_lob <= 6'h0;
      stq_21_bits_uop_imm_packed <= 20'h0;
      stq_21_bits_uop_csr_addr <= 12'h0;
      stq_21_bits_uop_rob_idx <= 7'h0;
      stq_21_bits_uop_ldq_idx <= 5'h0;
      stq_21_bits_uop_stq_idx <= 5'h0;
      stq_21_bits_uop_rxq_idx <= 2'h0;
      stq_21_bits_uop_pdst <= 7'h0;
      stq_21_bits_uop_prs1 <= 7'h0;
      stq_21_bits_uop_prs2 <= 7'h0;
      stq_21_bits_uop_prs3 <= 7'h0;
      stq_21_bits_uop_ppred <= 6'h0;
      stq_21_bits_uop_stale_pdst <= 7'h0;
      stq_21_bits_uop_exc_cause <= 64'h0;
      stq_21_bits_uop_mem_cmd <= 5'h0;
      stq_21_bits_uop_mem_size <= 2'h0;
      stq_21_bits_uop_ldst <= 6'h0;
      stq_21_bits_uop_lrs1 <= 6'h0;
      stq_21_bits_uop_lrs2 <= 6'h0;
      stq_21_bits_uop_lrs3 <= 6'h0;
      stq_21_bits_uop_dst_rtype <= 2'h2;
      stq_21_bits_uop_lrs1_rtype <= 2'h0;
      stq_21_bits_uop_lrs2_rtype <= 2'h0;
      stq_21_bits_uop_debug_fsrc <= 2'h0;
      stq_21_bits_uop_debug_tsrc <= 2'h0;
      stq_22_bits_uop_uopc <= 7'h0;
      stq_22_bits_uop_inst <= 32'h0;
      stq_22_bits_uop_debug_inst <= 32'h0;
      stq_22_bits_uop_debug_pc <= 40'h0;
      stq_22_bits_uop_iq_type <= 3'h0;
      stq_22_bits_uop_fu_code <= 10'h0;
      stq_22_bits_uop_ctrl_br_type <= 4'h0;
      stq_22_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_22_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_22_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_22_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_22_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_22_bits_uop_iw_state <= 2'h0;
      stq_22_bits_uop_br_mask <= 20'h0;
      stq_22_bits_uop_br_tag <= 5'h0;
      stq_22_bits_uop_ftq_idx <= 6'h0;
      stq_22_bits_uop_pc_lob <= 6'h0;
      stq_22_bits_uop_imm_packed <= 20'h0;
      stq_22_bits_uop_csr_addr <= 12'h0;
      stq_22_bits_uop_rob_idx <= 7'h0;
      stq_22_bits_uop_ldq_idx <= 5'h0;
      stq_22_bits_uop_stq_idx <= 5'h0;
      stq_22_bits_uop_rxq_idx <= 2'h0;
      stq_22_bits_uop_pdst <= 7'h0;
      stq_22_bits_uop_prs1 <= 7'h0;
      stq_22_bits_uop_prs2 <= 7'h0;
      stq_22_bits_uop_prs3 <= 7'h0;
      stq_22_bits_uop_ppred <= 6'h0;
      stq_22_bits_uop_stale_pdst <= 7'h0;
      stq_22_bits_uop_exc_cause <= 64'h0;
      stq_22_bits_uop_mem_cmd <= 5'h0;
      stq_22_bits_uop_mem_size <= 2'h0;
      stq_22_bits_uop_ldst <= 6'h0;
      stq_22_bits_uop_lrs1 <= 6'h0;
      stq_22_bits_uop_lrs2 <= 6'h0;
      stq_22_bits_uop_lrs3 <= 6'h0;
      stq_22_bits_uop_dst_rtype <= 2'h2;
      stq_22_bits_uop_lrs1_rtype <= 2'h0;
      stq_22_bits_uop_lrs2_rtype <= 2'h0;
      stq_22_bits_uop_debug_fsrc <= 2'h0;
      stq_22_bits_uop_debug_tsrc <= 2'h0;
      stq_23_bits_uop_uopc <= 7'h0;
      stq_23_bits_uop_inst <= 32'h0;
      stq_23_bits_uop_debug_inst <= 32'h0;
      stq_23_bits_uop_debug_pc <= 40'h0;
      stq_23_bits_uop_iq_type <= 3'h0;
      stq_23_bits_uop_fu_code <= 10'h0;
      stq_23_bits_uop_ctrl_br_type <= 4'h0;
      stq_23_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_23_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_23_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_23_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_23_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_23_bits_uop_iw_state <= 2'h0;
      stq_23_bits_uop_br_mask <= 20'h0;
      stq_23_bits_uop_br_tag <= 5'h0;
      stq_23_bits_uop_ftq_idx <= 6'h0;
      stq_23_bits_uop_pc_lob <= 6'h0;
      stq_23_bits_uop_imm_packed <= 20'h0;
      stq_23_bits_uop_csr_addr <= 12'h0;
      stq_23_bits_uop_rob_idx <= 7'h0;
      stq_23_bits_uop_ldq_idx <= 5'h0;
      stq_23_bits_uop_stq_idx <= 5'h0;
      stq_23_bits_uop_rxq_idx <= 2'h0;
      stq_23_bits_uop_pdst <= 7'h0;
      stq_23_bits_uop_prs1 <= 7'h0;
      stq_23_bits_uop_prs2 <= 7'h0;
      stq_23_bits_uop_prs3 <= 7'h0;
      stq_23_bits_uop_ppred <= 6'h0;
      stq_23_bits_uop_stale_pdst <= 7'h0;
      stq_23_bits_uop_exc_cause <= 64'h0;
      stq_23_bits_uop_mem_cmd <= 5'h0;
      stq_23_bits_uop_mem_size <= 2'h0;
      stq_23_bits_uop_ldst <= 6'h0;
      stq_23_bits_uop_lrs1 <= 6'h0;
      stq_23_bits_uop_lrs2 <= 6'h0;
      stq_23_bits_uop_lrs3 <= 6'h0;
      stq_23_bits_uop_dst_rtype <= 2'h2;
      stq_23_bits_uop_lrs1_rtype <= 2'h0;
      stq_23_bits_uop_lrs2_rtype <= 2'h0;
      stq_23_bits_uop_debug_fsrc <= 2'h0;
      stq_23_bits_uop_debug_tsrc <= 2'h0;
      stq_24_bits_uop_uopc <= 7'h0;
      stq_24_bits_uop_inst <= 32'h0;
      stq_24_bits_uop_debug_inst <= 32'h0;
      stq_24_bits_uop_debug_pc <= 40'h0;
      stq_24_bits_uop_iq_type <= 3'h0;
      stq_24_bits_uop_fu_code <= 10'h0;
      stq_24_bits_uop_ctrl_br_type <= 4'h0;
      stq_24_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_24_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_24_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_24_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_24_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_24_bits_uop_iw_state <= 2'h0;
      stq_24_bits_uop_br_mask <= 20'h0;
      stq_24_bits_uop_br_tag <= 5'h0;
      stq_24_bits_uop_ftq_idx <= 6'h0;
      stq_24_bits_uop_pc_lob <= 6'h0;
      stq_24_bits_uop_imm_packed <= 20'h0;
      stq_24_bits_uop_csr_addr <= 12'h0;
      stq_24_bits_uop_rob_idx <= 7'h0;
      stq_24_bits_uop_ldq_idx <= 5'h0;
      stq_24_bits_uop_stq_idx <= 5'h0;
      stq_24_bits_uop_rxq_idx <= 2'h0;
      stq_24_bits_uop_pdst <= 7'h0;
      stq_24_bits_uop_prs1 <= 7'h0;
      stq_24_bits_uop_prs2 <= 7'h0;
      stq_24_bits_uop_prs3 <= 7'h0;
      stq_24_bits_uop_ppred <= 6'h0;
      stq_24_bits_uop_stale_pdst <= 7'h0;
      stq_24_bits_uop_exc_cause <= 64'h0;
      stq_24_bits_uop_mem_cmd <= 5'h0;
      stq_24_bits_uop_mem_size <= 2'h0;
      stq_24_bits_uop_ldst <= 6'h0;
      stq_24_bits_uop_lrs1 <= 6'h0;
      stq_24_bits_uop_lrs2 <= 6'h0;
      stq_24_bits_uop_lrs3 <= 6'h0;
      stq_24_bits_uop_dst_rtype <= 2'h2;
      stq_24_bits_uop_lrs1_rtype <= 2'h0;
      stq_24_bits_uop_lrs2_rtype <= 2'h0;
      stq_24_bits_uop_debug_fsrc <= 2'h0;
      stq_24_bits_uop_debug_tsrc <= 2'h0;
      stq_25_bits_uop_uopc <= 7'h0;
      stq_25_bits_uop_inst <= 32'h0;
      stq_25_bits_uop_debug_inst <= 32'h0;
      stq_25_bits_uop_debug_pc <= 40'h0;
      stq_25_bits_uop_iq_type <= 3'h0;
      stq_25_bits_uop_fu_code <= 10'h0;
      stq_25_bits_uop_ctrl_br_type <= 4'h0;
      stq_25_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_25_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_25_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_25_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_25_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_25_bits_uop_iw_state <= 2'h0;
      stq_25_bits_uop_br_mask <= 20'h0;
      stq_25_bits_uop_br_tag <= 5'h0;
      stq_25_bits_uop_ftq_idx <= 6'h0;
      stq_25_bits_uop_pc_lob <= 6'h0;
      stq_25_bits_uop_imm_packed <= 20'h0;
      stq_25_bits_uop_csr_addr <= 12'h0;
      stq_25_bits_uop_rob_idx <= 7'h0;
      stq_25_bits_uop_ldq_idx <= 5'h0;
      stq_25_bits_uop_stq_idx <= 5'h0;
      stq_25_bits_uop_rxq_idx <= 2'h0;
      stq_25_bits_uop_pdst <= 7'h0;
      stq_25_bits_uop_prs1 <= 7'h0;
      stq_25_bits_uop_prs2 <= 7'h0;
      stq_25_bits_uop_prs3 <= 7'h0;
      stq_25_bits_uop_ppred <= 6'h0;
      stq_25_bits_uop_stale_pdst <= 7'h0;
      stq_25_bits_uop_exc_cause <= 64'h0;
      stq_25_bits_uop_mem_cmd <= 5'h0;
      stq_25_bits_uop_mem_size <= 2'h0;
      stq_25_bits_uop_ldst <= 6'h0;
      stq_25_bits_uop_lrs1 <= 6'h0;
      stq_25_bits_uop_lrs2 <= 6'h0;
      stq_25_bits_uop_lrs3 <= 6'h0;
      stq_25_bits_uop_dst_rtype <= 2'h2;
      stq_25_bits_uop_lrs1_rtype <= 2'h0;
      stq_25_bits_uop_lrs2_rtype <= 2'h0;
      stq_25_bits_uop_debug_fsrc <= 2'h0;
      stq_25_bits_uop_debug_tsrc <= 2'h0;
      stq_26_bits_uop_uopc <= 7'h0;
      stq_26_bits_uop_inst <= 32'h0;
      stq_26_bits_uop_debug_inst <= 32'h0;
      stq_26_bits_uop_debug_pc <= 40'h0;
      stq_26_bits_uop_iq_type <= 3'h0;
      stq_26_bits_uop_fu_code <= 10'h0;
      stq_26_bits_uop_ctrl_br_type <= 4'h0;
      stq_26_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_26_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_26_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_26_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_26_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_26_bits_uop_iw_state <= 2'h0;
      stq_26_bits_uop_br_mask <= 20'h0;
      stq_26_bits_uop_br_tag <= 5'h0;
      stq_26_bits_uop_ftq_idx <= 6'h0;
      stq_26_bits_uop_pc_lob <= 6'h0;
      stq_26_bits_uop_imm_packed <= 20'h0;
      stq_26_bits_uop_csr_addr <= 12'h0;
      stq_26_bits_uop_rob_idx <= 7'h0;
      stq_26_bits_uop_ldq_idx <= 5'h0;
      stq_26_bits_uop_stq_idx <= 5'h0;
      stq_26_bits_uop_rxq_idx <= 2'h0;
      stq_26_bits_uop_pdst <= 7'h0;
      stq_26_bits_uop_prs1 <= 7'h0;
      stq_26_bits_uop_prs2 <= 7'h0;
      stq_26_bits_uop_prs3 <= 7'h0;
      stq_26_bits_uop_ppred <= 6'h0;
      stq_26_bits_uop_stale_pdst <= 7'h0;
      stq_26_bits_uop_exc_cause <= 64'h0;
      stq_26_bits_uop_mem_cmd <= 5'h0;
      stq_26_bits_uop_mem_size <= 2'h0;
      stq_26_bits_uop_ldst <= 6'h0;
      stq_26_bits_uop_lrs1 <= 6'h0;
      stq_26_bits_uop_lrs2 <= 6'h0;
      stq_26_bits_uop_lrs3 <= 6'h0;
      stq_26_bits_uop_dst_rtype <= 2'h2;
      stq_26_bits_uop_lrs1_rtype <= 2'h0;
      stq_26_bits_uop_lrs2_rtype <= 2'h0;
      stq_26_bits_uop_debug_fsrc <= 2'h0;
      stq_26_bits_uop_debug_tsrc <= 2'h0;
      stq_27_bits_uop_uopc <= 7'h0;
      stq_27_bits_uop_inst <= 32'h0;
      stq_27_bits_uop_debug_inst <= 32'h0;
      stq_27_bits_uop_debug_pc <= 40'h0;
      stq_27_bits_uop_iq_type <= 3'h0;
      stq_27_bits_uop_fu_code <= 10'h0;
      stq_27_bits_uop_ctrl_br_type <= 4'h0;
      stq_27_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_27_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_27_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_27_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_27_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_27_bits_uop_iw_state <= 2'h0;
      stq_27_bits_uop_br_mask <= 20'h0;
      stq_27_bits_uop_br_tag <= 5'h0;
      stq_27_bits_uop_ftq_idx <= 6'h0;
      stq_27_bits_uop_pc_lob <= 6'h0;
      stq_27_bits_uop_imm_packed <= 20'h0;
      stq_27_bits_uop_csr_addr <= 12'h0;
      stq_27_bits_uop_rob_idx <= 7'h0;
      stq_27_bits_uop_ldq_idx <= 5'h0;
      stq_27_bits_uop_stq_idx <= 5'h0;
      stq_27_bits_uop_rxq_idx <= 2'h0;
      stq_27_bits_uop_pdst <= 7'h0;
      stq_27_bits_uop_prs1 <= 7'h0;
      stq_27_bits_uop_prs2 <= 7'h0;
      stq_27_bits_uop_prs3 <= 7'h0;
      stq_27_bits_uop_ppred <= 6'h0;
      stq_27_bits_uop_stale_pdst <= 7'h0;
      stq_27_bits_uop_exc_cause <= 64'h0;
      stq_27_bits_uop_mem_cmd <= 5'h0;
      stq_27_bits_uop_mem_size <= 2'h0;
      stq_27_bits_uop_ldst <= 6'h0;
      stq_27_bits_uop_lrs1 <= 6'h0;
      stq_27_bits_uop_lrs2 <= 6'h0;
      stq_27_bits_uop_lrs3 <= 6'h0;
      stq_27_bits_uop_dst_rtype <= 2'h2;
      stq_27_bits_uop_lrs1_rtype <= 2'h0;
      stq_27_bits_uop_lrs2_rtype <= 2'h0;
      stq_27_bits_uop_debug_fsrc <= 2'h0;
      stq_27_bits_uop_debug_tsrc <= 2'h0;
      stq_28_bits_uop_uopc <= 7'h0;
      stq_28_bits_uop_inst <= 32'h0;
      stq_28_bits_uop_debug_inst <= 32'h0;
      stq_28_bits_uop_debug_pc <= 40'h0;
      stq_28_bits_uop_iq_type <= 3'h0;
      stq_28_bits_uop_fu_code <= 10'h0;
      stq_28_bits_uop_ctrl_br_type <= 4'h0;
      stq_28_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_28_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_28_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_28_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_28_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_28_bits_uop_iw_state <= 2'h0;
      stq_28_bits_uop_br_mask <= 20'h0;
      stq_28_bits_uop_br_tag <= 5'h0;
      stq_28_bits_uop_ftq_idx <= 6'h0;
      stq_28_bits_uop_pc_lob <= 6'h0;
      stq_28_bits_uop_imm_packed <= 20'h0;
      stq_28_bits_uop_csr_addr <= 12'h0;
      stq_28_bits_uop_rob_idx <= 7'h0;
      stq_28_bits_uop_ldq_idx <= 5'h0;
      stq_28_bits_uop_stq_idx <= 5'h0;
      stq_28_bits_uop_rxq_idx <= 2'h0;
      stq_28_bits_uop_pdst <= 7'h0;
      stq_28_bits_uop_prs1 <= 7'h0;
      stq_28_bits_uop_prs2 <= 7'h0;
      stq_28_bits_uop_prs3 <= 7'h0;
      stq_28_bits_uop_ppred <= 6'h0;
      stq_28_bits_uop_stale_pdst <= 7'h0;
      stq_28_bits_uop_exc_cause <= 64'h0;
      stq_28_bits_uop_mem_cmd <= 5'h0;
      stq_28_bits_uop_mem_size <= 2'h0;
      stq_28_bits_uop_ldst <= 6'h0;
      stq_28_bits_uop_lrs1 <= 6'h0;
      stq_28_bits_uop_lrs2 <= 6'h0;
      stq_28_bits_uop_lrs3 <= 6'h0;
      stq_28_bits_uop_dst_rtype <= 2'h2;
      stq_28_bits_uop_lrs1_rtype <= 2'h0;
      stq_28_bits_uop_lrs2_rtype <= 2'h0;
      stq_28_bits_uop_debug_fsrc <= 2'h0;
      stq_28_bits_uop_debug_tsrc <= 2'h0;
      stq_29_bits_uop_uopc <= 7'h0;
      stq_29_bits_uop_inst <= 32'h0;
      stq_29_bits_uop_debug_inst <= 32'h0;
      stq_29_bits_uop_debug_pc <= 40'h0;
      stq_29_bits_uop_iq_type <= 3'h0;
      stq_29_bits_uop_fu_code <= 10'h0;
      stq_29_bits_uop_ctrl_br_type <= 4'h0;
      stq_29_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_29_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_29_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_29_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_29_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_29_bits_uop_iw_state <= 2'h0;
      stq_29_bits_uop_br_mask <= 20'h0;
      stq_29_bits_uop_br_tag <= 5'h0;
      stq_29_bits_uop_ftq_idx <= 6'h0;
      stq_29_bits_uop_pc_lob <= 6'h0;
      stq_29_bits_uop_imm_packed <= 20'h0;
      stq_29_bits_uop_csr_addr <= 12'h0;
      stq_29_bits_uop_rob_idx <= 7'h0;
      stq_29_bits_uop_ldq_idx <= 5'h0;
      stq_29_bits_uop_stq_idx <= 5'h0;
      stq_29_bits_uop_rxq_idx <= 2'h0;
      stq_29_bits_uop_pdst <= 7'h0;
      stq_29_bits_uop_prs1 <= 7'h0;
      stq_29_bits_uop_prs2 <= 7'h0;
      stq_29_bits_uop_prs3 <= 7'h0;
      stq_29_bits_uop_ppred <= 6'h0;
      stq_29_bits_uop_stale_pdst <= 7'h0;
      stq_29_bits_uop_exc_cause <= 64'h0;
      stq_29_bits_uop_mem_cmd <= 5'h0;
      stq_29_bits_uop_mem_size <= 2'h0;
      stq_29_bits_uop_ldst <= 6'h0;
      stq_29_bits_uop_lrs1 <= 6'h0;
      stq_29_bits_uop_lrs2 <= 6'h0;
      stq_29_bits_uop_lrs3 <= 6'h0;
      stq_29_bits_uop_dst_rtype <= 2'h2;
      stq_29_bits_uop_lrs1_rtype <= 2'h0;
      stq_29_bits_uop_lrs2_rtype <= 2'h0;
      stq_29_bits_uop_debug_fsrc <= 2'h0;
      stq_29_bits_uop_debug_tsrc <= 2'h0;
      stq_30_bits_uop_uopc <= 7'h0;
      stq_30_bits_uop_inst <= 32'h0;
      stq_30_bits_uop_debug_inst <= 32'h0;
      stq_30_bits_uop_debug_pc <= 40'h0;
      stq_30_bits_uop_iq_type <= 3'h0;
      stq_30_bits_uop_fu_code <= 10'h0;
      stq_30_bits_uop_ctrl_br_type <= 4'h0;
      stq_30_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_30_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_30_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_30_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_30_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_30_bits_uop_iw_state <= 2'h0;
      stq_30_bits_uop_br_mask <= 20'h0;
      stq_30_bits_uop_br_tag <= 5'h0;
      stq_30_bits_uop_ftq_idx <= 6'h0;
      stq_30_bits_uop_pc_lob <= 6'h0;
      stq_30_bits_uop_imm_packed <= 20'h0;
      stq_30_bits_uop_csr_addr <= 12'h0;
      stq_30_bits_uop_rob_idx <= 7'h0;
      stq_30_bits_uop_ldq_idx <= 5'h0;
      stq_30_bits_uop_stq_idx <= 5'h0;
      stq_30_bits_uop_rxq_idx <= 2'h0;
      stq_30_bits_uop_pdst <= 7'h0;
      stq_30_bits_uop_prs1 <= 7'h0;
      stq_30_bits_uop_prs2 <= 7'h0;
      stq_30_bits_uop_prs3 <= 7'h0;
      stq_30_bits_uop_ppred <= 6'h0;
      stq_30_bits_uop_stale_pdst <= 7'h0;
      stq_30_bits_uop_exc_cause <= 64'h0;
      stq_30_bits_uop_mem_cmd <= 5'h0;
      stq_30_bits_uop_mem_size <= 2'h0;
      stq_30_bits_uop_ldst <= 6'h0;
      stq_30_bits_uop_lrs1 <= 6'h0;
      stq_30_bits_uop_lrs2 <= 6'h0;
      stq_30_bits_uop_lrs3 <= 6'h0;
      stq_30_bits_uop_dst_rtype <= 2'h2;
      stq_30_bits_uop_lrs1_rtype <= 2'h0;
      stq_30_bits_uop_lrs2_rtype <= 2'h0;
      stq_30_bits_uop_debug_fsrc <= 2'h0;
      stq_30_bits_uop_debug_tsrc <= 2'h0;
      stq_31_bits_uop_uopc <= 7'h0;
      stq_31_bits_uop_inst <= 32'h0;
      stq_31_bits_uop_debug_inst <= 32'h0;
      stq_31_bits_uop_debug_pc <= 40'h0;
      stq_31_bits_uop_iq_type <= 3'h0;
      stq_31_bits_uop_fu_code <= 10'h0;
      stq_31_bits_uop_ctrl_br_type <= 4'h0;
      stq_31_bits_uop_ctrl_op1_sel <= 2'h0;
      stq_31_bits_uop_ctrl_op2_sel <= 3'h0;
      stq_31_bits_uop_ctrl_imm_sel <= 3'h0;
      stq_31_bits_uop_ctrl_op_fcn <= 4'h0;
      stq_31_bits_uop_ctrl_csr_cmd <= 3'h0;
      stq_31_bits_uop_iw_state <= 2'h0;
      stq_31_bits_uop_br_mask <= 20'h0;
      stq_31_bits_uop_br_tag <= 5'h0;
      stq_31_bits_uop_ftq_idx <= 6'h0;
      stq_31_bits_uop_pc_lob <= 6'h0;
      stq_31_bits_uop_imm_packed <= 20'h0;
      stq_31_bits_uop_csr_addr <= 12'h0;
      stq_31_bits_uop_rob_idx <= 7'h0;
      stq_31_bits_uop_ldq_idx <= 5'h0;
      stq_31_bits_uop_stq_idx <= 5'h0;
      stq_31_bits_uop_rxq_idx <= 2'h0;
      stq_31_bits_uop_pdst <= 7'h0;
      stq_31_bits_uop_prs1 <= 7'h0;
      stq_31_bits_uop_prs2 <= 7'h0;
      stq_31_bits_uop_prs3 <= 7'h0;
      stq_31_bits_uop_ppred <= 6'h0;
      stq_31_bits_uop_stale_pdst <= 7'h0;
      stq_31_bits_uop_exc_cause <= 64'h0;
      stq_31_bits_uop_mem_cmd <= 5'h0;
      stq_31_bits_uop_mem_size <= 2'h0;
      stq_31_bits_uop_ldst <= 6'h0;
      stq_31_bits_uop_lrs1 <= 6'h0;
      stq_31_bits_uop_lrs2 <= 6'h0;
      stq_31_bits_uop_lrs3 <= 6'h0;
      stq_31_bits_uop_dst_rtype <= 2'h2;
      stq_31_bits_uop_lrs1_rtype <= 2'h0;
      stq_31_bits_uop_lrs2_rtype <= 2'h0;
      stq_31_bits_uop_debug_fsrc <= 2'h0;
      stq_31_bits_uop_debug_tsrc <= 2'h0;
      stq_head <= 5'h0;
      stq_commit_head <= 5'h0;
      stq_execute_head <= 5'h0;
    end
    else begin
      if (_GEN_2454) begin
        if (_GEN_2134) begin
          if (_GEN_2037) begin
            if (_GEN_1653) begin
            end
            else begin
              stq_0_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_0_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_0_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_0_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_0_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_0_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_0_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_0_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_0_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_0_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_0_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_0_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_0_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_0_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_0_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_0_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_0_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_0_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_0_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_0_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_0_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_0_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_0_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_0_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_0_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_0_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_0_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_0_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_0_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_0_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_0_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_0_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_0_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_0_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_0_valid)
        stq_0_bits_uop_br_mask <= stq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2454) begin
        if (_GEN_2134) begin
          if (_GEN_2037) begin
            if (_GEN_1653) begin
            end
            else
              stq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_0_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_0_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2454) begin
        if (_GEN_2134) begin
          if (_GEN_2037) begin
            if (_GEN_1653) begin
            end
            else begin
              stq_0_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_0_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_0_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_0_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_0_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_0_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_0_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_0_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_0_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_0_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_0_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_0_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_0_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_0_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_0_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_0_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_0_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_0_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_0_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_0_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_0_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_0_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_0_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_0_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_0_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_0_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_0_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_0_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_0_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_0_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2805) begin
        if (_exe_tlb_uop_T_9)
          stq_0_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_0_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_0_bits_uop_pdst <= casez_tmp_246;
        else
          stq_0_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2678) begin
        if (_exe_tlb_uop_T_2)
          stq_0_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_0_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_0_bits_uop_pdst <= casez_tmp_246;
        else
          stq_0_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2454) begin
        if (_GEN_2134) begin
          if (_GEN_2037) begin
            if (_GEN_1653) begin
            end
            else
              stq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_0_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_0_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2454) begin
        if (_GEN_2134) begin
          if (_GEN_2037) begin
            if (_GEN_1653) begin
            end
            else begin
              stq_0_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_0_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_0_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
            end
          end
          else begin
            stq_0_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_0_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_0_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
          end
        end
        else begin
          stq_0_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_0_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_0_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
        end
      end
      else begin
        stq_0_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_0_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_0_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
      end
      if (dis_ld_val_3) begin
        if (_GEN_2134) begin
          if (dis_ld_val_1) begin
            if (_GEN_1653) begin
            end
            else
              stq_0_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5815)
            stq_0_bits_uop_ppred <= 6'h0;
        end
        else
          stq_0_bits_uop_ppred <= 6'h0;
        if (_GEN_2135) begin
          if (dis_ld_val_1) begin
            if (_GEN_1654) begin
            end
            else
              stq_1_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5816)
            stq_1_bits_uop_ppred <= 6'h0;
        end
        else
          stq_1_bits_uop_ppred <= 6'h0;
        if (_GEN_2136) begin
          if (dis_ld_val_1) begin
            if (_GEN_1655) begin
            end
            else
              stq_2_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5817)
            stq_2_bits_uop_ppred <= 6'h0;
        end
        else
          stq_2_bits_uop_ppred <= 6'h0;
        if (_GEN_2137) begin
          if (dis_ld_val_1) begin
            if (_GEN_1656) begin
            end
            else
              stq_3_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5818)
            stq_3_bits_uop_ppred <= 6'h0;
        end
        else
          stq_3_bits_uop_ppred <= 6'h0;
        if (_GEN_2138) begin
          if (dis_ld_val_1) begin
            if (_GEN_1657) begin
            end
            else
              stq_4_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5819)
            stq_4_bits_uop_ppred <= 6'h0;
        end
        else
          stq_4_bits_uop_ppred <= 6'h0;
        if (_GEN_2139) begin
          if (dis_ld_val_1) begin
            if (_GEN_1658) begin
            end
            else
              stq_5_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5820)
            stq_5_bits_uop_ppred <= 6'h0;
        end
        else
          stq_5_bits_uop_ppred <= 6'h0;
        if (_GEN_2140) begin
          if (dis_ld_val_1) begin
            if (_GEN_1659) begin
            end
            else
              stq_6_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5821)
            stq_6_bits_uop_ppred <= 6'h0;
        end
        else
          stq_6_bits_uop_ppred <= 6'h0;
        if (_GEN_2141) begin
          if (dis_ld_val_1) begin
            if (_GEN_1660) begin
            end
            else
              stq_7_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5822)
            stq_7_bits_uop_ppred <= 6'h0;
        end
        else
          stq_7_bits_uop_ppred <= 6'h0;
        if (_GEN_2142) begin
          if (dis_ld_val_1) begin
            if (_GEN_1661) begin
            end
            else
              stq_8_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5823)
            stq_8_bits_uop_ppred <= 6'h0;
        end
        else
          stq_8_bits_uop_ppred <= 6'h0;
        if (_GEN_2143) begin
          if (dis_ld_val_1) begin
            if (_GEN_1662) begin
            end
            else
              stq_9_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5824)
            stq_9_bits_uop_ppred <= 6'h0;
        end
        else
          stq_9_bits_uop_ppred <= 6'h0;
        if (_GEN_2144) begin
          if (dis_ld_val_1) begin
            if (_GEN_1663) begin
            end
            else
              stq_10_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5825)
            stq_10_bits_uop_ppred <= 6'h0;
        end
        else
          stq_10_bits_uop_ppred <= 6'h0;
        if (_GEN_2145) begin
          if (dis_ld_val_1) begin
            if (_GEN_1664) begin
            end
            else
              stq_11_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5826)
            stq_11_bits_uop_ppred <= 6'h0;
        end
        else
          stq_11_bits_uop_ppred <= 6'h0;
        if (_GEN_2146) begin
          if (dis_ld_val_1) begin
            if (_GEN_1665) begin
            end
            else
              stq_12_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5827)
            stq_12_bits_uop_ppred <= 6'h0;
        end
        else
          stq_12_bits_uop_ppred <= 6'h0;
        if (_GEN_2147) begin
          if (dis_ld_val_1) begin
            if (_GEN_1666) begin
            end
            else
              stq_13_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5828)
            stq_13_bits_uop_ppred <= 6'h0;
        end
        else
          stq_13_bits_uop_ppred <= 6'h0;
        if (_GEN_2148) begin
          if (dis_ld_val_1) begin
            if (_GEN_1667) begin
            end
            else
              stq_14_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5829)
            stq_14_bits_uop_ppred <= 6'h0;
        end
        else
          stq_14_bits_uop_ppred <= 6'h0;
        if (_GEN_2149) begin
          if (dis_ld_val_1) begin
            if (_GEN_1668) begin
            end
            else
              stq_15_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5830)
            stq_15_bits_uop_ppred <= 6'h0;
        end
        else
          stq_15_bits_uop_ppred <= 6'h0;
        if (_GEN_2150) begin
          if (dis_ld_val_1) begin
            if (_GEN_1669) begin
            end
            else
              stq_16_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5831)
            stq_16_bits_uop_ppred <= 6'h0;
        end
        else
          stq_16_bits_uop_ppred <= 6'h0;
        if (_GEN_2151) begin
          if (dis_ld_val_1) begin
            if (_GEN_1670) begin
            end
            else
              stq_17_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5832)
            stq_17_bits_uop_ppred <= 6'h0;
        end
        else
          stq_17_bits_uop_ppred <= 6'h0;
        if (_GEN_2152) begin
          if (dis_ld_val_1) begin
            if (_GEN_1671) begin
            end
            else
              stq_18_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5833)
            stq_18_bits_uop_ppred <= 6'h0;
        end
        else
          stq_18_bits_uop_ppred <= 6'h0;
        if (_GEN_2153) begin
          if (dis_ld_val_1) begin
            if (_GEN_1672) begin
            end
            else
              stq_19_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5834)
            stq_19_bits_uop_ppred <= 6'h0;
        end
        else
          stq_19_bits_uop_ppred <= 6'h0;
        if (_GEN_2154) begin
          if (dis_ld_val_1) begin
            if (_GEN_1673) begin
            end
            else
              stq_20_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5835)
            stq_20_bits_uop_ppred <= 6'h0;
        end
        else
          stq_20_bits_uop_ppred <= 6'h0;
        if (_GEN_2155) begin
          if (dis_ld_val_1) begin
            if (_GEN_1674) begin
            end
            else
              stq_21_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5836)
            stq_21_bits_uop_ppred <= 6'h0;
        end
        else
          stq_21_bits_uop_ppred <= 6'h0;
        if (_GEN_2156) begin
          if (dis_ld_val_1) begin
            if (_GEN_1675) begin
            end
            else
              stq_22_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5837)
            stq_22_bits_uop_ppred <= 6'h0;
        end
        else
          stq_22_bits_uop_ppred <= 6'h0;
        if (_GEN_2157) begin
          if (dis_ld_val_1) begin
            if (_GEN_1676) begin
            end
            else
              stq_23_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5838)
            stq_23_bits_uop_ppred <= 6'h0;
        end
        else
          stq_23_bits_uop_ppred <= 6'h0;
        if (_GEN_2158) begin
          if (dis_ld_val_1) begin
            if (_GEN_1677) begin
            end
            else
              stq_24_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5839)
            stq_24_bits_uop_ppred <= 6'h0;
        end
        else
          stq_24_bits_uop_ppred <= 6'h0;
        if (_GEN_2159) begin
          if (dis_ld_val_1) begin
            if (_GEN_1678) begin
            end
            else
              stq_25_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5840)
            stq_25_bits_uop_ppred <= 6'h0;
        end
        else
          stq_25_bits_uop_ppred <= 6'h0;
        if (_GEN_2160) begin
          if (dis_ld_val_1) begin
            if (_GEN_1679) begin
            end
            else
              stq_26_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5841)
            stq_26_bits_uop_ppred <= 6'h0;
        end
        else
          stq_26_bits_uop_ppred <= 6'h0;
        if (_GEN_2161) begin
          if (dis_ld_val_1) begin
            if (_GEN_1680) begin
            end
            else
              stq_27_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5842)
            stq_27_bits_uop_ppred <= 6'h0;
        end
        else
          stq_27_bits_uop_ppred <= 6'h0;
        if (_GEN_2162) begin
          if (dis_ld_val_1) begin
            if (_GEN_1681) begin
            end
            else
              stq_28_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5843)
            stq_28_bits_uop_ppred <= 6'h0;
        end
        else
          stq_28_bits_uop_ppred <= 6'h0;
        if (_GEN_2163) begin
          if (dis_ld_val_1) begin
            if (_GEN_1682) begin
            end
            else
              stq_29_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5844)
            stq_29_bits_uop_ppred <= 6'h0;
        end
        else
          stq_29_bits_uop_ppred <= 6'h0;
        if (_GEN_2164) begin
          if (dis_ld_val_1) begin
            if (_GEN_1683) begin
            end
            else
              stq_30_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5845)
            stq_30_bits_uop_ppred <= 6'h0;
        end
        else
          stq_30_bits_uop_ppred <= 6'h0;
        if (_GEN_2165) begin
          if (dis_ld_val_1) begin
            if (_GEN_1684) begin
            end
            else
              stq_31_bits_uop_ppred <= 6'h0;
          end
          else if (_GEN_5846)
            stq_31_bits_uop_ppred <= 6'h0;
        end
        else
          stq_31_bits_uop_ppred <= 6'h0;
      end
      else begin
        if (_GEN_2390 | ~_GEN_2134)
          stq_0_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1653) begin
          end
          else
            stq_0_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5815)
          stq_0_bits_uop_ppred <= 6'h0;
        if (_GEN_2392 | ~_GEN_2135)
          stq_1_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1654) begin
          end
          else
            stq_1_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5816)
          stq_1_bits_uop_ppred <= 6'h0;
        if (_GEN_2394 | ~_GEN_2136)
          stq_2_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1655) begin
          end
          else
            stq_2_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5817)
          stq_2_bits_uop_ppred <= 6'h0;
        if (_GEN_2396 | ~_GEN_2137)
          stq_3_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1656) begin
          end
          else
            stq_3_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5818)
          stq_3_bits_uop_ppred <= 6'h0;
        if (_GEN_2398 | ~_GEN_2138)
          stq_4_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1657) begin
          end
          else
            stq_4_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5819)
          stq_4_bits_uop_ppred <= 6'h0;
        if (_GEN_2400 | ~_GEN_2139)
          stq_5_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1658) begin
          end
          else
            stq_5_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5820)
          stq_5_bits_uop_ppred <= 6'h0;
        if (_GEN_2402 | ~_GEN_2140)
          stq_6_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1659) begin
          end
          else
            stq_6_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5821)
          stq_6_bits_uop_ppred <= 6'h0;
        if (_GEN_2404 | ~_GEN_2141)
          stq_7_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1660) begin
          end
          else
            stq_7_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5822)
          stq_7_bits_uop_ppred <= 6'h0;
        if (_GEN_2406 | ~_GEN_2142)
          stq_8_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1661) begin
          end
          else
            stq_8_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5823)
          stq_8_bits_uop_ppred <= 6'h0;
        if (_GEN_2408 | ~_GEN_2143)
          stq_9_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1662) begin
          end
          else
            stq_9_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5824)
          stq_9_bits_uop_ppred <= 6'h0;
        if (_GEN_2410 | ~_GEN_2144)
          stq_10_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1663) begin
          end
          else
            stq_10_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5825)
          stq_10_bits_uop_ppred <= 6'h0;
        if (_GEN_2412 | ~_GEN_2145)
          stq_11_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1664) begin
          end
          else
            stq_11_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5826)
          stq_11_bits_uop_ppred <= 6'h0;
        if (_GEN_2414 | ~_GEN_2146)
          stq_12_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1665) begin
          end
          else
            stq_12_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5827)
          stq_12_bits_uop_ppred <= 6'h0;
        if (_GEN_2416 | ~_GEN_2147)
          stq_13_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1666) begin
          end
          else
            stq_13_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5828)
          stq_13_bits_uop_ppred <= 6'h0;
        if (_GEN_2418 | ~_GEN_2148)
          stq_14_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1667) begin
          end
          else
            stq_14_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5829)
          stq_14_bits_uop_ppred <= 6'h0;
        if (_GEN_2420 | ~_GEN_2149)
          stq_15_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1668) begin
          end
          else
            stq_15_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5830)
          stq_15_bits_uop_ppred <= 6'h0;
        if (_GEN_2422 | ~_GEN_2150)
          stq_16_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1669) begin
          end
          else
            stq_16_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5831)
          stq_16_bits_uop_ppred <= 6'h0;
        if (_GEN_2424 | ~_GEN_2151)
          stq_17_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1670) begin
          end
          else
            stq_17_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5832)
          stq_17_bits_uop_ppred <= 6'h0;
        if (_GEN_2426 | ~_GEN_2152)
          stq_18_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1671) begin
          end
          else
            stq_18_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5833)
          stq_18_bits_uop_ppred <= 6'h0;
        if (_GEN_2428 | ~_GEN_2153)
          stq_19_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1672) begin
          end
          else
            stq_19_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5834)
          stq_19_bits_uop_ppred <= 6'h0;
        if (_GEN_2430 | ~_GEN_2154)
          stq_20_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1673) begin
          end
          else
            stq_20_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5835)
          stq_20_bits_uop_ppred <= 6'h0;
        if (_GEN_2432 | ~_GEN_2155)
          stq_21_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1674) begin
          end
          else
            stq_21_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5836)
          stq_21_bits_uop_ppred <= 6'h0;
        if (_GEN_2434 | ~_GEN_2156)
          stq_22_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1675) begin
          end
          else
            stq_22_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5837)
          stq_22_bits_uop_ppred <= 6'h0;
        if (_GEN_2436 | ~_GEN_2157)
          stq_23_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1676) begin
          end
          else
            stq_23_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5838)
          stq_23_bits_uop_ppred <= 6'h0;
        if (_GEN_2438 | ~_GEN_2158)
          stq_24_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1677) begin
          end
          else
            stq_24_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5839)
          stq_24_bits_uop_ppred <= 6'h0;
        if (_GEN_2440 | ~_GEN_2159)
          stq_25_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1678) begin
          end
          else
            stq_25_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5840)
          stq_25_bits_uop_ppred <= 6'h0;
        if (_GEN_2442 | ~_GEN_2160)
          stq_26_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1679) begin
          end
          else
            stq_26_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5841)
          stq_26_bits_uop_ppred <= 6'h0;
        if (_GEN_2444 | ~_GEN_2161)
          stq_27_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1680) begin
          end
          else
            stq_27_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5842)
          stq_27_bits_uop_ppred <= 6'h0;
        if (_GEN_2446 | ~_GEN_2162)
          stq_28_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1681) begin
          end
          else
            stq_28_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5843)
          stq_28_bits_uop_ppred <= 6'h0;
        if (_GEN_2448 | ~_GEN_2163)
          stq_29_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1682) begin
          end
          else
            stq_29_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5844)
          stq_29_bits_uop_ppred <= 6'h0;
        if (_GEN_2450 | ~_GEN_2164)
          stq_30_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1683) begin
          end
          else
            stq_30_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5845)
          stq_30_bits_uop_ppred <= 6'h0;
        if (_GEN_2452 | ~_GEN_2165)
          stq_31_bits_uop_ppred <= 6'h0;
        else if (dis_ld_val_1) begin
          if (_GEN_1684) begin
          end
          else
            stq_31_bits_uop_ppred <= 6'h0;
        end
        else if (_GEN_5846)
          stq_31_bits_uop_ppred <= 6'h0;
      end
      if (_GEN_2454) begin
        if (_GEN_2134) begin
          if (_GEN_2037) begin
            if (_GEN_1653) begin
            end
            else begin
              stq_0_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_0_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_0_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_0_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_0_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_0_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_0_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_0_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_0_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_0_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_0_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_0_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_0_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_0_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_0_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_0_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_0_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_0_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_0_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_0_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_0_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_0_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_0_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_0_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_0_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_0_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_0_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_0_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_0_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_0_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_0_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_0_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_0_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_0_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2455) begin
        if (_GEN_2135) begin
          if (_GEN_2038) begin
            if (_GEN_1654) begin
            end
            else begin
              stq_1_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_1_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_1_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_1_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_1_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_1_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_1_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_1_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_1_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_1_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_1_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_1_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_1_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_1_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_1_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_1_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_1_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_1_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_1_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_1_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_1_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_1_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_1_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_1_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_1_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_1_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_1_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_1_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_1_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_1_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_1_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_1_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_1_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_1_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_1_valid)
        stq_1_bits_uop_br_mask <= stq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2455) begin
        if (_GEN_2135) begin
          if (_GEN_2038) begin
            if (_GEN_1654) begin
            end
            else
              stq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_1_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_1_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2455) begin
        if (_GEN_2135) begin
          if (_GEN_2038) begin
            if (_GEN_1654) begin
            end
            else begin
              stq_1_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_1_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_1_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_1_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_1_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_1_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_1_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_1_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_1_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_1_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_1_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_1_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_1_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_1_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_1_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_1_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_1_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_1_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_1_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_1_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_1_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_1_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_1_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_1_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_1_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_1_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_1_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_1_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_1_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_1_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2807) begin
        if (_exe_tlb_uop_T_9)
          stq_1_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_1_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_1_bits_uop_pdst <= casez_tmp_246;
        else
          stq_1_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2679) begin
        if (_exe_tlb_uop_T_2)
          stq_1_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_1_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_1_bits_uop_pdst <= casez_tmp_246;
        else
          stq_1_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2455) begin
        if (_GEN_2135) begin
          if (_GEN_2038) begin
            if (_GEN_1654) begin
            end
            else
              stq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_1_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_1_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2455) begin
        if (_GEN_2135) begin
          if (_GEN_2038) begin
            if (_GEN_1654) begin
            end
            else begin
              stq_1_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_1_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_1_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_1_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_1_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_1_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_1_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_1_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_1_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_1_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_1_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_1_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_1_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_1_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_1_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_1_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_1_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_1_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_1_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_1_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_1_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_1_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_1_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_1_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_1_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_1_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_1_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_1_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_1_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_1_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_1_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_1_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_1_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_1_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_1_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_1_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_1_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_1_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_1_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_1_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_1_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_1_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_1_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_1_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_1_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_1_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2456) begin
        if (_GEN_2136) begin
          if (_GEN_2039) begin
            if (_GEN_1655) begin
            end
            else begin
              stq_2_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_2_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_2_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_2_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_2_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_2_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_2_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_2_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_2_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_2_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_2_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_2_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_2_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_2_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_2_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_2_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_2_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_2_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_2_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_2_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_2_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_2_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_2_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_2_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_2_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_2_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_2_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_2_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_2_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_2_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_2_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_2_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_2_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_2_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_2_valid)
        stq_2_bits_uop_br_mask <= stq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2456) begin
        if (_GEN_2136) begin
          if (_GEN_2039) begin
            if (_GEN_1655) begin
            end
            else
              stq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_2_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_2_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2456) begin
        if (_GEN_2136) begin
          if (_GEN_2039) begin
            if (_GEN_1655) begin
            end
            else begin
              stq_2_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_2_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_2_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_2_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_2_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_2_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_2_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_2_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_2_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_2_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_2_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_2_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_2_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_2_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_2_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_2_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_2_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_2_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_2_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_2_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_2_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_2_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_2_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_2_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_2_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_2_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_2_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_2_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_2_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_2_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2809) begin
        if (_exe_tlb_uop_T_9)
          stq_2_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_2_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_2_bits_uop_pdst <= casez_tmp_246;
        else
          stq_2_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2680) begin
        if (_exe_tlb_uop_T_2)
          stq_2_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_2_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_2_bits_uop_pdst <= casez_tmp_246;
        else
          stq_2_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2456) begin
        if (_GEN_2136) begin
          if (_GEN_2039) begin
            if (_GEN_1655) begin
            end
            else
              stq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_2_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_2_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2456) begin
        if (_GEN_2136) begin
          if (_GEN_2039) begin
            if (_GEN_1655) begin
            end
            else begin
              stq_2_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_2_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_2_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_2_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_2_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_2_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_2_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_2_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_2_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_2_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_2_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_2_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_2_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_2_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_2_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_2_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_2_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_2_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_2_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_2_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_2_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_2_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_2_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_2_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_2_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_2_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_2_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_2_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_2_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_2_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_2_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_2_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_2_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_2_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_2_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_2_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_2_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_2_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_2_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_2_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_2_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_2_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_2_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_2_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_2_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_2_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2457) begin
        if (_GEN_2137) begin
          if (_GEN_2040) begin
            if (_GEN_1656) begin
            end
            else begin
              stq_3_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_3_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_3_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_3_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_3_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_3_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_3_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_3_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_3_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_3_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_3_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_3_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_3_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_3_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_3_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_3_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_3_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_3_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_3_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_3_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_3_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_3_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_3_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_3_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_3_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_3_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_3_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_3_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_3_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_3_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_3_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_3_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_3_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_3_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_3_valid)
        stq_3_bits_uop_br_mask <= stq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2457) begin
        if (_GEN_2137) begin
          if (_GEN_2040) begin
            if (_GEN_1656) begin
            end
            else
              stq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_3_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_3_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2457) begin
        if (_GEN_2137) begin
          if (_GEN_2040) begin
            if (_GEN_1656) begin
            end
            else begin
              stq_3_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_3_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_3_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_3_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_3_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_3_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_3_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_3_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_3_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_3_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_3_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_3_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_3_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_3_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_3_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_3_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_3_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_3_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_3_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_3_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_3_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_3_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_3_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_3_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_3_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_3_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_3_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_3_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_3_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_3_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2811) begin
        if (_exe_tlb_uop_T_9)
          stq_3_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_3_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_3_bits_uop_pdst <= casez_tmp_246;
        else
          stq_3_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2681) begin
        if (_exe_tlb_uop_T_2)
          stq_3_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_3_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_3_bits_uop_pdst <= casez_tmp_246;
        else
          stq_3_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2457) begin
        if (_GEN_2137) begin
          if (_GEN_2040) begin
            if (_GEN_1656) begin
            end
            else
              stq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_3_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_3_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2457) begin
        if (_GEN_2137) begin
          if (_GEN_2040) begin
            if (_GEN_1656) begin
            end
            else begin
              stq_3_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_3_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_3_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_3_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_3_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_3_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_3_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_3_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_3_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_3_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_3_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_3_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_3_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_3_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_3_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_3_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_3_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_3_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_3_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_3_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_3_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_3_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_3_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_3_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_3_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_3_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_3_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_3_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_3_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_3_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_3_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_3_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_3_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_3_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_3_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_3_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_3_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_3_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_3_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_3_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_3_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_3_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_3_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_3_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_3_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_3_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2458) begin
        if (_GEN_2138) begin
          if (_GEN_2041) begin
            if (_GEN_1657) begin
            end
            else begin
              stq_4_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_4_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_4_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_4_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_4_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_4_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_4_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_4_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_4_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_4_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_4_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_4_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_4_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_4_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_4_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_4_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_4_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_4_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_4_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_4_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_4_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_4_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_4_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_4_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_4_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_4_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_4_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_4_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_4_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_4_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_4_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_4_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_4_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_4_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_4_valid)
        stq_4_bits_uop_br_mask <= stq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2458) begin
        if (_GEN_2138) begin
          if (_GEN_2041) begin
            if (_GEN_1657) begin
            end
            else
              stq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_4_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_4_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2458) begin
        if (_GEN_2138) begin
          if (_GEN_2041) begin
            if (_GEN_1657) begin
            end
            else begin
              stq_4_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_4_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_4_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_4_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_4_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_4_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_4_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_4_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_4_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_4_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_4_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_4_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_4_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_4_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_4_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_4_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_4_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_4_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_4_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_4_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_4_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_4_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_4_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_4_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_4_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_4_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_4_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_4_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_4_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_4_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2813) begin
        if (_exe_tlb_uop_T_9)
          stq_4_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_4_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_4_bits_uop_pdst <= casez_tmp_246;
        else
          stq_4_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2682) begin
        if (_exe_tlb_uop_T_2)
          stq_4_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_4_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_4_bits_uop_pdst <= casez_tmp_246;
        else
          stq_4_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2458) begin
        if (_GEN_2138) begin
          if (_GEN_2041) begin
            if (_GEN_1657) begin
            end
            else
              stq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_4_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_4_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2458) begin
        if (_GEN_2138) begin
          if (_GEN_2041) begin
            if (_GEN_1657) begin
            end
            else begin
              stq_4_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_4_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_4_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_4_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_4_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_4_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_4_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_4_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_4_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_4_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_4_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_4_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_4_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_4_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_4_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_4_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_4_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_4_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_4_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_4_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_4_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_4_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_4_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_4_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_4_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_4_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_4_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_4_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_4_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_4_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_4_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_4_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_4_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_4_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_4_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_4_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_4_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_4_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_4_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_4_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_4_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_4_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_4_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_4_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_4_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_4_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2459) begin
        if (_GEN_2139) begin
          if (_GEN_2042) begin
            if (_GEN_1658) begin
            end
            else begin
              stq_5_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_5_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_5_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_5_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_5_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_5_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_5_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_5_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_5_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_5_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_5_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_5_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_5_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_5_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_5_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_5_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_5_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_5_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_5_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_5_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_5_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_5_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_5_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_5_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_5_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_5_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_5_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_5_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_5_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_5_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_5_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_5_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_5_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_5_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_5_valid)
        stq_5_bits_uop_br_mask <= stq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2459) begin
        if (_GEN_2139) begin
          if (_GEN_2042) begin
            if (_GEN_1658) begin
            end
            else
              stq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_5_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_5_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2459) begin
        if (_GEN_2139) begin
          if (_GEN_2042) begin
            if (_GEN_1658) begin
            end
            else begin
              stq_5_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_5_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_5_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_5_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_5_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_5_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_5_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_5_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_5_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_5_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_5_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_5_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_5_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_5_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_5_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_5_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_5_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_5_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_5_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_5_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_5_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_5_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_5_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_5_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_5_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_5_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_5_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_5_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_5_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_5_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2815) begin
        if (_exe_tlb_uop_T_9)
          stq_5_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_5_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_5_bits_uop_pdst <= casez_tmp_246;
        else
          stq_5_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2683) begin
        if (_exe_tlb_uop_T_2)
          stq_5_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_5_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_5_bits_uop_pdst <= casez_tmp_246;
        else
          stq_5_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2459) begin
        if (_GEN_2139) begin
          if (_GEN_2042) begin
            if (_GEN_1658) begin
            end
            else
              stq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_5_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_5_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2459) begin
        if (_GEN_2139) begin
          if (_GEN_2042) begin
            if (_GEN_1658) begin
            end
            else begin
              stq_5_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_5_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_5_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_5_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_5_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_5_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_5_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_5_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_5_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_5_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_5_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_5_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_5_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_5_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_5_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_5_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_5_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_5_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_5_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_5_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_5_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_5_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_5_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_5_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_5_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_5_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_5_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_5_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_5_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_5_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_5_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_5_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_5_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_5_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_5_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_5_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_5_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_5_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_5_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_5_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_5_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_5_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_5_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_5_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_5_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_5_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2460) begin
        if (_GEN_2140) begin
          if (_GEN_2043) begin
            if (_GEN_1659) begin
            end
            else begin
              stq_6_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_6_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_6_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_6_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_6_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_6_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_6_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_6_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_6_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_6_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_6_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_6_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_6_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_6_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_6_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_6_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_6_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_6_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_6_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_6_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_6_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_6_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_6_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_6_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_6_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_6_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_6_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_6_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_6_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_6_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_6_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_6_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_6_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_6_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_6_valid)
        stq_6_bits_uop_br_mask <= stq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2460) begin
        if (_GEN_2140) begin
          if (_GEN_2043) begin
            if (_GEN_1659) begin
            end
            else
              stq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_6_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_6_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2460) begin
        if (_GEN_2140) begin
          if (_GEN_2043) begin
            if (_GEN_1659) begin
            end
            else begin
              stq_6_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_6_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_6_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_6_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_6_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_6_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_6_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_6_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_6_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_6_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_6_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_6_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_6_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_6_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_6_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_6_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_6_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_6_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_6_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_6_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_6_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_6_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_6_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_6_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_6_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_6_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_6_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_6_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_6_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_6_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2817) begin
        if (_exe_tlb_uop_T_9)
          stq_6_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_6_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_6_bits_uop_pdst <= casez_tmp_246;
        else
          stq_6_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2684) begin
        if (_exe_tlb_uop_T_2)
          stq_6_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_6_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_6_bits_uop_pdst <= casez_tmp_246;
        else
          stq_6_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2460) begin
        if (_GEN_2140) begin
          if (_GEN_2043) begin
            if (_GEN_1659) begin
            end
            else
              stq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_6_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_6_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2460) begin
        if (_GEN_2140) begin
          if (_GEN_2043) begin
            if (_GEN_1659) begin
            end
            else begin
              stq_6_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_6_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_6_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_6_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_6_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_6_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_6_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_6_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_6_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_6_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_6_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_6_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_6_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_6_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_6_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_6_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_6_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_6_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_6_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_6_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_6_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_6_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_6_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_6_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_6_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_6_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_6_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_6_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_6_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_6_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_6_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_6_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_6_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_6_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_6_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_6_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_6_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_6_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_6_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_6_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_6_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_6_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_6_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_6_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_6_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_6_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2461) begin
        if (_GEN_2141) begin
          if (_GEN_2044) begin
            if (_GEN_1660) begin
            end
            else begin
              stq_7_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_7_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_7_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_7_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_7_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_7_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_7_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_7_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_7_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_7_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_7_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_7_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_7_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_7_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_7_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_7_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_7_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_7_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_7_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_7_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_7_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_7_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_7_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_7_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_7_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_7_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_7_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_7_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_7_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_7_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_7_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_7_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_7_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_7_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_7_valid)
        stq_7_bits_uop_br_mask <= stq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2461) begin
        if (_GEN_2141) begin
          if (_GEN_2044) begin
            if (_GEN_1660) begin
            end
            else
              stq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_7_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_7_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2461) begin
        if (_GEN_2141) begin
          if (_GEN_2044) begin
            if (_GEN_1660) begin
            end
            else begin
              stq_7_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_7_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_7_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_7_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_7_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_7_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_7_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_7_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_7_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_7_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_7_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_7_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_7_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_7_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_7_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_7_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_7_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_7_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_7_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_7_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_7_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_7_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_7_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_7_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_7_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_7_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_7_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_7_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_7_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_7_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2819) begin
        if (_exe_tlb_uop_T_9)
          stq_7_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_7_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_7_bits_uop_pdst <= casez_tmp_246;
        else
          stq_7_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2685) begin
        if (_exe_tlb_uop_T_2)
          stq_7_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_7_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_7_bits_uop_pdst <= casez_tmp_246;
        else
          stq_7_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2461) begin
        if (_GEN_2141) begin
          if (_GEN_2044) begin
            if (_GEN_1660) begin
            end
            else
              stq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_7_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_7_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2461) begin
        if (_GEN_2141) begin
          if (_GEN_2044) begin
            if (_GEN_1660) begin
            end
            else begin
              stq_7_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_7_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_7_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_7_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_7_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_7_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_7_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_7_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_7_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_7_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_7_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_7_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_7_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_7_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_7_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_7_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_7_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_7_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_7_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_7_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_7_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_7_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_7_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_7_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_7_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_7_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_7_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_7_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_7_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_7_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_7_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_7_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_7_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_7_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_7_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_7_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_7_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_7_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_7_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_7_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_7_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_7_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_7_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_7_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_7_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_7_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2462) begin
        if (_GEN_2142) begin
          if (_GEN_2045) begin
            if (_GEN_1661) begin
            end
            else begin
              stq_8_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_8_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_8_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_8_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_8_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_8_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_8_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_8_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_8_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_8_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_8_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_8_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_8_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_8_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_8_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_8_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_8_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_8_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_8_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_8_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_8_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_8_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_8_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_8_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_8_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_8_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_8_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_8_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_8_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_8_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_8_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_8_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_8_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_8_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_8_valid)
        stq_8_bits_uop_br_mask <= stq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2462) begin
        if (_GEN_2142) begin
          if (_GEN_2045) begin
            if (_GEN_1661) begin
            end
            else
              stq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_8_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_8_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2462) begin
        if (_GEN_2142) begin
          if (_GEN_2045) begin
            if (_GEN_1661) begin
            end
            else begin
              stq_8_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_8_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_8_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_8_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_8_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_8_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_8_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_8_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_8_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_8_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_8_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_8_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_8_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_8_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_8_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_8_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_8_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_8_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_8_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_8_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_8_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_8_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_8_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_8_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_8_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_8_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_8_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_8_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_8_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_8_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2821) begin
        if (_exe_tlb_uop_T_9)
          stq_8_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_8_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_8_bits_uop_pdst <= casez_tmp_246;
        else
          stq_8_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2686) begin
        if (_exe_tlb_uop_T_2)
          stq_8_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_8_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_8_bits_uop_pdst <= casez_tmp_246;
        else
          stq_8_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2462) begin
        if (_GEN_2142) begin
          if (_GEN_2045) begin
            if (_GEN_1661) begin
            end
            else
              stq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_8_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_8_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2462) begin
        if (_GEN_2142) begin
          if (_GEN_2045) begin
            if (_GEN_1661) begin
            end
            else begin
              stq_8_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_8_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_8_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_8_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_8_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_8_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_8_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_8_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_8_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_8_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_8_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_8_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_8_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_8_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_8_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_8_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_8_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_8_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_8_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_8_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_8_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_8_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_8_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_8_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_8_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_8_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_8_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_8_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_8_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_8_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_8_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_8_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_8_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_8_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_8_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_8_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_8_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_8_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_8_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_8_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_8_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_8_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_8_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_8_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_8_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_8_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2463) begin
        if (_GEN_2143) begin
          if (_GEN_2046) begin
            if (_GEN_1662) begin
            end
            else begin
              stq_9_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_9_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_9_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_9_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_9_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_9_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_9_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_9_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_9_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_9_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_9_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_9_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_9_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_9_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_9_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_9_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_9_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_9_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_9_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_9_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_9_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_9_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_9_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_9_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_9_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_9_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_9_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_9_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_9_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_9_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_9_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_9_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_9_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_9_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_9_valid)
        stq_9_bits_uop_br_mask <= stq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2463) begin
        if (_GEN_2143) begin
          if (_GEN_2046) begin
            if (_GEN_1662) begin
            end
            else
              stq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_9_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_9_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2463) begin
        if (_GEN_2143) begin
          if (_GEN_2046) begin
            if (_GEN_1662) begin
            end
            else begin
              stq_9_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_9_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_9_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_9_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_9_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_9_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_9_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_9_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_9_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_9_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_9_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_9_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_9_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_9_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_9_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_9_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_9_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_9_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_9_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_9_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_9_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_9_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_9_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_9_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_9_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_9_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_9_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_9_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_9_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_9_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2823) begin
        if (_exe_tlb_uop_T_9)
          stq_9_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_9_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_9_bits_uop_pdst <= casez_tmp_246;
        else
          stq_9_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2687) begin
        if (_exe_tlb_uop_T_2)
          stq_9_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_9_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_9_bits_uop_pdst <= casez_tmp_246;
        else
          stq_9_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2463) begin
        if (_GEN_2143) begin
          if (_GEN_2046) begin
            if (_GEN_1662) begin
            end
            else
              stq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_9_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_9_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2463) begin
        if (_GEN_2143) begin
          if (_GEN_2046) begin
            if (_GEN_1662) begin
            end
            else begin
              stq_9_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_9_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_9_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_9_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_9_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_9_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_9_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_9_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_9_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_9_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_9_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_9_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_9_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_9_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_9_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_9_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_9_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_9_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_9_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_9_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_9_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_9_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_9_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_9_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_9_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_9_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_9_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_9_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_9_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_9_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_9_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_9_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_9_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_9_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_9_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_9_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_9_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_9_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_9_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_9_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_9_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_9_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_9_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_9_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_9_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_9_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2464) begin
        if (_GEN_2144) begin
          if (_GEN_2047) begin
            if (_GEN_1663) begin
            end
            else begin
              stq_10_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_10_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_10_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_10_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_10_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_10_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_10_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_10_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_10_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_10_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_10_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_10_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_10_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_10_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_10_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_10_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_10_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_10_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_10_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_10_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_10_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_10_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_10_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_10_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_10_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_10_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_10_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_10_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_10_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_10_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_10_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_10_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_10_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_10_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_10_valid)
        stq_10_bits_uop_br_mask <= stq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2464) begin
        if (_GEN_2144) begin
          if (_GEN_2047) begin
            if (_GEN_1663) begin
            end
            else
              stq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_10_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_10_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2464) begin
        if (_GEN_2144) begin
          if (_GEN_2047) begin
            if (_GEN_1663) begin
            end
            else begin
              stq_10_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_10_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_10_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_10_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_10_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_10_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_10_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_10_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_10_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_10_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_10_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_10_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_10_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_10_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_10_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_10_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_10_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_10_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_10_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_10_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_10_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_10_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_10_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_10_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_10_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_10_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_10_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_10_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_10_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_10_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2825) begin
        if (_exe_tlb_uop_T_9)
          stq_10_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_10_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_10_bits_uop_pdst <= casez_tmp_246;
        else
          stq_10_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2688) begin
        if (_exe_tlb_uop_T_2)
          stq_10_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_10_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_10_bits_uop_pdst <= casez_tmp_246;
        else
          stq_10_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2464) begin
        if (_GEN_2144) begin
          if (_GEN_2047) begin
            if (_GEN_1663) begin
            end
            else
              stq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_10_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_10_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2464) begin
        if (_GEN_2144) begin
          if (_GEN_2047) begin
            if (_GEN_1663) begin
            end
            else begin
              stq_10_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_10_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_10_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_10_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_10_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_10_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_10_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_10_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_10_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_10_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_10_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_10_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_10_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_10_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_10_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_10_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_10_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_10_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_10_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_10_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_10_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_10_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_10_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_10_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_10_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_10_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_10_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_10_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_10_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_10_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_10_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_10_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_10_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_10_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_10_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_10_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_10_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_10_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_10_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_10_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_10_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_10_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_10_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_10_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_10_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_10_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2465) begin
        if (_GEN_2145) begin
          if (_GEN_2048) begin
            if (_GEN_1664) begin
            end
            else begin
              stq_11_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_11_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_11_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_11_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_11_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_11_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_11_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_11_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_11_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_11_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_11_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_11_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_11_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_11_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_11_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_11_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_11_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_11_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_11_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_11_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_11_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_11_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_11_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_11_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_11_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_11_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_11_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_11_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_11_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_11_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_11_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_11_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_11_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_11_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_11_valid)
        stq_11_bits_uop_br_mask <= stq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2465) begin
        if (_GEN_2145) begin
          if (_GEN_2048) begin
            if (_GEN_1664) begin
            end
            else
              stq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_11_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_11_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2465) begin
        if (_GEN_2145) begin
          if (_GEN_2048) begin
            if (_GEN_1664) begin
            end
            else begin
              stq_11_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_11_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_11_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_11_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_11_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_11_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_11_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_11_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_11_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_11_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_11_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_11_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_11_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_11_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_11_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_11_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_11_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_11_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_11_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_11_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_11_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_11_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_11_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_11_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_11_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_11_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_11_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_11_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_11_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_11_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2827) begin
        if (_exe_tlb_uop_T_9)
          stq_11_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_11_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_11_bits_uop_pdst <= casez_tmp_246;
        else
          stq_11_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2689) begin
        if (_exe_tlb_uop_T_2)
          stq_11_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_11_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_11_bits_uop_pdst <= casez_tmp_246;
        else
          stq_11_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2465) begin
        if (_GEN_2145) begin
          if (_GEN_2048) begin
            if (_GEN_1664) begin
            end
            else
              stq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_11_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_11_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2465) begin
        if (_GEN_2145) begin
          if (_GEN_2048) begin
            if (_GEN_1664) begin
            end
            else begin
              stq_11_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_11_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_11_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_11_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_11_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_11_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_11_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_11_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_11_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_11_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_11_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_11_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_11_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_11_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_11_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_11_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_11_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_11_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_11_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_11_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_11_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_11_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_11_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_11_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_11_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_11_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_11_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_11_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_11_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_11_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_11_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_11_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_11_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_11_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_11_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_11_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_11_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_11_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_11_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_11_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_11_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_11_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_11_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_11_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_11_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_11_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2466) begin
        if (_GEN_2146) begin
          if (_GEN_2049) begin
            if (_GEN_1665) begin
            end
            else begin
              stq_12_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_12_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_12_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_12_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_12_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_12_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_12_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_12_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_12_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_12_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_12_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_12_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_12_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_12_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_12_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_12_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_12_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_12_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_12_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_12_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_12_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_12_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_12_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_12_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_12_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_12_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_12_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_12_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_12_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_12_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_12_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_12_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_12_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_12_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_12_valid)
        stq_12_bits_uop_br_mask <= stq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2466) begin
        if (_GEN_2146) begin
          if (_GEN_2049) begin
            if (_GEN_1665) begin
            end
            else
              stq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_12_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_12_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2466) begin
        if (_GEN_2146) begin
          if (_GEN_2049) begin
            if (_GEN_1665) begin
            end
            else begin
              stq_12_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_12_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_12_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_12_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_12_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_12_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_12_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_12_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_12_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_12_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_12_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_12_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_12_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_12_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_12_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_12_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_12_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_12_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_12_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_12_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_12_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_12_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_12_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_12_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_12_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_12_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_12_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_12_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_12_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_12_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2829) begin
        if (_exe_tlb_uop_T_9)
          stq_12_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_12_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_12_bits_uop_pdst <= casez_tmp_246;
        else
          stq_12_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2690) begin
        if (_exe_tlb_uop_T_2)
          stq_12_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_12_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_12_bits_uop_pdst <= casez_tmp_246;
        else
          stq_12_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2466) begin
        if (_GEN_2146) begin
          if (_GEN_2049) begin
            if (_GEN_1665) begin
            end
            else
              stq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_12_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_12_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2466) begin
        if (_GEN_2146) begin
          if (_GEN_2049) begin
            if (_GEN_1665) begin
            end
            else begin
              stq_12_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_12_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_12_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_12_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_12_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_12_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_12_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_12_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_12_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_12_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_12_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_12_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_12_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_12_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_12_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_12_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_12_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_12_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_12_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_12_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_12_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_12_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_12_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_12_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_12_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_12_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_12_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_12_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_12_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_12_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_12_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_12_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_12_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_12_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_12_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_12_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_12_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_12_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_12_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_12_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_12_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_12_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_12_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_12_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_12_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_12_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2467) begin
        if (_GEN_2147) begin
          if (_GEN_2050) begin
            if (_GEN_1666) begin
            end
            else begin
              stq_13_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_13_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_13_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_13_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_13_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_13_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_13_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_13_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_13_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_13_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_13_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_13_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_13_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_13_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_13_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_13_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_13_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_13_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_13_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_13_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_13_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_13_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_13_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_13_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_13_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_13_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_13_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_13_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_13_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_13_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_13_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_13_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_13_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_13_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_13_valid)
        stq_13_bits_uop_br_mask <= stq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2467) begin
        if (_GEN_2147) begin
          if (_GEN_2050) begin
            if (_GEN_1666) begin
            end
            else
              stq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_13_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_13_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2467) begin
        if (_GEN_2147) begin
          if (_GEN_2050) begin
            if (_GEN_1666) begin
            end
            else begin
              stq_13_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_13_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_13_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_13_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_13_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_13_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_13_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_13_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_13_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_13_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_13_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_13_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_13_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_13_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_13_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_13_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_13_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_13_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_13_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_13_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_13_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_13_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_13_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_13_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_13_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_13_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_13_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_13_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_13_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_13_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2831) begin
        if (_exe_tlb_uop_T_9)
          stq_13_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_13_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_13_bits_uop_pdst <= casez_tmp_246;
        else
          stq_13_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2691) begin
        if (_exe_tlb_uop_T_2)
          stq_13_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_13_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_13_bits_uop_pdst <= casez_tmp_246;
        else
          stq_13_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2467) begin
        if (_GEN_2147) begin
          if (_GEN_2050) begin
            if (_GEN_1666) begin
            end
            else
              stq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_13_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_13_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2467) begin
        if (_GEN_2147) begin
          if (_GEN_2050) begin
            if (_GEN_1666) begin
            end
            else begin
              stq_13_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_13_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_13_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_13_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_13_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_13_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_13_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_13_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_13_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_13_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_13_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_13_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_13_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_13_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_13_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_13_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_13_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_13_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_13_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_13_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_13_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_13_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_13_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_13_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_13_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_13_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_13_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_13_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_13_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_13_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_13_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_13_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_13_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_13_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_13_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_13_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_13_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_13_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_13_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_13_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_13_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_13_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_13_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_13_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_13_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_13_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2468) begin
        if (_GEN_2148) begin
          if (_GEN_2051) begin
            if (_GEN_1667) begin
            end
            else begin
              stq_14_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_14_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_14_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_14_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_14_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_14_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_14_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_14_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_14_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_14_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_14_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_14_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_14_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_14_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_14_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_14_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_14_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_14_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_14_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_14_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_14_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_14_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_14_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_14_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_14_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_14_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_14_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_14_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_14_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_14_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_14_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_14_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_14_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_14_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_14_valid)
        stq_14_bits_uop_br_mask <= stq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2468) begin
        if (_GEN_2148) begin
          if (_GEN_2051) begin
            if (_GEN_1667) begin
            end
            else
              stq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_14_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_14_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2468) begin
        if (_GEN_2148) begin
          if (_GEN_2051) begin
            if (_GEN_1667) begin
            end
            else begin
              stq_14_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_14_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_14_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_14_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_14_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_14_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_14_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_14_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_14_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_14_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_14_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_14_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_14_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_14_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_14_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_14_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_14_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_14_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_14_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_14_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_14_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_14_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_14_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_14_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_14_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_14_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_14_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_14_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_14_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_14_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2833) begin
        if (_exe_tlb_uop_T_9)
          stq_14_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_14_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_14_bits_uop_pdst <= casez_tmp_246;
        else
          stq_14_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2692) begin
        if (_exe_tlb_uop_T_2)
          stq_14_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_14_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_14_bits_uop_pdst <= casez_tmp_246;
        else
          stq_14_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2468) begin
        if (_GEN_2148) begin
          if (_GEN_2051) begin
            if (_GEN_1667) begin
            end
            else
              stq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_14_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_14_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2468) begin
        if (_GEN_2148) begin
          if (_GEN_2051) begin
            if (_GEN_1667) begin
            end
            else begin
              stq_14_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_14_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_14_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_14_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_14_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_14_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_14_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_14_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_14_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_14_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_14_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_14_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_14_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_14_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_14_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_14_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_14_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_14_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_14_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_14_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_14_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_14_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_14_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_14_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_14_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_14_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_14_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_14_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_14_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_14_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_14_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_14_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_14_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_14_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_14_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_14_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_14_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_14_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_14_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_14_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_14_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_14_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_14_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_14_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_14_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_14_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2469) begin
        if (_GEN_2149) begin
          if (_GEN_2052) begin
            if (_GEN_1668) begin
            end
            else begin
              stq_15_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_15_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_15_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_15_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_15_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_15_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_15_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_15_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_15_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_15_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_15_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_15_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_15_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_15_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_15_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_15_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_15_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_15_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_15_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_15_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_15_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_15_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_15_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_15_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_15_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_15_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_15_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_15_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_15_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_15_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_15_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_15_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_15_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_15_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_15_valid)
        stq_15_bits_uop_br_mask <= stq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2469) begin
        if (_GEN_2149) begin
          if (_GEN_2052) begin
            if (_GEN_1668) begin
            end
            else
              stq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_15_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_15_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2469) begin
        if (_GEN_2149) begin
          if (_GEN_2052) begin
            if (_GEN_1668) begin
            end
            else begin
              stq_15_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_15_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_15_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_15_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_15_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_15_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_15_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_15_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_15_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_15_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_15_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_15_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_15_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_15_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_15_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_15_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_15_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_15_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_15_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_15_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_15_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_15_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_15_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_15_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_15_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_15_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_15_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_15_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_15_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_15_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2835) begin
        if (_exe_tlb_uop_T_9)
          stq_15_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_15_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_15_bits_uop_pdst <= casez_tmp_246;
        else
          stq_15_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2693) begin
        if (_exe_tlb_uop_T_2)
          stq_15_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_15_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_15_bits_uop_pdst <= casez_tmp_246;
        else
          stq_15_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2469) begin
        if (_GEN_2149) begin
          if (_GEN_2052) begin
            if (_GEN_1668) begin
            end
            else
              stq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_15_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_15_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2469) begin
        if (_GEN_2149) begin
          if (_GEN_2052) begin
            if (_GEN_1668) begin
            end
            else begin
              stq_15_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_15_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_15_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_15_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_15_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_15_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_15_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_15_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_15_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_15_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_15_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_15_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_15_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_15_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_15_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_15_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_15_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_15_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_15_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_15_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_15_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_15_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_15_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_15_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_15_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_15_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_15_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_15_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_15_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_15_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_15_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_15_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_15_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_15_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_15_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_15_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_15_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_15_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_15_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_15_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_15_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_15_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_15_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_15_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_15_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_15_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2470) begin
        if (_GEN_2150) begin
          if (_GEN_2053) begin
            if (_GEN_1669) begin
            end
            else begin
              stq_16_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_16_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_16_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_16_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_16_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_16_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_16_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_16_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_16_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_16_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_16_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_16_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_16_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_16_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_16_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_16_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_16_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_16_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_16_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_16_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_16_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_16_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_16_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_16_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_16_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_16_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_16_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_16_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_16_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_16_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_16_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_16_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_16_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_16_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_16_valid)
        stq_16_bits_uop_br_mask <= stq_16_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2470) begin
        if (_GEN_2150) begin
          if (_GEN_2053) begin
            if (_GEN_1669) begin
            end
            else
              stq_16_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_16_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_16_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_16_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2470) begin
        if (_GEN_2150) begin
          if (_GEN_2053) begin
            if (_GEN_1669) begin
            end
            else begin
              stq_16_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_16_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_16_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_16_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_16_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_16_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_16_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_16_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_16_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_16_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_16_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_16_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_16_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_16_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_16_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_16_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_16_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_16_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_16_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_16_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_16_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_16_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_16_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_16_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_16_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_16_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_16_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_16_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_16_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_16_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_16_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_16_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_16_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_16_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_16_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_16_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2837) begin
        if (_exe_tlb_uop_T_9)
          stq_16_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_16_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_16_bits_uop_pdst <= casez_tmp_246;
        else
          stq_16_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2694) begin
        if (_exe_tlb_uop_T_2)
          stq_16_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_16_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_16_bits_uop_pdst <= casez_tmp_246;
        else
          stq_16_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2470) begin
        if (_GEN_2150) begin
          if (_GEN_2053) begin
            if (_GEN_1669) begin
            end
            else
              stq_16_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_16_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_16_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_16_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2470) begin
        if (_GEN_2150) begin
          if (_GEN_2053) begin
            if (_GEN_1669) begin
            end
            else begin
              stq_16_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_16_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_16_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_16_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_16_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_16_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_16_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_16_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_16_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_16_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_16_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_16_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_16_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_16_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_16_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_16_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_16_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_16_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_16_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_16_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_16_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_16_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_16_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_16_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_16_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_16_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_16_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_16_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_16_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_16_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_16_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_16_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_16_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_16_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_16_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_16_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_16_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_16_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_16_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_16_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_16_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_16_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_16_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_16_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_16_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_16_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_16_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_16_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_16_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_16_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_16_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_16_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_16_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_16_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_16_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_16_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_16_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_16_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2471) begin
        if (_GEN_2151) begin
          if (_GEN_2054) begin
            if (_GEN_1670) begin
            end
            else begin
              stq_17_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_17_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_17_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_17_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_17_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_17_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_17_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_17_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_17_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_17_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_17_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_17_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_17_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_17_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_17_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_17_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_17_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_17_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_17_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_17_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_17_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_17_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_17_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_17_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_17_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_17_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_17_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_17_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_17_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_17_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_17_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_17_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_17_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_17_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_17_valid)
        stq_17_bits_uop_br_mask <= stq_17_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2471) begin
        if (_GEN_2151) begin
          if (_GEN_2054) begin
            if (_GEN_1670) begin
            end
            else
              stq_17_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_17_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_17_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_17_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2471) begin
        if (_GEN_2151) begin
          if (_GEN_2054) begin
            if (_GEN_1670) begin
            end
            else begin
              stq_17_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_17_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_17_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_17_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_17_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_17_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_17_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_17_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_17_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_17_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_17_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_17_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_17_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_17_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_17_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_17_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_17_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_17_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_17_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_17_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_17_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_17_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_17_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_17_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_17_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_17_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_17_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_17_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_17_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_17_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_17_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_17_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_17_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_17_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_17_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_17_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2839) begin
        if (_exe_tlb_uop_T_9)
          stq_17_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_17_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_17_bits_uop_pdst <= casez_tmp_246;
        else
          stq_17_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2695) begin
        if (_exe_tlb_uop_T_2)
          stq_17_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_17_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_17_bits_uop_pdst <= casez_tmp_246;
        else
          stq_17_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2471) begin
        if (_GEN_2151) begin
          if (_GEN_2054) begin
            if (_GEN_1670) begin
            end
            else
              stq_17_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_17_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_17_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_17_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2471) begin
        if (_GEN_2151) begin
          if (_GEN_2054) begin
            if (_GEN_1670) begin
            end
            else begin
              stq_17_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_17_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_17_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_17_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_17_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_17_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_17_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_17_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_17_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_17_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_17_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_17_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_17_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_17_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_17_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_17_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_17_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_17_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_17_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_17_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_17_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_17_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_17_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_17_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_17_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_17_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_17_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_17_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_17_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_17_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_17_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_17_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_17_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_17_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_17_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_17_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_17_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_17_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_17_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_17_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_17_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_17_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_17_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_17_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_17_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_17_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_17_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_17_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_17_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_17_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_17_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_17_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_17_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_17_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_17_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_17_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_17_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_17_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2472) begin
        if (_GEN_2152) begin
          if (_GEN_2055) begin
            if (_GEN_1671) begin
            end
            else begin
              stq_18_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_18_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_18_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_18_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_18_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_18_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_18_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_18_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_18_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_18_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_18_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_18_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_18_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_18_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_18_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_18_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_18_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_18_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_18_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_18_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_18_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_18_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_18_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_18_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_18_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_18_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_18_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_18_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_18_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_18_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_18_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_18_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_18_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_18_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_18_valid)
        stq_18_bits_uop_br_mask <= stq_18_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2472) begin
        if (_GEN_2152) begin
          if (_GEN_2055) begin
            if (_GEN_1671) begin
            end
            else
              stq_18_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_18_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_18_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_18_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2472) begin
        if (_GEN_2152) begin
          if (_GEN_2055) begin
            if (_GEN_1671) begin
            end
            else begin
              stq_18_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_18_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_18_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_18_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_18_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_18_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_18_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_18_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_18_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_18_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_18_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_18_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_18_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_18_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_18_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_18_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_18_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_18_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_18_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_18_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_18_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_18_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_18_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_18_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_18_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_18_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_18_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_18_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_18_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_18_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_18_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_18_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_18_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_18_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_18_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_18_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2841) begin
        if (_exe_tlb_uop_T_9)
          stq_18_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_18_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_18_bits_uop_pdst <= casez_tmp_246;
        else
          stq_18_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2696) begin
        if (_exe_tlb_uop_T_2)
          stq_18_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_18_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_18_bits_uop_pdst <= casez_tmp_246;
        else
          stq_18_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2472) begin
        if (_GEN_2152) begin
          if (_GEN_2055) begin
            if (_GEN_1671) begin
            end
            else
              stq_18_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_18_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_18_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_18_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2472) begin
        if (_GEN_2152) begin
          if (_GEN_2055) begin
            if (_GEN_1671) begin
            end
            else begin
              stq_18_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_18_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_18_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_18_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_18_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_18_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_18_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_18_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_18_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_18_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_18_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_18_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_18_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_18_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_18_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_18_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_18_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_18_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_18_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_18_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_18_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_18_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_18_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_18_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_18_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_18_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_18_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_18_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_18_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_18_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_18_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_18_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_18_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_18_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_18_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_18_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_18_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_18_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_18_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_18_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_18_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_18_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_18_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_18_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_18_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_18_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_18_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_18_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_18_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_18_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_18_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_18_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_18_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_18_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_18_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_18_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_18_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_18_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2473) begin
        if (_GEN_2153) begin
          if (_GEN_2056) begin
            if (_GEN_1672) begin
            end
            else begin
              stq_19_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_19_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_19_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_19_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_19_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_19_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_19_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_19_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_19_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_19_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_19_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_19_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_19_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_19_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_19_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_19_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_19_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_19_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_19_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_19_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_19_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_19_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_19_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_19_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_19_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_19_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_19_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_19_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_19_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_19_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_19_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_19_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_19_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_19_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_19_valid)
        stq_19_bits_uop_br_mask <= stq_19_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2473) begin
        if (_GEN_2153) begin
          if (_GEN_2056) begin
            if (_GEN_1672) begin
            end
            else
              stq_19_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_19_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_19_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_19_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2473) begin
        if (_GEN_2153) begin
          if (_GEN_2056) begin
            if (_GEN_1672) begin
            end
            else begin
              stq_19_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_19_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_19_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_19_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_19_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_19_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_19_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_19_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_19_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_19_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_19_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_19_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_19_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_19_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_19_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_19_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_19_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_19_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_19_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_19_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_19_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_19_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_19_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_19_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_19_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_19_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_19_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_19_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_19_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_19_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_19_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_19_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_19_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_19_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_19_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_19_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2843) begin
        if (_exe_tlb_uop_T_9)
          stq_19_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_19_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_19_bits_uop_pdst <= casez_tmp_246;
        else
          stq_19_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2697) begin
        if (_exe_tlb_uop_T_2)
          stq_19_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_19_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_19_bits_uop_pdst <= casez_tmp_246;
        else
          stq_19_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2473) begin
        if (_GEN_2153) begin
          if (_GEN_2056) begin
            if (_GEN_1672) begin
            end
            else
              stq_19_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_19_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_19_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_19_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2473) begin
        if (_GEN_2153) begin
          if (_GEN_2056) begin
            if (_GEN_1672) begin
            end
            else begin
              stq_19_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_19_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_19_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_19_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_19_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_19_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_19_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_19_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_19_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_19_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_19_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_19_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_19_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_19_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_19_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_19_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_19_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_19_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_19_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_19_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_19_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_19_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_19_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_19_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_19_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_19_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_19_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_19_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_19_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_19_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_19_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_19_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_19_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_19_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_19_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_19_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_19_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_19_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_19_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_19_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_19_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_19_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_19_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_19_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_19_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_19_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_19_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_19_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_19_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_19_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_19_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_19_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_19_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_19_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_19_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_19_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_19_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_19_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2474) begin
        if (_GEN_2154) begin
          if (_GEN_2057) begin
            if (_GEN_1673) begin
            end
            else begin
              stq_20_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_20_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_20_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_20_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_20_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_20_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_20_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_20_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_20_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_20_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_20_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_20_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_20_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_20_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_20_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_20_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_20_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_20_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_20_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_20_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_20_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_20_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_20_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_20_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_20_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_20_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_20_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_20_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_20_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_20_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_20_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_20_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_20_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_20_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_20_valid)
        stq_20_bits_uop_br_mask <= stq_20_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2474) begin
        if (_GEN_2154) begin
          if (_GEN_2057) begin
            if (_GEN_1673) begin
            end
            else
              stq_20_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_20_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_20_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_20_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2474) begin
        if (_GEN_2154) begin
          if (_GEN_2057) begin
            if (_GEN_1673) begin
            end
            else begin
              stq_20_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_20_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_20_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_20_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_20_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_20_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_20_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_20_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_20_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_20_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_20_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_20_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_20_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_20_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_20_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_20_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_20_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_20_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_20_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_20_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_20_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_20_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_20_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_20_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_20_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_20_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_20_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_20_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_20_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_20_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_20_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_20_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_20_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_20_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_20_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_20_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2845) begin
        if (_exe_tlb_uop_T_9)
          stq_20_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_20_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_20_bits_uop_pdst <= casez_tmp_246;
        else
          stq_20_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2698) begin
        if (_exe_tlb_uop_T_2)
          stq_20_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_20_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_20_bits_uop_pdst <= casez_tmp_246;
        else
          stq_20_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2474) begin
        if (_GEN_2154) begin
          if (_GEN_2057) begin
            if (_GEN_1673) begin
            end
            else
              stq_20_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_20_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_20_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_20_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2474) begin
        if (_GEN_2154) begin
          if (_GEN_2057) begin
            if (_GEN_1673) begin
            end
            else begin
              stq_20_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_20_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_20_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_20_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_20_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_20_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_20_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_20_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_20_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_20_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_20_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_20_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_20_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_20_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_20_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_20_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_20_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_20_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_20_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_20_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_20_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_20_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_20_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_20_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_20_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_20_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_20_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_20_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_20_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_20_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_20_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_20_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_20_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_20_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_20_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_20_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_20_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_20_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_20_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_20_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_20_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_20_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_20_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_20_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_20_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_20_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_20_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_20_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_20_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_20_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_20_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_20_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_20_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_20_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_20_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_20_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_20_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_20_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2475) begin
        if (_GEN_2155) begin
          if (_GEN_2058) begin
            if (_GEN_1674) begin
            end
            else begin
              stq_21_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_21_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_21_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_21_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_21_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_21_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_21_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_21_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_21_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_21_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_21_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_21_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_21_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_21_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_21_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_21_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_21_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_21_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_21_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_21_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_21_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_21_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_21_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_21_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_21_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_21_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_21_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_21_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_21_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_21_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_21_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_21_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_21_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_21_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_21_valid)
        stq_21_bits_uop_br_mask <= stq_21_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2475) begin
        if (_GEN_2155) begin
          if (_GEN_2058) begin
            if (_GEN_1674) begin
            end
            else
              stq_21_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_21_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_21_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_21_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2475) begin
        if (_GEN_2155) begin
          if (_GEN_2058) begin
            if (_GEN_1674) begin
            end
            else begin
              stq_21_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_21_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_21_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_21_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_21_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_21_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_21_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_21_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_21_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_21_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_21_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_21_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_21_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_21_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_21_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_21_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_21_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_21_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_21_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_21_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_21_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_21_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_21_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_21_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_21_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_21_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_21_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_21_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_21_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_21_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_21_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_21_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_21_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_21_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_21_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_21_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2847) begin
        if (_exe_tlb_uop_T_9)
          stq_21_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_21_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_21_bits_uop_pdst <= casez_tmp_246;
        else
          stq_21_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2699) begin
        if (_exe_tlb_uop_T_2)
          stq_21_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_21_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_21_bits_uop_pdst <= casez_tmp_246;
        else
          stq_21_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2475) begin
        if (_GEN_2155) begin
          if (_GEN_2058) begin
            if (_GEN_1674) begin
            end
            else
              stq_21_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_21_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_21_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_21_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2475) begin
        if (_GEN_2155) begin
          if (_GEN_2058) begin
            if (_GEN_1674) begin
            end
            else begin
              stq_21_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_21_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_21_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_21_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_21_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_21_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_21_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_21_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_21_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_21_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_21_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_21_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_21_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_21_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_21_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_21_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_21_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_21_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_21_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_21_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_21_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_21_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_21_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_21_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_21_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_21_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_21_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_21_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_21_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_21_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_21_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_21_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_21_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_21_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_21_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_21_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_21_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_21_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_21_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_21_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_21_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_21_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_21_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_21_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_21_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_21_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_21_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_21_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_21_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_21_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_21_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_21_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_21_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_21_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_21_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_21_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_21_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_21_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2476) begin
        if (_GEN_2156) begin
          if (_GEN_2059) begin
            if (_GEN_1675) begin
            end
            else begin
              stq_22_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_22_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_22_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_22_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_22_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_22_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_22_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_22_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_22_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_22_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_22_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_22_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_22_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_22_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_22_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_22_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_22_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_22_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_22_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_22_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_22_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_22_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_22_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_22_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_22_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_22_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_22_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_22_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_22_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_22_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_22_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_22_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_22_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_22_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_22_valid)
        stq_22_bits_uop_br_mask <= stq_22_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2476) begin
        if (_GEN_2156) begin
          if (_GEN_2059) begin
            if (_GEN_1675) begin
            end
            else
              stq_22_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_22_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_22_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_22_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2476) begin
        if (_GEN_2156) begin
          if (_GEN_2059) begin
            if (_GEN_1675) begin
            end
            else begin
              stq_22_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_22_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_22_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_22_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_22_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_22_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_22_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_22_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_22_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_22_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_22_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_22_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_22_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_22_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_22_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_22_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_22_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_22_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_22_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_22_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_22_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_22_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_22_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_22_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_22_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_22_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_22_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_22_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_22_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_22_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_22_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_22_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_22_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_22_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_22_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_22_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2849) begin
        if (_exe_tlb_uop_T_9)
          stq_22_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_22_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_22_bits_uop_pdst <= casez_tmp_246;
        else
          stq_22_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2700) begin
        if (_exe_tlb_uop_T_2)
          stq_22_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_22_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_22_bits_uop_pdst <= casez_tmp_246;
        else
          stq_22_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2476) begin
        if (_GEN_2156) begin
          if (_GEN_2059) begin
            if (_GEN_1675) begin
            end
            else
              stq_22_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_22_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_22_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_22_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2476) begin
        if (_GEN_2156) begin
          if (_GEN_2059) begin
            if (_GEN_1675) begin
            end
            else begin
              stq_22_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_22_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_22_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_22_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_22_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_22_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_22_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_22_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_22_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_22_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_22_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_22_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_22_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_22_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_22_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_22_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_22_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_22_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_22_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_22_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_22_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_22_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_22_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_22_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_22_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_22_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_22_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_22_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_22_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_22_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_22_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_22_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_22_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_22_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_22_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_22_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_22_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_22_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_22_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_22_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_22_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_22_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_22_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_22_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_22_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_22_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_22_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_22_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_22_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_22_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_22_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_22_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_22_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_22_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_22_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_22_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_22_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_22_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2477) begin
        if (_GEN_2157) begin
          if (_GEN_2060) begin
            if (_GEN_1676) begin
            end
            else begin
              stq_23_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_23_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_23_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_23_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_23_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_23_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_23_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_23_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_23_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_23_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_23_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_23_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_23_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_23_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_23_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_23_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_23_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_23_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_23_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_23_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_23_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_23_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_23_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_23_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_23_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_23_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_23_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_23_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_23_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_23_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_23_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_23_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_23_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_23_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_23_valid)
        stq_23_bits_uop_br_mask <= stq_23_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2477) begin
        if (_GEN_2157) begin
          if (_GEN_2060) begin
            if (_GEN_1676) begin
            end
            else
              stq_23_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_23_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_23_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_23_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2477) begin
        if (_GEN_2157) begin
          if (_GEN_2060) begin
            if (_GEN_1676) begin
            end
            else begin
              stq_23_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_23_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_23_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_23_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_23_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_23_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_23_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_23_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_23_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_23_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_23_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_23_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_23_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_23_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_23_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_23_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_23_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_23_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_23_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_23_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_23_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_23_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_23_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_23_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_23_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_23_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_23_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_23_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_23_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_23_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_23_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_23_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_23_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_23_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_23_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_23_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2851) begin
        if (_exe_tlb_uop_T_9)
          stq_23_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_23_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_23_bits_uop_pdst <= casez_tmp_246;
        else
          stq_23_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2701) begin
        if (_exe_tlb_uop_T_2)
          stq_23_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_23_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_23_bits_uop_pdst <= casez_tmp_246;
        else
          stq_23_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2477) begin
        if (_GEN_2157) begin
          if (_GEN_2060) begin
            if (_GEN_1676) begin
            end
            else
              stq_23_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_23_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_23_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_23_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2477) begin
        if (_GEN_2157) begin
          if (_GEN_2060) begin
            if (_GEN_1676) begin
            end
            else begin
              stq_23_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_23_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_23_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_23_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_23_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_23_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_23_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_23_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_23_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_23_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_23_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_23_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_23_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_23_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_23_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_23_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_23_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_23_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_23_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_23_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_23_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_23_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_23_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_23_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_23_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_23_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_23_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_23_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_23_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_23_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_23_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_23_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_23_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_23_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_23_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_23_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_23_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_23_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_23_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_23_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_23_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_23_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_23_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_23_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_23_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_23_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_23_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_23_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_23_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_23_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_23_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_23_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_23_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_23_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_23_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_23_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_23_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_23_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2478) begin
        if (_GEN_2158) begin
          if (_GEN_2061) begin
            if (_GEN_1677) begin
            end
            else begin
              stq_24_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_24_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_24_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_24_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_24_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_24_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_24_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_24_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_24_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_24_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_24_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_24_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_24_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_24_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_24_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_24_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_24_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_24_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_24_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_24_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_24_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_24_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_24_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_24_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_24_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_24_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_24_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_24_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_24_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_24_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_24_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_24_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_24_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_24_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_24_valid)
        stq_24_bits_uop_br_mask <= stq_24_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2478) begin
        if (_GEN_2158) begin
          if (_GEN_2061) begin
            if (_GEN_1677) begin
            end
            else
              stq_24_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_24_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_24_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_24_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2478) begin
        if (_GEN_2158) begin
          if (_GEN_2061) begin
            if (_GEN_1677) begin
            end
            else begin
              stq_24_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_24_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_24_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_24_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_24_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_24_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_24_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_24_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_24_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_24_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_24_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_24_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_24_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_24_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_24_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_24_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_24_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_24_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_24_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_24_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_24_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_24_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_24_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_24_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_24_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_24_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_24_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_24_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_24_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_24_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_24_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_24_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_24_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_24_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_24_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_24_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2853) begin
        if (_exe_tlb_uop_T_9)
          stq_24_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_24_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_24_bits_uop_pdst <= casez_tmp_246;
        else
          stq_24_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2702) begin
        if (_exe_tlb_uop_T_2)
          stq_24_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_24_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_24_bits_uop_pdst <= casez_tmp_246;
        else
          stq_24_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2478) begin
        if (_GEN_2158) begin
          if (_GEN_2061) begin
            if (_GEN_1677) begin
            end
            else
              stq_24_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_24_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_24_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_24_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2478) begin
        if (_GEN_2158) begin
          if (_GEN_2061) begin
            if (_GEN_1677) begin
            end
            else begin
              stq_24_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_24_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_24_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_24_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_24_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_24_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_24_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_24_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_24_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_24_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_24_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_24_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_24_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_24_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_24_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_24_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_24_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_24_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_24_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_24_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_24_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_24_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_24_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_24_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_24_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_24_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_24_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_24_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_24_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_24_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_24_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_24_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_24_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_24_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_24_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_24_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_24_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_24_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_24_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_24_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_24_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_24_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_24_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_24_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_24_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_24_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_24_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_24_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_24_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_24_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_24_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_24_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_24_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_24_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_24_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_24_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_24_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_24_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2479) begin
        if (_GEN_2159) begin
          if (_GEN_2062) begin
            if (_GEN_1678) begin
            end
            else begin
              stq_25_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_25_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_25_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_25_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_25_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_25_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_25_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_25_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_25_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_25_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_25_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_25_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_25_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_25_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_25_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_25_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_25_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_25_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_25_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_25_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_25_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_25_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_25_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_25_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_25_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_25_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_25_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_25_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_25_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_25_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_25_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_25_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_25_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_25_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_25_valid)
        stq_25_bits_uop_br_mask <= stq_25_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2479) begin
        if (_GEN_2159) begin
          if (_GEN_2062) begin
            if (_GEN_1678) begin
            end
            else
              stq_25_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_25_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_25_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_25_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2479) begin
        if (_GEN_2159) begin
          if (_GEN_2062) begin
            if (_GEN_1678) begin
            end
            else begin
              stq_25_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_25_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_25_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_25_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_25_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_25_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_25_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_25_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_25_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_25_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_25_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_25_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_25_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_25_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_25_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_25_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_25_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_25_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_25_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_25_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_25_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_25_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_25_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_25_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_25_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_25_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_25_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_25_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_25_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_25_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_25_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_25_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_25_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_25_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_25_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_25_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2855) begin
        if (_exe_tlb_uop_T_9)
          stq_25_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_25_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_25_bits_uop_pdst <= casez_tmp_246;
        else
          stq_25_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2703) begin
        if (_exe_tlb_uop_T_2)
          stq_25_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_25_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_25_bits_uop_pdst <= casez_tmp_246;
        else
          stq_25_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2479) begin
        if (_GEN_2159) begin
          if (_GEN_2062) begin
            if (_GEN_1678) begin
            end
            else
              stq_25_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_25_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_25_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_25_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2479) begin
        if (_GEN_2159) begin
          if (_GEN_2062) begin
            if (_GEN_1678) begin
            end
            else begin
              stq_25_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_25_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_25_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_25_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_25_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_25_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_25_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_25_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_25_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_25_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_25_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_25_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_25_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_25_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_25_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_25_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_25_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_25_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_25_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_25_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_25_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_25_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_25_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_25_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_25_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_25_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_25_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_25_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_25_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_25_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_25_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_25_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_25_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_25_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_25_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_25_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_25_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_25_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_25_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_25_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_25_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_25_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_25_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_25_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_25_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_25_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_25_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_25_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_25_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_25_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_25_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_25_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_25_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_25_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_25_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_25_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_25_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_25_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2480) begin
        if (_GEN_2160) begin
          if (_GEN_2063) begin
            if (_GEN_1679) begin
            end
            else begin
              stq_26_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_26_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_26_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_26_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_26_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_26_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_26_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_26_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_26_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_26_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_26_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_26_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_26_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_26_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_26_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_26_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_26_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_26_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_26_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_26_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_26_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_26_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_26_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_26_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_26_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_26_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_26_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_26_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_26_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_26_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_26_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_26_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_26_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_26_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_26_valid)
        stq_26_bits_uop_br_mask <= stq_26_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2480) begin
        if (_GEN_2160) begin
          if (_GEN_2063) begin
            if (_GEN_1679) begin
            end
            else
              stq_26_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_26_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_26_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_26_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2480) begin
        if (_GEN_2160) begin
          if (_GEN_2063) begin
            if (_GEN_1679) begin
            end
            else begin
              stq_26_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_26_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_26_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_26_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_26_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_26_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_26_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_26_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_26_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_26_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_26_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_26_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_26_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_26_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_26_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_26_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_26_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_26_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_26_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_26_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_26_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_26_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_26_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_26_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_26_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_26_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_26_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_26_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_26_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_26_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_26_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_26_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_26_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_26_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_26_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_26_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2857) begin
        if (_exe_tlb_uop_T_9)
          stq_26_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_26_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_26_bits_uop_pdst <= casez_tmp_246;
        else
          stq_26_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2704) begin
        if (_exe_tlb_uop_T_2)
          stq_26_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_26_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_26_bits_uop_pdst <= casez_tmp_246;
        else
          stq_26_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2480) begin
        if (_GEN_2160) begin
          if (_GEN_2063) begin
            if (_GEN_1679) begin
            end
            else
              stq_26_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_26_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_26_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_26_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2480) begin
        if (_GEN_2160) begin
          if (_GEN_2063) begin
            if (_GEN_1679) begin
            end
            else begin
              stq_26_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_26_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_26_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_26_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_26_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_26_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_26_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_26_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_26_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_26_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_26_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_26_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_26_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_26_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_26_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_26_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_26_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_26_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_26_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_26_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_26_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_26_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_26_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_26_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_26_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_26_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_26_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_26_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_26_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_26_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_26_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_26_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_26_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_26_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_26_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_26_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_26_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_26_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_26_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_26_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_26_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_26_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_26_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_26_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_26_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_26_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_26_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_26_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_26_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_26_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_26_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_26_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_26_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_26_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_26_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_26_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_26_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_26_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2481) begin
        if (_GEN_2161) begin
          if (_GEN_2064) begin
            if (_GEN_1680) begin
            end
            else begin
              stq_27_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_27_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_27_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_27_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_27_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_27_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_27_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_27_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_27_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_27_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_27_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_27_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_27_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_27_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_27_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_27_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_27_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_27_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_27_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_27_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_27_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_27_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_27_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_27_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_27_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_27_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_27_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_27_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_27_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_27_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_27_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_27_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_27_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_27_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_27_valid)
        stq_27_bits_uop_br_mask <= stq_27_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2481) begin
        if (_GEN_2161) begin
          if (_GEN_2064) begin
            if (_GEN_1680) begin
            end
            else
              stq_27_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_27_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_27_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_27_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2481) begin
        if (_GEN_2161) begin
          if (_GEN_2064) begin
            if (_GEN_1680) begin
            end
            else begin
              stq_27_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_27_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_27_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_27_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_27_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_27_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_27_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_27_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_27_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_27_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_27_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_27_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_27_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_27_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_27_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_27_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_27_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_27_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_27_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_27_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_27_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_27_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_27_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_27_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_27_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_27_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_27_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_27_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_27_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_27_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_27_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_27_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_27_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_27_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_27_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_27_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2859) begin
        if (_exe_tlb_uop_T_9)
          stq_27_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_27_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_27_bits_uop_pdst <= casez_tmp_246;
        else
          stq_27_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2705) begin
        if (_exe_tlb_uop_T_2)
          stq_27_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_27_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_27_bits_uop_pdst <= casez_tmp_246;
        else
          stq_27_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2481) begin
        if (_GEN_2161) begin
          if (_GEN_2064) begin
            if (_GEN_1680) begin
            end
            else
              stq_27_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_27_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_27_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_27_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2481) begin
        if (_GEN_2161) begin
          if (_GEN_2064) begin
            if (_GEN_1680) begin
            end
            else begin
              stq_27_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_27_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_27_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_27_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_27_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_27_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_27_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_27_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_27_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_27_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_27_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_27_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_27_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_27_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_27_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_27_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_27_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_27_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_27_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_27_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_27_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_27_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_27_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_27_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_27_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_27_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_27_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_27_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_27_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_27_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_27_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_27_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_27_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_27_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_27_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_27_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_27_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_27_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_27_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_27_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_27_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_27_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_27_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_27_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_27_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_27_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_27_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_27_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_27_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_27_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_27_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_27_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_27_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_27_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_27_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_27_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_27_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_27_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2482) begin
        if (_GEN_2162) begin
          if (_GEN_2065) begin
            if (_GEN_1681) begin
            end
            else begin
              stq_28_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_28_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_28_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_28_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_28_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_28_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_28_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_28_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_28_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_28_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_28_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_28_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_28_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_28_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_28_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_28_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_28_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_28_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_28_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_28_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_28_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_28_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_28_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_28_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_28_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_28_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_28_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_28_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_28_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_28_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_28_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_28_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_28_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_28_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_28_valid)
        stq_28_bits_uop_br_mask <= stq_28_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2482) begin
        if (_GEN_2162) begin
          if (_GEN_2065) begin
            if (_GEN_1681) begin
            end
            else
              stq_28_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_28_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_28_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_28_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2482) begin
        if (_GEN_2162) begin
          if (_GEN_2065) begin
            if (_GEN_1681) begin
            end
            else begin
              stq_28_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_28_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_28_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_28_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_28_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_28_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_28_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_28_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_28_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_28_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_28_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_28_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_28_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_28_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_28_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_28_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_28_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_28_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_28_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_28_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_28_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_28_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_28_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_28_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_28_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_28_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_28_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_28_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_28_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_28_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_28_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_28_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_28_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_28_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_28_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_28_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2861) begin
        if (_exe_tlb_uop_T_9)
          stq_28_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_28_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_28_bits_uop_pdst <= casez_tmp_246;
        else
          stq_28_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2706) begin
        if (_exe_tlb_uop_T_2)
          stq_28_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_28_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_28_bits_uop_pdst <= casez_tmp_246;
        else
          stq_28_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2482) begin
        if (_GEN_2162) begin
          if (_GEN_2065) begin
            if (_GEN_1681) begin
            end
            else
              stq_28_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_28_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_28_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_28_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2482) begin
        if (_GEN_2162) begin
          if (_GEN_2065) begin
            if (_GEN_1681) begin
            end
            else begin
              stq_28_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_28_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_28_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_28_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_28_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_28_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_28_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_28_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_28_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_28_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_28_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_28_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_28_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_28_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_28_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_28_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_28_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_28_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_28_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_28_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_28_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_28_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_28_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_28_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_28_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_28_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_28_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_28_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_28_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_28_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_28_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_28_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_28_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_28_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_28_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_28_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_28_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_28_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_28_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_28_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_28_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_28_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_28_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_28_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_28_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_28_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_28_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_28_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_28_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_28_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_28_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_28_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_28_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_28_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_28_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_28_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_28_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_28_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2483) begin
        if (_GEN_2163) begin
          if (_GEN_2066) begin
            if (_GEN_1682) begin
            end
            else begin
              stq_29_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_29_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_29_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_29_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_29_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_29_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_29_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_29_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_29_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_29_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_29_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_29_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_29_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_29_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_29_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_29_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_29_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_29_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_29_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_29_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_29_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_29_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_29_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_29_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_29_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_29_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_29_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_29_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_29_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_29_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_29_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_29_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_29_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_29_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_29_valid)
        stq_29_bits_uop_br_mask <= stq_29_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2483) begin
        if (_GEN_2163) begin
          if (_GEN_2066) begin
            if (_GEN_1682) begin
            end
            else
              stq_29_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_29_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_29_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_29_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2483) begin
        if (_GEN_2163) begin
          if (_GEN_2066) begin
            if (_GEN_1682) begin
            end
            else begin
              stq_29_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_29_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_29_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_29_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_29_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_29_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_29_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_29_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_29_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_29_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_29_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_29_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_29_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_29_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_29_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_29_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_29_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_29_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_29_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_29_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_29_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_29_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_29_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_29_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_29_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_29_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_29_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_29_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_29_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_29_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_29_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_29_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_29_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_29_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_29_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_29_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2863) begin
        if (_exe_tlb_uop_T_9)
          stq_29_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_29_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_29_bits_uop_pdst <= casez_tmp_246;
        else
          stq_29_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2707) begin
        if (_exe_tlb_uop_T_2)
          stq_29_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_29_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_29_bits_uop_pdst <= casez_tmp_246;
        else
          stq_29_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2483) begin
        if (_GEN_2163) begin
          if (_GEN_2066) begin
            if (_GEN_1682) begin
            end
            else
              stq_29_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_29_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_29_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_29_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2483) begin
        if (_GEN_2163) begin
          if (_GEN_2066) begin
            if (_GEN_1682) begin
            end
            else begin
              stq_29_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_29_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_29_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_29_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_29_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_29_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_29_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_29_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_29_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_29_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_29_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_29_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_29_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_29_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_29_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_29_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_29_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_29_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_29_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_29_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_29_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_29_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_29_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_29_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_29_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_29_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_29_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_29_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_29_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_29_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_29_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_29_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_29_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_29_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_29_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_29_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_29_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_29_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_29_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_29_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_29_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_29_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_29_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_29_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_29_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_29_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_29_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_29_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_29_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_29_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_29_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_29_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_29_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_29_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_29_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_29_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_29_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_29_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2484) begin
        if (_GEN_2164) begin
          if (_GEN_2067) begin
            if (_GEN_1683) begin
            end
            else begin
              stq_30_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_30_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_30_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_30_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_30_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_30_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_30_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_30_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_30_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_30_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_30_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_30_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_30_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_30_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_30_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_30_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_30_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_30_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_30_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_30_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_30_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_30_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_30_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_30_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_30_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_30_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_30_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_30_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_30_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_30_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_30_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_30_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_30_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_30_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_30_valid)
        stq_30_bits_uop_br_mask <= stq_30_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2484) begin
        if (_GEN_2164) begin
          if (_GEN_2067) begin
            if (_GEN_1683) begin
            end
            else
              stq_30_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_30_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_30_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_30_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2484) begin
        if (_GEN_2164) begin
          if (_GEN_2067) begin
            if (_GEN_1683) begin
            end
            else begin
              stq_30_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_30_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_30_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_30_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_30_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_30_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_30_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_30_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_30_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_30_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_30_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_30_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_30_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_30_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_30_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_30_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_30_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_30_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_30_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_30_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_30_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_30_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_30_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_30_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_30_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_30_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_30_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_30_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_30_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_30_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_30_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_30_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_30_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_30_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_30_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_30_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2865) begin
        if (_exe_tlb_uop_T_9)
          stq_30_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_30_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_30_bits_uop_pdst <= casez_tmp_246;
        else
          stq_30_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2708) begin
        if (_exe_tlb_uop_T_2)
          stq_30_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_30_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_30_bits_uop_pdst <= casez_tmp_246;
        else
          stq_30_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2484) begin
        if (_GEN_2164) begin
          if (_GEN_2067) begin
            if (_GEN_1683) begin
            end
            else
              stq_30_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_30_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_30_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_30_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2484) begin
        if (_GEN_2164) begin
          if (_GEN_2067) begin
            if (_GEN_1683) begin
            end
            else begin
              stq_30_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_30_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_30_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_30_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_30_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_30_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_30_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_30_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_30_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_30_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_30_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_30_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_30_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_30_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_30_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_30_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_30_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_30_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_30_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_30_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_30_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_30_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_30_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_30_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_30_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_30_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_30_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_30_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_30_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_30_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_30_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_30_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_30_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_30_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_30_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_30_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_30_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_30_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_30_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_30_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_30_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_30_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_30_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_30_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_30_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_30_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_30_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_30_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_30_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_30_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_30_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_30_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_30_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_30_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_30_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_30_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_30_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_30_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (_GEN_2485) begin
        if (_GEN_2165) begin
          if (_GEN_2068) begin
            if (_GEN_1684) begin
            end
            else begin
              stq_31_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
              stq_31_bits_uop_inst <= io_core_dis_uops_0_bits_inst;
              stq_31_bits_uop_debug_inst <= io_core_dis_uops_0_bits_debug_inst;
              stq_31_bits_uop_debug_pc <= io_core_dis_uops_0_bits_debug_pc;
              stq_31_bits_uop_iq_type <= io_core_dis_uops_0_bits_iq_type;
              stq_31_bits_uop_fu_code <= io_core_dis_uops_0_bits_fu_code;
              stq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_0_bits_ctrl_br_type;
              stq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_0_bits_ctrl_op1_sel;
              stq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_0_bits_ctrl_op2_sel;
              stq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_0_bits_ctrl_imm_sel;
              stq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_0_bits_ctrl_op_fcn;
              stq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_0_bits_ctrl_csr_cmd;
              stq_31_bits_uop_iw_state <= io_core_dis_uops_0_bits_iw_state;
            end
          end
          else begin
            stq_31_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
            stq_31_bits_uop_inst <= io_core_dis_uops_1_bits_inst;
            stq_31_bits_uop_debug_inst <= io_core_dis_uops_1_bits_debug_inst;
            stq_31_bits_uop_debug_pc <= io_core_dis_uops_1_bits_debug_pc;
            stq_31_bits_uop_iq_type <= io_core_dis_uops_1_bits_iq_type;
            stq_31_bits_uop_fu_code <= io_core_dis_uops_1_bits_fu_code;
            stq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_1_bits_ctrl_br_type;
            stq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_1_bits_ctrl_op1_sel;
            stq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_1_bits_ctrl_op2_sel;
            stq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_1_bits_ctrl_imm_sel;
            stq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_1_bits_ctrl_op_fcn;
            stq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_1_bits_ctrl_csr_cmd;
            stq_31_bits_uop_iw_state <= io_core_dis_uops_1_bits_iw_state;
          end
        end
        else begin
          stq_31_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
          stq_31_bits_uop_inst <= io_core_dis_uops_2_bits_inst;
          stq_31_bits_uop_debug_inst <= io_core_dis_uops_2_bits_debug_inst;
          stq_31_bits_uop_debug_pc <= io_core_dis_uops_2_bits_debug_pc;
          stq_31_bits_uop_iq_type <= io_core_dis_uops_2_bits_iq_type;
          stq_31_bits_uop_fu_code <= io_core_dis_uops_2_bits_fu_code;
          stq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_2_bits_ctrl_br_type;
          stq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_2_bits_ctrl_op1_sel;
          stq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_2_bits_ctrl_op2_sel;
          stq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_2_bits_ctrl_imm_sel;
          stq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_2_bits_ctrl_op_fcn;
          stq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_2_bits_ctrl_csr_cmd;
          stq_31_bits_uop_iw_state <= io_core_dis_uops_2_bits_iw_state;
        end
      end
      else begin
        stq_31_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
        stq_31_bits_uop_inst <= io_core_dis_uops_3_bits_inst;
        stq_31_bits_uop_debug_inst <= io_core_dis_uops_3_bits_debug_inst;
        stq_31_bits_uop_debug_pc <= io_core_dis_uops_3_bits_debug_pc;
        stq_31_bits_uop_iq_type <= io_core_dis_uops_3_bits_iq_type;
        stq_31_bits_uop_fu_code <= io_core_dis_uops_3_bits_fu_code;
        stq_31_bits_uop_ctrl_br_type <= io_core_dis_uops_3_bits_ctrl_br_type;
        stq_31_bits_uop_ctrl_op1_sel <= io_core_dis_uops_3_bits_ctrl_op1_sel;
        stq_31_bits_uop_ctrl_op2_sel <= io_core_dis_uops_3_bits_ctrl_op2_sel;
        stq_31_bits_uop_ctrl_imm_sel <= io_core_dis_uops_3_bits_ctrl_imm_sel;
        stq_31_bits_uop_ctrl_op_fcn <= io_core_dis_uops_3_bits_ctrl_op_fcn;
        stq_31_bits_uop_ctrl_csr_cmd <= io_core_dis_uops_3_bits_ctrl_csr_cmd;
        stq_31_bits_uop_iw_state <= io_core_dis_uops_3_bits_iw_state;
      end
      if (stq_31_valid)
        stq_31_bits_uop_br_mask <= stq_31_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_2485) begin
        if (_GEN_2165) begin
          if (_GEN_2068) begin
            if (_GEN_1684) begin
            end
            else
              stq_31_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_31_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_31_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_31_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_2485) begin
        if (_GEN_2165) begin
          if (_GEN_2068) begin
            if (_GEN_1684) begin
            end
            else begin
              stq_31_bits_uop_br_tag <= io_core_dis_uops_0_bits_br_tag;
              stq_31_bits_uop_ftq_idx <= io_core_dis_uops_0_bits_ftq_idx;
              stq_31_bits_uop_pc_lob <= io_core_dis_uops_0_bits_pc_lob;
              stq_31_bits_uop_imm_packed <= io_core_dis_uops_0_bits_imm_packed;
              stq_31_bits_uop_csr_addr <= io_core_dis_uops_0_bits_csr_addr;
              stq_31_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_31_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_31_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
              stq_31_bits_uop_rxq_idx <= io_core_dis_uops_0_bits_rxq_idx;
            end
          end
          else begin
            stq_31_bits_uop_br_tag <= io_core_dis_uops_1_bits_br_tag;
            stq_31_bits_uop_ftq_idx <= io_core_dis_uops_1_bits_ftq_idx;
            stq_31_bits_uop_pc_lob <= io_core_dis_uops_1_bits_pc_lob;
            stq_31_bits_uop_imm_packed <= io_core_dis_uops_1_bits_imm_packed;
            stq_31_bits_uop_csr_addr <= io_core_dis_uops_1_bits_csr_addr;
            stq_31_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_31_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_31_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
            stq_31_bits_uop_rxq_idx <= io_core_dis_uops_1_bits_rxq_idx;
          end
        end
        else begin
          stq_31_bits_uop_br_tag <= io_core_dis_uops_2_bits_br_tag;
          stq_31_bits_uop_ftq_idx <= io_core_dis_uops_2_bits_ftq_idx;
          stq_31_bits_uop_pc_lob <= io_core_dis_uops_2_bits_pc_lob;
          stq_31_bits_uop_imm_packed <= io_core_dis_uops_2_bits_imm_packed;
          stq_31_bits_uop_csr_addr <= io_core_dis_uops_2_bits_csr_addr;
          stq_31_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_31_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_31_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
          stq_31_bits_uop_rxq_idx <= io_core_dis_uops_2_bits_rxq_idx;
        end
      end
      else begin
        stq_31_bits_uop_br_tag <= io_core_dis_uops_3_bits_br_tag;
        stq_31_bits_uop_ftq_idx <= io_core_dis_uops_3_bits_ftq_idx;
        stq_31_bits_uop_pc_lob <= io_core_dis_uops_3_bits_pc_lob;
        stq_31_bits_uop_imm_packed <= io_core_dis_uops_3_bits_imm_packed;
        stq_31_bits_uop_csr_addr <= io_core_dis_uops_3_bits_csr_addr;
        stq_31_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_31_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_31_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
        stq_31_bits_uop_rxq_idx <= io_core_dis_uops_3_bits_rxq_idx;
      end
      if (_GEN_2867) begin
        if (_exe_tlb_uop_T_9)
          stq_31_bits_uop_pdst <= _mem_incoming_uop_WIRE_1_pdst;
        else if (will_fire_load_retry_1_will_fire)
          stq_31_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_1_will_fire)
          stq_31_bits_uop_pdst <= casez_tmp_246;
        else
          stq_31_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2709) begin
        if (_exe_tlb_uop_T_2)
          stq_31_bits_uop_pdst <= _mem_incoming_uop_WIRE_0_pdst;
        else if (will_fire_load_retry_0_will_fire)
          stq_31_bits_uop_pdst <= casez_tmp_160;
        else if (will_fire_sta_retry_0_will_fire)
          stq_31_bits_uop_pdst <= casez_tmp_246;
        else
          stq_31_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_2485) begin
        if (_GEN_2165) begin
          if (_GEN_2068) begin
            if (_GEN_1684) begin
            end
            else
              stq_31_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_31_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_31_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_31_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_2485) begin
        if (_GEN_2165) begin
          if (_GEN_2068) begin
            if (_GEN_1684) begin
            end
            else begin
              stq_31_bits_uop_prs1 <= io_core_dis_uops_0_bits_prs1;
              stq_31_bits_uop_prs2 <= io_core_dis_uops_0_bits_prs2;
              stq_31_bits_uop_prs3 <= io_core_dis_uops_0_bits_prs3;
              stq_31_bits_uop_stale_pdst <= io_core_dis_uops_0_bits_stale_pdst;
              stq_31_bits_uop_exc_cause <= io_core_dis_uops_0_bits_exc_cause;
              stq_31_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_31_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_31_bits_uop_ldst <= io_core_dis_uops_0_bits_ldst;
              stq_31_bits_uop_lrs1 <= io_core_dis_uops_0_bits_lrs1;
              stq_31_bits_uop_lrs2 <= io_core_dis_uops_0_bits_lrs2;
              stq_31_bits_uop_lrs3 <= io_core_dis_uops_0_bits_lrs3;
              stq_31_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
              stq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_0_bits_lrs1_rtype;
              stq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_0_bits_lrs2_rtype;
              stq_31_bits_uop_debug_fsrc <= io_core_dis_uops_0_bits_debug_fsrc;
              stq_31_bits_uop_debug_tsrc <= io_core_dis_uops_0_bits_debug_tsrc;
            end
          end
          else begin
            stq_31_bits_uop_prs1 <= io_core_dis_uops_1_bits_prs1;
            stq_31_bits_uop_prs2 <= io_core_dis_uops_1_bits_prs2;
            stq_31_bits_uop_prs3 <= io_core_dis_uops_1_bits_prs3;
            stq_31_bits_uop_stale_pdst <= io_core_dis_uops_1_bits_stale_pdst;
            stq_31_bits_uop_exc_cause <= io_core_dis_uops_1_bits_exc_cause;
            stq_31_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_31_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_31_bits_uop_ldst <= io_core_dis_uops_1_bits_ldst;
            stq_31_bits_uop_lrs1 <= io_core_dis_uops_1_bits_lrs1;
            stq_31_bits_uop_lrs2 <= io_core_dis_uops_1_bits_lrs2;
            stq_31_bits_uop_lrs3 <= io_core_dis_uops_1_bits_lrs3;
            stq_31_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
            stq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_1_bits_lrs1_rtype;
            stq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_1_bits_lrs2_rtype;
            stq_31_bits_uop_debug_fsrc <= io_core_dis_uops_1_bits_debug_fsrc;
            stq_31_bits_uop_debug_tsrc <= io_core_dis_uops_1_bits_debug_tsrc;
          end
        end
        else begin
          stq_31_bits_uop_prs1 <= io_core_dis_uops_2_bits_prs1;
          stq_31_bits_uop_prs2 <= io_core_dis_uops_2_bits_prs2;
          stq_31_bits_uop_prs3 <= io_core_dis_uops_2_bits_prs3;
          stq_31_bits_uop_stale_pdst <= io_core_dis_uops_2_bits_stale_pdst;
          stq_31_bits_uop_exc_cause <= io_core_dis_uops_2_bits_exc_cause;
          stq_31_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_31_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_31_bits_uop_ldst <= io_core_dis_uops_2_bits_ldst;
          stq_31_bits_uop_lrs1 <= io_core_dis_uops_2_bits_lrs1;
          stq_31_bits_uop_lrs2 <= io_core_dis_uops_2_bits_lrs2;
          stq_31_bits_uop_lrs3 <= io_core_dis_uops_2_bits_lrs3;
          stq_31_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
          stq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_2_bits_lrs1_rtype;
          stq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_2_bits_lrs2_rtype;
          stq_31_bits_uop_debug_fsrc <= io_core_dis_uops_2_bits_debug_fsrc;
          stq_31_bits_uop_debug_tsrc <= io_core_dis_uops_2_bits_debug_tsrc;
        end
      end
      else begin
        stq_31_bits_uop_prs1 <= io_core_dis_uops_3_bits_prs1;
        stq_31_bits_uop_prs2 <= io_core_dis_uops_3_bits_prs2;
        stq_31_bits_uop_prs3 <= io_core_dis_uops_3_bits_prs3;
        stq_31_bits_uop_stale_pdst <= io_core_dis_uops_3_bits_stale_pdst;
        stq_31_bits_uop_exc_cause <= io_core_dis_uops_3_bits_exc_cause;
        stq_31_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_31_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_31_bits_uop_ldst <= io_core_dis_uops_3_bits_ldst;
        stq_31_bits_uop_lrs1 <= io_core_dis_uops_3_bits_lrs1;
        stq_31_bits_uop_lrs2 <= io_core_dis_uops_3_bits_lrs2;
        stq_31_bits_uop_lrs3 <= io_core_dis_uops_3_bits_lrs3;
        stq_31_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
        stq_31_bits_uop_lrs1_rtype <= io_core_dis_uops_3_bits_lrs1_rtype;
        stq_31_bits_uop_lrs2_rtype <= io_core_dis_uops_3_bits_lrs2_rtype;
        stq_31_bits_uop_debug_fsrc <= io_core_dis_uops_3_bits_debug_fsrc;
        stq_31_bits_uop_debug_tsrc <= io_core_dis_uops_3_bits_debug_tsrc;
      end
      if (clear_store)
        stq_head <= stq_head + 5'h1;
      if (commit_store_3)
        stq_commit_head <= _GEN_1555 + 5'h1;
      else if (commit_store_2)
        stq_commit_head <= _GEN_1554;
      else if (commit_store_1)
        stq_commit_head <= _GEN_1549;
      else if (commit_store)
        stq_commit_head <= _GEN_1544;
      if (clear_store & casez_tmp_544)
        stq_execute_head <= stq_execute_head + 5'h1;
      else if (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | io_dmem_nack_1_bits_uop_uses_ldq | io_dmem_nack_1_bits_uop_stq_idx < stq_head ^ _GEN_1587 ^ io_dmem_nack_1_bits_uop_stq_idx >= stq_execute_head) begin
        if (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | io_dmem_nack_0_bits_uop_uses_ldq | io_dmem_nack_0_bits_uop_stq_idx < stq_head ^ _GEN_1587 ^ io_dmem_nack_0_bits_uop_stq_idx >= stq_execute_head) begin
          if (_GEN_281 | ~will_fire_store_commit_1_will_fire) begin
            if (_GEN_275 | ~(will_fire_store_commit_0_will_fire & dmem_req_fire_0)) begin
            end
            else
              stq_execute_head <= stq_execute_head + 5'h1;
          end
          else if (dmem_req_fire_1)
            stq_execute_head <= stq_execute_head + 5'h1;
        end
        else
          stq_execute_head <= io_dmem_nack_0_bits_uop_stq_idx;
      end
      else
        stq_execute_head <= io_dmem_nack_1_bits_uop_stq_idx;
    end
    stq_0_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_0_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_0_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_0_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_0_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_0_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_0_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_0_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_0_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_0_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_0_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_0_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_0_bits_uop_taken <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_0_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_0_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_0_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_0_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2454 & _GEN_2134 & _GEN_2037 & _GEN_1653 & stq_0_bits_uop_ppred_busy;
    stq_0_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h0 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h0 | (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_0_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_0_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_0_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_0_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_0_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_0_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_0_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_0_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_0_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_0_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_0_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_0_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_0_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_0_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_0_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_0_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_0_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_0_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_0_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_0_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2454 ? (_GEN_2134 ? (_GEN_2037 ? (_GEN_1653 ? stq_0_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_0_bits_addr_valid <= ~_GEN_5752 & (clear_store ? ~_GEN_5654 & _GEN_2806 : ~_GEN_5208 & _GEN_2806);
    if (_GEN_2805) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_0_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_0_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_0_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_0_bits_addr_bits <= casez_tmp_290;
        else
          stq_0_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_0_bits_addr_bits <= _GEN_280;
      stq_0_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2678) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_0_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_0_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_0_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_0_bits_addr_bits <= casez_tmp_290;
        else
          stq_0_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_0_bits_addr_bits <= _GEN_274;
      stq_0_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_0_bits_data_valid <= ~_GEN_5752 & (clear_store ? ~_GEN_5654 & _GEN_2870 : ~_GEN_5208 & _GEN_2870);
    if (_stq_bits_data_bits_T_2 & _GEN_2869)
      stq_0_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2710)
      stq_0_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_0_bits_committed <= ~_GEN_5716 & (commit_store_3 ? _GEN_5590 | _GEN_5496 | _GEN_5401 : _GEN_5496 | _GEN_5401);
    stq_0_bits_succeeded <= ~_GEN_5716 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h0 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h0 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2583)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2583)) & _GEN_2454 & _GEN_2134 & _GEN_2037 & _GEN_1653 & stq_0_bits_succeeded);
    stq_1_valid <= ~_GEN_5754 & (clear_store ? ~_GEN_5656 & _GEN_2393 : ~_GEN_5209 & _GEN_2393);
    stq_1_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_1_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_1_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_1_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_1_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_1_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_1_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_1_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_1_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_1_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_1_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_1_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_1_bits_uop_taken <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_1_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_1_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_1_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_1_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2455 & _GEN_2135 & _GEN_2038 & _GEN_1654 & stq_1_bits_uop_ppred_busy;
    stq_1_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1 | (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_1_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_1_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_1_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_1_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_1_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_1_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_1_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_1_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_1_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_1_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_1_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_1_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_1_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_1_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_1_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_1_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_1_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_1_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_1_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_1_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2455 ? (_GEN_2135 ? (_GEN_2038 ? (_GEN_1654 ? stq_1_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_1_bits_addr_valid <= ~_GEN_5754 & (clear_store ? ~_GEN_5656 & _GEN_2808 : ~_GEN_5209 & _GEN_2808);
    if (_GEN_2807) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_1_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_1_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_1_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_1_bits_addr_bits <= casez_tmp_290;
        else
          stq_1_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_1_bits_addr_bits <= _GEN_280;
      stq_1_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2679) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_1_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_1_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_1_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_1_bits_addr_bits <= casez_tmp_290;
        else
          stq_1_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_1_bits_addr_bits <= _GEN_274;
      stq_1_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_1_bits_data_valid <= ~_GEN_5754 & (clear_store ? ~_GEN_5656 & _GEN_2872 : ~_GEN_5209 & _GEN_2872);
    if (_stq_bits_data_bits_T_2 & _GEN_2871)
      stq_1_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2711)
      stq_1_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_1_bits_committed <= ~_GEN_5717 & (commit_store_3 ? _GEN_5591 | _GEN_5498 | _GEN_5403 : _GEN_5498 | _GEN_5403);
    stq_1_bits_succeeded <= ~_GEN_5717 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2584)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2584)) & _GEN_2455 & _GEN_2135 & _GEN_2038 & _GEN_1654 & stq_1_bits_succeeded);
    stq_2_valid <= ~_GEN_5756 & (clear_store ? ~_GEN_5658 & _GEN_2395 : ~_GEN_5210 & _GEN_2395);
    stq_2_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_2_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_2_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_2_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_2_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_2_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_2_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_2_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_2_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_2_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_2_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_2_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_2_bits_uop_taken <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_2_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_2_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_2_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_2_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2456 & _GEN_2136 & _GEN_2039 & _GEN_1655 & stq_2_bits_uop_ppred_busy;
    stq_2_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h2 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h2 | (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_2_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_2_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_2_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_2_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_2_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_2_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_2_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_2_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_2_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_2_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_2_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_2_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_2_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_2_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_2_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_2_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_2_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_2_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_2_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_2_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2456 ? (_GEN_2136 ? (_GEN_2039 ? (_GEN_1655 ? stq_2_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_2_bits_addr_valid <= ~_GEN_5756 & (clear_store ? ~_GEN_5658 & _GEN_2810 : ~_GEN_5210 & _GEN_2810);
    if (_GEN_2809) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_2_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_2_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_2_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_2_bits_addr_bits <= casez_tmp_290;
        else
          stq_2_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_2_bits_addr_bits <= _GEN_280;
      stq_2_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2680) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_2_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_2_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_2_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_2_bits_addr_bits <= casez_tmp_290;
        else
          stq_2_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_2_bits_addr_bits <= _GEN_274;
      stq_2_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_2_bits_data_valid <= ~_GEN_5756 & (clear_store ? ~_GEN_5658 & _GEN_2874 : ~_GEN_5210 & _GEN_2874);
    if (_stq_bits_data_bits_T_2 & _GEN_2873)
      stq_2_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2712)
      stq_2_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_2_bits_committed <= ~_GEN_5718 & (commit_store_3 ? _GEN_5592 | _GEN_5500 | _GEN_5405 : _GEN_5500 | _GEN_5405);
    stq_2_bits_succeeded <= ~_GEN_5718 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h2 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h2 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2585)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2585)) & _GEN_2456 & _GEN_2136 & _GEN_2039 & _GEN_1655 & stq_2_bits_succeeded);
    stq_3_valid <= ~_GEN_5758 & (clear_store ? ~_GEN_5660 & _GEN_2397 : ~_GEN_5211 & _GEN_2397);
    stq_3_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_3_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_3_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_3_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_3_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_3_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_3_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_3_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_3_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_3_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_3_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_3_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_3_bits_uop_taken <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_3_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_3_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_3_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_3_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2457 & _GEN_2137 & _GEN_2040 & _GEN_1656 & stq_3_bits_uop_ppred_busy;
    stq_3_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h3 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h3 | (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_3_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_3_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_3_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_3_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_3_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_3_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_3_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_3_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_3_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_3_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_3_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_3_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_3_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_3_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_3_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_3_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_3_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_3_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_3_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_3_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2457 ? (_GEN_2137 ? (_GEN_2040 ? (_GEN_1656 ? stq_3_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_3_bits_addr_valid <= ~_GEN_5758 & (clear_store ? ~_GEN_5660 & _GEN_2812 : ~_GEN_5211 & _GEN_2812);
    if (_GEN_2811) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_3_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_3_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_3_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_3_bits_addr_bits <= casez_tmp_290;
        else
          stq_3_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_3_bits_addr_bits <= _GEN_280;
      stq_3_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2681) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_3_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_3_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_3_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_3_bits_addr_bits <= casez_tmp_290;
        else
          stq_3_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_3_bits_addr_bits <= _GEN_274;
      stq_3_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_3_bits_data_valid <= ~_GEN_5758 & (clear_store ? ~_GEN_5660 & _GEN_2876 : ~_GEN_5211 & _GEN_2876);
    if (_stq_bits_data_bits_T_2 & _GEN_2875)
      stq_3_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2713)
      stq_3_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_3_bits_committed <= ~_GEN_5719 & (commit_store_3 ? _GEN_5593 | _GEN_5502 | _GEN_5407 : _GEN_5502 | _GEN_5407);
    stq_3_bits_succeeded <= ~_GEN_5719 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h3 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h3 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2586)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2586)) & _GEN_2457 & _GEN_2137 & _GEN_2040 & _GEN_1656 & stq_3_bits_succeeded);
    stq_4_valid <= ~_GEN_5760 & (clear_store ? ~_GEN_5662 & _GEN_2399 : ~_GEN_5212 & _GEN_2399);
    stq_4_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_4_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_4_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_4_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_4_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_4_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_4_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_4_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_4_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_4_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_4_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_4_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_4_bits_uop_taken <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_4_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_4_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_4_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_4_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2458 & _GEN_2138 & _GEN_2041 & _GEN_1657 & stq_4_bits_uop_ppred_busy;
    stq_4_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h4 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h4 | (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_4_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_4_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_4_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_4_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_4_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_4_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_4_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_4_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_4_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_4_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_4_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_4_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_4_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_4_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_4_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_4_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_4_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_4_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_4_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_4_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2458 ? (_GEN_2138 ? (_GEN_2041 ? (_GEN_1657 ? stq_4_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_4_bits_addr_valid <= ~_GEN_5760 & (clear_store ? ~_GEN_5662 & _GEN_2814 : ~_GEN_5212 & _GEN_2814);
    if (_GEN_2813) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_4_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_4_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_4_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_4_bits_addr_bits <= casez_tmp_290;
        else
          stq_4_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_4_bits_addr_bits <= _GEN_280;
      stq_4_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2682) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_4_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_4_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_4_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_4_bits_addr_bits <= casez_tmp_290;
        else
          stq_4_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_4_bits_addr_bits <= _GEN_274;
      stq_4_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_4_bits_data_valid <= ~_GEN_5760 & (clear_store ? ~_GEN_5662 & _GEN_2878 : ~_GEN_5212 & _GEN_2878);
    if (_stq_bits_data_bits_T_2 & _GEN_2877)
      stq_4_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2714)
      stq_4_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_4_bits_committed <= ~_GEN_5720 & (commit_store_3 ? _GEN_5594 | _GEN_5504 | _GEN_5409 : _GEN_5504 | _GEN_5409);
    stq_4_bits_succeeded <= ~_GEN_5720 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h4 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h4 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2587)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2587)) & _GEN_2458 & _GEN_2138 & _GEN_2041 & _GEN_1657 & stq_4_bits_succeeded);
    stq_5_valid <= ~_GEN_5762 & (clear_store ? ~_GEN_5664 & _GEN_2401 : ~_GEN_5213 & _GEN_2401);
    stq_5_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_5_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_5_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_5_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_5_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_5_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_5_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_5_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_5_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_5_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_5_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_5_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_5_bits_uop_taken <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_5_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_5_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_5_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_5_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2459 & _GEN_2139 & _GEN_2042 & _GEN_1658 & stq_5_bits_uop_ppred_busy;
    stq_5_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h5 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h5 | (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_5_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_5_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_5_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_5_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_5_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_5_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_5_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_5_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_5_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_5_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_5_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_5_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_5_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_5_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_5_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_5_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_5_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_5_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_5_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_5_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2459 ? (_GEN_2139 ? (_GEN_2042 ? (_GEN_1658 ? stq_5_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_5_bits_addr_valid <= ~_GEN_5762 & (clear_store ? ~_GEN_5664 & _GEN_2816 : ~_GEN_5213 & _GEN_2816);
    if (_GEN_2815) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_5_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_5_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_5_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_5_bits_addr_bits <= casez_tmp_290;
        else
          stq_5_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_5_bits_addr_bits <= _GEN_280;
      stq_5_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2683) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_5_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_5_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_5_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_5_bits_addr_bits <= casez_tmp_290;
        else
          stq_5_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_5_bits_addr_bits <= _GEN_274;
      stq_5_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_5_bits_data_valid <= ~_GEN_5762 & (clear_store ? ~_GEN_5664 & _GEN_2880 : ~_GEN_5213 & _GEN_2880);
    if (_stq_bits_data_bits_T_2 & _GEN_2879)
      stq_5_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2715)
      stq_5_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_5_bits_committed <= ~_GEN_5721 & (commit_store_3 ? _GEN_5595 | _GEN_5506 | _GEN_5411 : _GEN_5506 | _GEN_5411);
    stq_5_bits_succeeded <= ~_GEN_5721 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h5 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h5 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2588)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2588)) & _GEN_2459 & _GEN_2139 & _GEN_2042 & _GEN_1658 & stq_5_bits_succeeded);
    stq_6_valid <= ~_GEN_5764 & (clear_store ? ~_GEN_5666 & _GEN_2403 : ~_GEN_5214 & _GEN_2403);
    stq_6_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_6_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_6_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_6_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_6_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_6_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_6_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_6_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_6_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_6_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_6_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_6_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_6_bits_uop_taken <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_6_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_6_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_6_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_6_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2460 & _GEN_2140 & _GEN_2043 & _GEN_1659 & stq_6_bits_uop_ppred_busy;
    stq_6_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h6 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h6 | (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_6_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_6_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_6_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_6_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_6_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_6_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_6_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_6_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_6_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_6_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_6_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_6_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_6_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_6_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_6_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_6_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_6_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_6_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_6_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_6_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2460 ? (_GEN_2140 ? (_GEN_2043 ? (_GEN_1659 ? stq_6_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_6_bits_addr_valid <= ~_GEN_5764 & (clear_store ? ~_GEN_5666 & _GEN_2818 : ~_GEN_5214 & _GEN_2818);
    if (_GEN_2817) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_6_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_6_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_6_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_6_bits_addr_bits <= casez_tmp_290;
        else
          stq_6_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_6_bits_addr_bits <= _GEN_280;
      stq_6_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2684) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_6_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_6_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_6_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_6_bits_addr_bits <= casez_tmp_290;
        else
          stq_6_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_6_bits_addr_bits <= _GEN_274;
      stq_6_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_6_bits_data_valid <= ~_GEN_5764 & (clear_store ? ~_GEN_5666 & _GEN_2882 : ~_GEN_5214 & _GEN_2882);
    if (_stq_bits_data_bits_T_2 & _GEN_2881)
      stq_6_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2716)
      stq_6_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_6_bits_committed <= ~_GEN_5722 & (commit_store_3 ? _GEN_5596 | _GEN_5508 | _GEN_5413 : _GEN_5508 | _GEN_5413);
    stq_6_bits_succeeded <= ~_GEN_5722 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h6 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h6 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2589)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2589)) & _GEN_2460 & _GEN_2140 & _GEN_2043 & _GEN_1659 & stq_6_bits_succeeded);
    stq_7_valid <= ~_GEN_5766 & (clear_store ? ~_GEN_5668 & _GEN_2405 : ~_GEN_5215 & _GEN_2405);
    stq_7_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_7_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_7_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_7_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_7_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_7_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_7_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_7_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_7_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_7_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_7_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_7_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_7_bits_uop_taken <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_7_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_7_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_7_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_7_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2461 & _GEN_2141 & _GEN_2044 & _GEN_1660 & stq_7_bits_uop_ppred_busy;
    stq_7_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h7 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h7 | (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_7_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_7_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_7_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_7_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_7_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_7_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_7_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_7_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_7_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_7_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_7_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_7_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_7_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_7_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_7_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_7_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_7_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_7_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_7_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_7_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2461 ? (_GEN_2141 ? (_GEN_2044 ? (_GEN_1660 ? stq_7_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_7_bits_addr_valid <= ~_GEN_5766 & (clear_store ? ~_GEN_5668 & _GEN_2820 : ~_GEN_5215 & _GEN_2820);
    if (_GEN_2819) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_7_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_7_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_7_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_7_bits_addr_bits <= casez_tmp_290;
        else
          stq_7_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_7_bits_addr_bits <= _GEN_280;
      stq_7_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2685) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_7_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_7_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_7_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_7_bits_addr_bits <= casez_tmp_290;
        else
          stq_7_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_7_bits_addr_bits <= _GEN_274;
      stq_7_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_7_bits_data_valid <= ~_GEN_5766 & (clear_store ? ~_GEN_5668 & _GEN_2884 : ~_GEN_5215 & _GEN_2884);
    if (_stq_bits_data_bits_T_2 & _GEN_2883)
      stq_7_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2717)
      stq_7_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_7_bits_committed <= ~_GEN_5723 & (commit_store_3 ? _GEN_5597 | _GEN_5510 | _GEN_5415 : _GEN_5510 | _GEN_5415);
    stq_7_bits_succeeded <= ~_GEN_5723 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h7 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h7 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2590)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2590)) & _GEN_2461 & _GEN_2141 & _GEN_2044 & _GEN_1660 & stq_7_bits_succeeded);
    stq_8_valid <= ~_GEN_5768 & (clear_store ? ~_GEN_5670 & _GEN_2407 : ~_GEN_5216 & _GEN_2407);
    stq_8_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_8_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_8_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_8_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_8_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_8_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_8_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_8_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_8_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_8_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_8_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_8_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_8_bits_uop_taken <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_8_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_8_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_8_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_8_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2462 & _GEN_2142 & _GEN_2045 & _GEN_1661 & stq_8_bits_uop_ppred_busy;
    stq_8_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h8 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h8 | (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_8_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_8_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_8_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_8_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_8_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_8_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_8_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_8_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_8_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_8_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_8_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_8_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_8_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_8_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_8_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_8_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_8_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_8_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_8_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_8_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2462 ? (_GEN_2142 ? (_GEN_2045 ? (_GEN_1661 ? stq_8_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_8_bits_addr_valid <= ~_GEN_5768 & (clear_store ? ~_GEN_5670 & _GEN_2822 : ~_GEN_5216 & _GEN_2822);
    if (_GEN_2821) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_8_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_8_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_8_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_8_bits_addr_bits <= casez_tmp_290;
        else
          stq_8_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_8_bits_addr_bits <= _GEN_280;
      stq_8_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2686) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_8_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_8_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_8_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_8_bits_addr_bits <= casez_tmp_290;
        else
          stq_8_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_8_bits_addr_bits <= _GEN_274;
      stq_8_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_8_bits_data_valid <= ~_GEN_5768 & (clear_store ? ~_GEN_5670 & _GEN_2886 : ~_GEN_5216 & _GEN_2886);
    if (_stq_bits_data_bits_T_2 & _GEN_2885)
      stq_8_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2718)
      stq_8_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_8_bits_committed <= ~_GEN_5724 & (commit_store_3 ? _GEN_5598 | _GEN_5512 | _GEN_5417 : _GEN_5512 | _GEN_5417);
    stq_8_bits_succeeded <= ~_GEN_5724 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h8 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h8 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2591)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2591)) & _GEN_2462 & _GEN_2142 & _GEN_2045 & _GEN_1661 & stq_8_bits_succeeded);
    stq_9_valid <= ~_GEN_5770 & (clear_store ? ~_GEN_5672 & _GEN_2409 : ~_GEN_5217 & _GEN_2409);
    stq_9_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_9_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_9_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_9_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_9_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_9_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_9_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_9_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_9_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_9_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_9_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_9_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_9_bits_uop_taken <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_9_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_9_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_9_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_9_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2463 & _GEN_2143 & _GEN_2046 & _GEN_1662 & stq_9_bits_uop_ppred_busy;
    stq_9_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h9 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h9 | (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_9_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_9_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_9_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_9_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_9_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_9_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_9_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_9_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_9_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_9_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_9_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_9_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_9_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_9_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_9_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_9_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_9_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_9_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_9_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_9_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2463 ? (_GEN_2143 ? (_GEN_2046 ? (_GEN_1662 ? stq_9_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_9_bits_addr_valid <= ~_GEN_5770 & (clear_store ? ~_GEN_5672 & _GEN_2824 : ~_GEN_5217 & _GEN_2824);
    if (_GEN_2823) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_9_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_9_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_9_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_9_bits_addr_bits <= casez_tmp_290;
        else
          stq_9_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_9_bits_addr_bits <= _GEN_280;
      stq_9_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2687) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_9_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_9_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_9_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_9_bits_addr_bits <= casez_tmp_290;
        else
          stq_9_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_9_bits_addr_bits <= _GEN_274;
      stq_9_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_9_bits_data_valid <= ~_GEN_5770 & (clear_store ? ~_GEN_5672 & _GEN_2888 : ~_GEN_5217 & _GEN_2888);
    if (_stq_bits_data_bits_T_2 & _GEN_2887)
      stq_9_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2719)
      stq_9_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_9_bits_committed <= ~_GEN_5725 & (commit_store_3 ? _GEN_5599 | _GEN_5514 | _GEN_5419 : _GEN_5514 | _GEN_5419);
    stq_9_bits_succeeded <= ~_GEN_5725 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h9 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h9 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2592)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2592)) & _GEN_2463 & _GEN_2143 & _GEN_2046 & _GEN_1662 & stq_9_bits_succeeded);
    stq_10_valid <= ~_GEN_5772 & (clear_store ? ~_GEN_5674 & _GEN_2411 : ~_GEN_5218 & _GEN_2411);
    stq_10_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_10_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_10_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_10_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_10_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_10_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_10_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_10_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_10_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_10_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_10_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_10_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_10_bits_uop_taken <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_10_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_10_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_10_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_10_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2464 & _GEN_2144 & _GEN_2047 & _GEN_1663 & stq_10_bits_uop_ppred_busy;
    stq_10_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hA | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hA | (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_10_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_10_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_10_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_10_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_10_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_10_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_10_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_10_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_10_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_10_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_10_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_10_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_10_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_10_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_10_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_10_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_10_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_10_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_10_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_10_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2464 ? (_GEN_2144 ? (_GEN_2047 ? (_GEN_1663 ? stq_10_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_10_bits_addr_valid <= ~_GEN_5772 & (clear_store ? ~_GEN_5674 & _GEN_2826 : ~_GEN_5218 & _GEN_2826);
    if (_GEN_2825) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_10_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_10_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_10_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_10_bits_addr_bits <= casez_tmp_290;
        else
          stq_10_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_10_bits_addr_bits <= _GEN_280;
      stq_10_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2688) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_10_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_10_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_10_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_10_bits_addr_bits <= casez_tmp_290;
        else
          stq_10_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_10_bits_addr_bits <= _GEN_274;
      stq_10_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_10_bits_data_valid <= ~_GEN_5772 & (clear_store ? ~_GEN_5674 & _GEN_2890 : ~_GEN_5218 & _GEN_2890);
    if (_stq_bits_data_bits_T_2 & _GEN_2889)
      stq_10_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2720)
      stq_10_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_10_bits_committed <= ~_GEN_5726 & (commit_store_3 ? _GEN_5600 | _GEN_5516 | _GEN_5421 : _GEN_5516 | _GEN_5421);
    stq_10_bits_succeeded <= ~_GEN_5726 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hA | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hA | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2593)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2593)) & _GEN_2464 & _GEN_2144 & _GEN_2047 & _GEN_1663 & stq_10_bits_succeeded);
    stq_11_valid <= ~_GEN_5774 & (clear_store ? ~_GEN_5676 & _GEN_2413 : ~_GEN_5219 & _GEN_2413);
    stq_11_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_11_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_11_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_11_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_11_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_11_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_11_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_11_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_11_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_11_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_11_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_11_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_11_bits_uop_taken <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_11_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_11_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_11_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_11_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2465 & _GEN_2145 & _GEN_2048 & _GEN_1664 & stq_11_bits_uop_ppred_busy;
    stq_11_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hB | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hB | (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_11_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_11_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_11_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_11_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_11_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_11_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_11_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_11_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_11_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_11_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_11_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_11_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_11_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_11_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_11_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_11_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_11_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_11_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_11_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_11_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2465 ? (_GEN_2145 ? (_GEN_2048 ? (_GEN_1664 ? stq_11_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_11_bits_addr_valid <= ~_GEN_5774 & (clear_store ? ~_GEN_5676 & _GEN_2828 : ~_GEN_5219 & _GEN_2828);
    if (_GEN_2827) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_11_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_11_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_11_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_11_bits_addr_bits <= casez_tmp_290;
        else
          stq_11_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_11_bits_addr_bits <= _GEN_280;
      stq_11_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2689) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_11_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_11_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_11_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_11_bits_addr_bits <= casez_tmp_290;
        else
          stq_11_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_11_bits_addr_bits <= _GEN_274;
      stq_11_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_11_bits_data_valid <= ~_GEN_5774 & (clear_store ? ~_GEN_5676 & _GEN_2892 : ~_GEN_5219 & _GEN_2892);
    if (_stq_bits_data_bits_T_2 & _GEN_2891)
      stq_11_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2721)
      stq_11_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_11_bits_committed <= ~_GEN_5727 & (commit_store_3 ? _GEN_5601 | _GEN_5518 | _GEN_5423 : _GEN_5518 | _GEN_5423);
    stq_11_bits_succeeded <= ~_GEN_5727 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hB | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hB | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2594)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2594)) & _GEN_2465 & _GEN_2145 & _GEN_2048 & _GEN_1664 & stq_11_bits_succeeded);
    stq_12_valid <= ~_GEN_5776 & (clear_store ? ~_GEN_5678 & _GEN_2415 : ~_GEN_5220 & _GEN_2415);
    stq_12_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_12_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_12_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_12_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_12_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_12_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_12_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_12_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_12_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_12_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_12_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_12_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_12_bits_uop_taken <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_12_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_12_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_12_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_12_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2466 & _GEN_2146 & _GEN_2049 & _GEN_1665 & stq_12_bits_uop_ppred_busy;
    stq_12_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hC | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hC | (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_12_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_12_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_12_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_12_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_12_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_12_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_12_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_12_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_12_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_12_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_12_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_12_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_12_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_12_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_12_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_12_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_12_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_12_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_12_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_12_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2466 ? (_GEN_2146 ? (_GEN_2049 ? (_GEN_1665 ? stq_12_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_12_bits_addr_valid <= ~_GEN_5776 & (clear_store ? ~_GEN_5678 & _GEN_2830 : ~_GEN_5220 & _GEN_2830);
    if (_GEN_2829) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_12_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_12_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_12_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_12_bits_addr_bits <= casez_tmp_290;
        else
          stq_12_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_12_bits_addr_bits <= _GEN_280;
      stq_12_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2690) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_12_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_12_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_12_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_12_bits_addr_bits <= casez_tmp_290;
        else
          stq_12_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_12_bits_addr_bits <= _GEN_274;
      stq_12_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_12_bits_data_valid <= ~_GEN_5776 & (clear_store ? ~_GEN_5678 & _GEN_2894 : ~_GEN_5220 & _GEN_2894);
    if (_stq_bits_data_bits_T_2 & _GEN_2893)
      stq_12_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2722)
      stq_12_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_12_bits_committed <= ~_GEN_5728 & (commit_store_3 ? _GEN_5602 | _GEN_5520 | _GEN_5425 : _GEN_5520 | _GEN_5425);
    stq_12_bits_succeeded <= ~_GEN_5728 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hC | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hC | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2595)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2595)) & _GEN_2466 & _GEN_2146 & _GEN_2049 & _GEN_1665 & stq_12_bits_succeeded);
    stq_13_valid <= ~_GEN_5778 & (clear_store ? ~_GEN_5680 & _GEN_2417 : ~_GEN_5221 & _GEN_2417);
    stq_13_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_13_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_13_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_13_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_13_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_13_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_13_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_13_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_13_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_13_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_13_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_13_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_13_bits_uop_taken <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_13_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_13_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_13_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_13_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2467 & _GEN_2147 & _GEN_2050 & _GEN_1666 & stq_13_bits_uop_ppred_busy;
    stq_13_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hD | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hD | (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_13_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_13_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_13_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_13_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_13_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_13_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_13_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_13_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_13_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_13_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_13_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_13_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_13_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_13_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_13_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_13_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_13_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_13_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_13_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_13_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2467 ? (_GEN_2147 ? (_GEN_2050 ? (_GEN_1666 ? stq_13_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_13_bits_addr_valid <= ~_GEN_5778 & (clear_store ? ~_GEN_5680 & _GEN_2832 : ~_GEN_5221 & _GEN_2832);
    if (_GEN_2831) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_13_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_13_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_13_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_13_bits_addr_bits <= casez_tmp_290;
        else
          stq_13_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_13_bits_addr_bits <= _GEN_280;
      stq_13_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2691) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_13_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_13_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_13_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_13_bits_addr_bits <= casez_tmp_290;
        else
          stq_13_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_13_bits_addr_bits <= _GEN_274;
      stq_13_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_13_bits_data_valid <= ~_GEN_5778 & (clear_store ? ~_GEN_5680 & _GEN_2896 : ~_GEN_5221 & _GEN_2896);
    if (_stq_bits_data_bits_T_2 & _GEN_2895)
      stq_13_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2723)
      stq_13_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_13_bits_committed <= ~_GEN_5729 & (commit_store_3 ? _GEN_5603 | _GEN_5522 | _GEN_5427 : _GEN_5522 | _GEN_5427);
    stq_13_bits_succeeded <= ~_GEN_5729 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hD | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hD | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2596)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2596)) & _GEN_2467 & _GEN_2147 & _GEN_2050 & _GEN_1666 & stq_13_bits_succeeded);
    stq_14_valid <= ~_GEN_5780 & (clear_store ? ~_GEN_5682 & _GEN_2419 : ~_GEN_5222 & _GEN_2419);
    stq_14_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_14_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_14_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_14_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_14_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_14_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_14_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_14_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_14_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_14_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_14_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_14_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_14_bits_uop_taken <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_14_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_14_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_14_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_14_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2468 & _GEN_2148 & _GEN_2051 & _GEN_1667 & stq_14_bits_uop_ppred_busy;
    stq_14_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hE | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hE | (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_14_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_14_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_14_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_14_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_14_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_14_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_14_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_14_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_14_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_14_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_14_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_14_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_14_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_14_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_14_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_14_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_14_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_14_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_14_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_14_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2468 ? (_GEN_2148 ? (_GEN_2051 ? (_GEN_1667 ? stq_14_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_14_bits_addr_valid <= ~_GEN_5780 & (clear_store ? ~_GEN_5682 & _GEN_2834 : ~_GEN_5222 & _GEN_2834);
    if (_GEN_2833) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_14_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_14_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_14_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_14_bits_addr_bits <= casez_tmp_290;
        else
          stq_14_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_14_bits_addr_bits <= _GEN_280;
      stq_14_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2692) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_14_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_14_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_14_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_14_bits_addr_bits <= casez_tmp_290;
        else
          stq_14_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_14_bits_addr_bits <= _GEN_274;
      stq_14_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_14_bits_data_valid <= ~_GEN_5780 & (clear_store ? ~_GEN_5682 & _GEN_2898 : ~_GEN_5222 & _GEN_2898);
    if (_stq_bits_data_bits_T_2 & _GEN_2897)
      stq_14_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2724)
      stq_14_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_14_bits_committed <= ~_GEN_5730 & (commit_store_3 ? _GEN_5604 | _GEN_5524 | _GEN_5429 : _GEN_5524 | _GEN_5429);
    stq_14_bits_succeeded <= ~_GEN_5730 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hE | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hE | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2597)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2597)) & _GEN_2468 & _GEN_2148 & _GEN_2051 & _GEN_1667 & stq_14_bits_succeeded);
    stq_15_valid <= ~_GEN_5782 & (clear_store ? ~_GEN_5684 & _GEN_2421 : ~_GEN_5223 & _GEN_2421);
    stq_15_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_15_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_15_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_15_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_15_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_15_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_15_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_15_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_15_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_15_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_15_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_15_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_15_bits_uop_taken <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_15_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_15_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_15_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_15_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2469 & _GEN_2149 & _GEN_2052 & _GEN_1668 & stq_15_bits_uop_ppred_busy;
    stq_15_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hF | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hF | (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_15_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_15_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_15_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_15_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_15_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_15_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_15_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_15_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_15_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_15_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_15_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_15_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_15_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_15_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_15_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_15_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_15_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_15_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_15_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_15_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2469 ? (_GEN_2149 ? (_GEN_2052 ? (_GEN_1668 ? stq_15_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_15_bits_addr_valid <= ~_GEN_5782 & (clear_store ? ~_GEN_5684 & _GEN_2836 : ~_GEN_5223 & _GEN_2836);
    if (_GEN_2835) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_15_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_15_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_15_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_15_bits_addr_bits <= casez_tmp_290;
        else
          stq_15_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_15_bits_addr_bits <= _GEN_280;
      stq_15_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2693) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_15_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_15_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_15_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_15_bits_addr_bits <= casez_tmp_290;
        else
          stq_15_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_15_bits_addr_bits <= _GEN_274;
      stq_15_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_15_bits_data_valid <= ~_GEN_5782 & (clear_store ? ~_GEN_5684 & _GEN_2900 : ~_GEN_5223 & _GEN_2900);
    if (_stq_bits_data_bits_T_2 & _GEN_2899)
      stq_15_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2725)
      stq_15_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_15_bits_committed <= ~_GEN_5731 & (commit_store_3 ? _GEN_5605 | _GEN_5526 | _GEN_5431 : _GEN_5526 | _GEN_5431);
    stq_15_bits_succeeded <= ~_GEN_5731 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hF | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hF | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2598)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2598)) & _GEN_2469 & _GEN_2149 & _GEN_2052 & _GEN_1668 & stq_15_bits_succeeded);
    stq_16_valid <= ~_GEN_5784 & (clear_store ? ~_GEN_5686 & _GEN_2423 : ~_GEN_5224 & _GEN_2423);
    stq_16_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_16_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_16_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_16_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_16_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_16_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_16_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_16_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_16_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_16_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_16_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_16_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_16_bits_uop_taken <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_16_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_16_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_16_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_16_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2470 & _GEN_2150 & _GEN_2053 & _GEN_1669 & stq_16_bits_uop_ppred_busy;
    stq_16_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h10 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h10 | (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_16_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_16_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_16_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_16_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_16_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_16_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_16_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_16_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_16_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_16_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_16_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_16_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_16_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_16_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_16_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_16_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_16_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_16_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_16_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_16_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2470 ? (_GEN_2150 ? (_GEN_2053 ? (_GEN_1669 ? stq_16_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_16_bits_addr_valid <= ~_GEN_5784 & (clear_store ? ~_GEN_5686 & _GEN_2838 : ~_GEN_5224 & _GEN_2838);
    if (_GEN_2837) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_16_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_16_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_16_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_16_bits_addr_bits <= casez_tmp_290;
        else
          stq_16_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_16_bits_addr_bits <= _GEN_280;
      stq_16_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2694) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_16_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_16_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_16_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_16_bits_addr_bits <= casez_tmp_290;
        else
          stq_16_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_16_bits_addr_bits <= _GEN_274;
      stq_16_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_16_bits_data_valid <= ~_GEN_5784 & (clear_store ? ~_GEN_5686 & _GEN_2902 : ~_GEN_5224 & _GEN_2902);
    if (_stq_bits_data_bits_T_2 & _GEN_2901)
      stq_16_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2726)
      stq_16_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_16_bits_committed <= ~_GEN_5732 & (commit_store_3 ? _GEN_5606 | _GEN_5528 | _GEN_5433 : _GEN_5528 | _GEN_5433);
    stq_16_bits_succeeded <= ~_GEN_5732 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h10 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h10 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2599)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2599)) & _GEN_2470 & _GEN_2150 & _GEN_2053 & _GEN_1669 & stq_16_bits_succeeded);
    stq_17_valid <= ~_GEN_5786 & (clear_store ? ~_GEN_5688 & _GEN_2425 : ~_GEN_5225 & _GEN_2425);
    stq_17_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_17_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_17_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_17_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_17_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_17_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_17_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_17_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_17_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_17_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_17_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_17_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_17_bits_uop_taken <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_17_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_17_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_17_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_17_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2471 & _GEN_2151 & _GEN_2054 & _GEN_1670 & stq_17_bits_uop_ppred_busy;
    stq_17_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h11 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h11 | (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_17_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_17_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_17_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_17_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_17_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_17_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_17_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_17_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_17_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_17_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_17_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_17_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_17_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_17_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_17_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_17_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_17_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_17_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_17_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_17_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2471 ? (_GEN_2151 ? (_GEN_2054 ? (_GEN_1670 ? stq_17_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_17_bits_addr_valid <= ~_GEN_5786 & (clear_store ? ~_GEN_5688 & _GEN_2840 : ~_GEN_5225 & _GEN_2840);
    if (_GEN_2839) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_17_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_17_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_17_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_17_bits_addr_bits <= casez_tmp_290;
        else
          stq_17_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_17_bits_addr_bits <= _GEN_280;
      stq_17_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2695) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_17_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_17_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_17_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_17_bits_addr_bits <= casez_tmp_290;
        else
          stq_17_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_17_bits_addr_bits <= _GEN_274;
      stq_17_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_17_bits_data_valid <= ~_GEN_5786 & (clear_store ? ~_GEN_5688 & _GEN_2904 : ~_GEN_5225 & _GEN_2904);
    if (_stq_bits_data_bits_T_2 & _GEN_2903)
      stq_17_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2727)
      stq_17_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_17_bits_committed <= ~_GEN_5733 & (commit_store_3 ? _GEN_5607 | _GEN_5530 | _GEN_5435 : _GEN_5530 | _GEN_5435);
    stq_17_bits_succeeded <= ~_GEN_5733 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h11 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h11 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2600)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2600)) & _GEN_2471 & _GEN_2151 & _GEN_2054 & _GEN_1670 & stq_17_bits_succeeded);
    stq_18_valid <= ~_GEN_5788 & (clear_store ? ~_GEN_5690 & _GEN_2427 : ~_GEN_5226 & _GEN_2427);
    stq_18_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_18_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_18_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_18_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_18_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_18_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_18_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_18_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_18_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_18_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_18_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_18_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_18_bits_uop_taken <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_18_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_18_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_18_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_18_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2472 & _GEN_2152 & _GEN_2055 & _GEN_1671 & stq_18_bits_uop_ppred_busy;
    stq_18_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h12 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h12 | (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_18_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_18_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_18_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_18_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_18_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_18_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_18_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_18_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_18_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_18_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_18_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_18_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_18_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_18_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_18_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_18_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_18_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_18_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_18_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_18_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2472 ? (_GEN_2152 ? (_GEN_2055 ? (_GEN_1671 ? stq_18_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_18_bits_addr_valid <= ~_GEN_5788 & (clear_store ? ~_GEN_5690 & _GEN_2842 : ~_GEN_5226 & _GEN_2842);
    if (_GEN_2841) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_18_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_18_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_18_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_18_bits_addr_bits <= casez_tmp_290;
        else
          stq_18_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_18_bits_addr_bits <= _GEN_280;
      stq_18_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2696) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_18_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_18_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_18_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_18_bits_addr_bits <= casez_tmp_290;
        else
          stq_18_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_18_bits_addr_bits <= _GEN_274;
      stq_18_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_18_bits_data_valid <= ~_GEN_5788 & (clear_store ? ~_GEN_5690 & _GEN_2906 : ~_GEN_5226 & _GEN_2906);
    if (_stq_bits_data_bits_T_2 & _GEN_2905)
      stq_18_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2728)
      stq_18_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_18_bits_committed <= ~_GEN_5734 & (commit_store_3 ? _GEN_5608 | _GEN_5532 | _GEN_5437 : _GEN_5532 | _GEN_5437);
    stq_18_bits_succeeded <= ~_GEN_5734 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h12 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h12 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2601)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2601)) & _GEN_2472 & _GEN_2152 & _GEN_2055 & _GEN_1671 & stq_18_bits_succeeded);
    stq_19_valid <= ~_GEN_5790 & (clear_store ? ~_GEN_5692 & _GEN_2429 : ~_GEN_5227 & _GEN_2429);
    stq_19_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_19_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_19_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_19_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_19_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_19_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_19_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_19_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_19_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_19_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_19_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_19_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_19_bits_uop_taken <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_19_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_19_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_19_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_19_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2473 & _GEN_2153 & _GEN_2056 & _GEN_1672 & stq_19_bits_uop_ppred_busy;
    stq_19_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h13 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h13 | (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_19_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_19_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_19_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_19_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_19_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_19_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_19_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_19_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_19_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_19_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_19_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_19_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_19_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_19_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_19_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_19_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_19_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_19_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_19_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_19_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2473 ? (_GEN_2153 ? (_GEN_2056 ? (_GEN_1672 ? stq_19_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_19_bits_addr_valid <= ~_GEN_5790 & (clear_store ? ~_GEN_5692 & _GEN_2844 : ~_GEN_5227 & _GEN_2844);
    if (_GEN_2843) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_19_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_19_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_19_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_19_bits_addr_bits <= casez_tmp_290;
        else
          stq_19_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_19_bits_addr_bits <= _GEN_280;
      stq_19_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2697) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_19_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_19_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_19_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_19_bits_addr_bits <= casez_tmp_290;
        else
          stq_19_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_19_bits_addr_bits <= _GEN_274;
      stq_19_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_19_bits_data_valid <= ~_GEN_5790 & (clear_store ? ~_GEN_5692 & _GEN_2908 : ~_GEN_5227 & _GEN_2908);
    if (_stq_bits_data_bits_T_2 & _GEN_2907)
      stq_19_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2729)
      stq_19_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_19_bits_committed <= ~_GEN_5735 & (commit_store_3 ? _GEN_5609 | _GEN_5534 | _GEN_5439 : _GEN_5534 | _GEN_5439);
    stq_19_bits_succeeded <= ~_GEN_5735 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h13 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h13 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2602)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2602)) & _GEN_2473 & _GEN_2153 & _GEN_2056 & _GEN_1672 & stq_19_bits_succeeded);
    stq_20_valid <= ~_GEN_5792 & (clear_store ? ~_GEN_5694 & _GEN_2431 : ~_GEN_5228 & _GEN_2431);
    stq_20_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_20_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_20_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_20_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_20_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_20_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_20_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_20_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_20_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_20_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_20_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_20_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_20_bits_uop_taken <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_20_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_20_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_20_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_20_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2474 & _GEN_2154 & _GEN_2057 & _GEN_1673 & stq_20_bits_uop_ppred_busy;
    stq_20_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h14 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h14 | (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_20_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_20_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_20_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_20_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_20_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_20_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_20_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_20_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_20_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_20_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_20_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_20_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_20_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_20_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_20_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_20_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_20_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_20_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_20_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_20_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2474 ? (_GEN_2154 ? (_GEN_2057 ? (_GEN_1673 ? stq_20_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_20_bits_addr_valid <= ~_GEN_5792 & (clear_store ? ~_GEN_5694 & _GEN_2846 : ~_GEN_5228 & _GEN_2846);
    if (_GEN_2845) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_20_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_20_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_20_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_20_bits_addr_bits <= casez_tmp_290;
        else
          stq_20_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_20_bits_addr_bits <= _GEN_280;
      stq_20_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2698) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_20_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_20_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_20_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_20_bits_addr_bits <= casez_tmp_290;
        else
          stq_20_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_20_bits_addr_bits <= _GEN_274;
      stq_20_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_20_bits_data_valid <= ~_GEN_5792 & (clear_store ? ~_GEN_5694 & _GEN_2910 : ~_GEN_5228 & _GEN_2910);
    if (_stq_bits_data_bits_T_2 & _GEN_2909)
      stq_20_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2730)
      stq_20_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_20_bits_committed <= ~_GEN_5736 & (commit_store_3 ? _GEN_5610 | _GEN_5536 | _GEN_5441 : _GEN_5536 | _GEN_5441);
    stq_20_bits_succeeded <= ~_GEN_5736 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h14 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h14 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2603)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2603)) & _GEN_2474 & _GEN_2154 & _GEN_2057 & _GEN_1673 & stq_20_bits_succeeded);
    stq_21_valid <= ~_GEN_5794 & (clear_store ? ~_GEN_5696 & _GEN_2433 : ~_GEN_5229 & _GEN_2433);
    stq_21_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_21_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_21_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_21_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_21_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_21_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_21_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_21_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_21_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_21_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_21_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_21_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_21_bits_uop_taken <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_21_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_21_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_21_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_21_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2475 & _GEN_2155 & _GEN_2058 & _GEN_1674 & stq_21_bits_uop_ppred_busy;
    stq_21_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h15 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h15 | (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_21_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_21_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_21_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_21_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_21_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_21_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_21_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_21_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_21_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_21_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_21_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_21_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_21_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_21_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_21_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_21_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_21_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_21_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_21_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_21_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2475 ? (_GEN_2155 ? (_GEN_2058 ? (_GEN_1674 ? stq_21_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_21_bits_addr_valid <= ~_GEN_5794 & (clear_store ? ~_GEN_5696 & _GEN_2848 : ~_GEN_5229 & _GEN_2848);
    if (_GEN_2847) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_21_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_21_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_21_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_21_bits_addr_bits <= casez_tmp_290;
        else
          stq_21_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_21_bits_addr_bits <= _GEN_280;
      stq_21_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2699) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_21_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_21_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_21_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_21_bits_addr_bits <= casez_tmp_290;
        else
          stq_21_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_21_bits_addr_bits <= _GEN_274;
      stq_21_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_21_bits_data_valid <= ~_GEN_5794 & (clear_store ? ~_GEN_5696 & _GEN_2912 : ~_GEN_5229 & _GEN_2912);
    if (_stq_bits_data_bits_T_2 & _GEN_2911)
      stq_21_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2731)
      stq_21_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_21_bits_committed <= ~_GEN_5737 & (commit_store_3 ? _GEN_5611 | _GEN_5538 | _GEN_5443 : _GEN_5538 | _GEN_5443);
    stq_21_bits_succeeded <= ~_GEN_5737 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h15 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h15 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2604)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2604)) & _GEN_2475 & _GEN_2155 & _GEN_2058 & _GEN_1674 & stq_21_bits_succeeded);
    stq_22_valid <= ~_GEN_5796 & (clear_store ? ~_GEN_5698 & _GEN_2435 : ~_GEN_5230 & _GEN_2435);
    stq_22_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_22_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_22_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_22_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_22_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_22_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_22_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_22_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_22_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_22_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_22_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_22_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_22_bits_uop_taken <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_22_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_22_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_22_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_22_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2476 & _GEN_2156 & _GEN_2059 & _GEN_1675 & stq_22_bits_uop_ppred_busy;
    stq_22_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h16 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h16 | (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_22_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_22_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_22_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_22_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_22_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_22_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_22_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_22_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_22_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_22_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_22_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_22_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_22_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_22_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_22_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_22_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_22_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_22_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_22_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_22_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2476 ? (_GEN_2156 ? (_GEN_2059 ? (_GEN_1675 ? stq_22_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_22_bits_addr_valid <= ~_GEN_5796 & (clear_store ? ~_GEN_5698 & _GEN_2850 : ~_GEN_5230 & _GEN_2850);
    if (_GEN_2849) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_22_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_22_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_22_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_22_bits_addr_bits <= casez_tmp_290;
        else
          stq_22_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_22_bits_addr_bits <= _GEN_280;
      stq_22_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2700) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_22_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_22_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_22_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_22_bits_addr_bits <= casez_tmp_290;
        else
          stq_22_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_22_bits_addr_bits <= _GEN_274;
      stq_22_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_22_bits_data_valid <= ~_GEN_5796 & (clear_store ? ~_GEN_5698 & _GEN_2914 : ~_GEN_5230 & _GEN_2914);
    if (_stq_bits_data_bits_T_2 & _GEN_2913)
      stq_22_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2732)
      stq_22_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_22_bits_committed <= ~_GEN_5738 & (commit_store_3 ? _GEN_5612 | _GEN_5540 | _GEN_5445 : _GEN_5540 | _GEN_5445);
    stq_22_bits_succeeded <= ~_GEN_5738 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h16 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h16 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2605)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2605)) & _GEN_2476 & _GEN_2156 & _GEN_2059 & _GEN_1675 & stq_22_bits_succeeded);
    stq_23_valid <= ~_GEN_5798 & (clear_store ? ~_GEN_5700 & _GEN_2437 : ~_GEN_5231 & _GEN_2437);
    stq_23_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_23_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_23_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_23_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_23_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_23_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_23_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_23_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_23_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_23_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_23_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_23_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_23_bits_uop_taken <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_23_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_23_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_23_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_23_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2477 & _GEN_2157 & _GEN_2060 & _GEN_1676 & stq_23_bits_uop_ppred_busy;
    stq_23_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h17 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h17 | (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_23_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_23_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_23_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_23_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_23_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_23_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_23_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_23_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_23_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_23_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_23_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_23_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_23_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_23_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_23_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_23_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_23_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_23_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_23_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_23_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2477 ? (_GEN_2157 ? (_GEN_2060 ? (_GEN_1676 ? stq_23_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_23_bits_addr_valid <= ~_GEN_5798 & (clear_store ? ~_GEN_5700 & _GEN_2852 : ~_GEN_5231 & _GEN_2852);
    if (_GEN_2851) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_23_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_23_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_23_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_23_bits_addr_bits <= casez_tmp_290;
        else
          stq_23_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_23_bits_addr_bits <= _GEN_280;
      stq_23_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2701) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_23_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_23_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_23_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_23_bits_addr_bits <= casez_tmp_290;
        else
          stq_23_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_23_bits_addr_bits <= _GEN_274;
      stq_23_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_23_bits_data_valid <= ~_GEN_5798 & (clear_store ? ~_GEN_5700 & _GEN_2916 : ~_GEN_5231 & _GEN_2916);
    if (_stq_bits_data_bits_T_2 & _GEN_2915)
      stq_23_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2733)
      stq_23_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_23_bits_committed <= ~_GEN_5739 & (commit_store_3 ? _GEN_5613 | _GEN_5542 | _GEN_5447 : _GEN_5542 | _GEN_5447);
    stq_23_bits_succeeded <= ~_GEN_5739 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h17 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h17 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2606)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2606)) & _GEN_2477 & _GEN_2157 & _GEN_2060 & _GEN_1676 & stq_23_bits_succeeded);
    stq_24_valid <= ~_GEN_5800 & (clear_store ? ~_GEN_5702 & _GEN_2439 : ~_GEN_5232 & _GEN_2439);
    stq_24_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_24_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_24_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_24_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_24_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_24_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_24_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_24_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_24_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_24_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_24_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_24_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_24_bits_uop_taken <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_24_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_24_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_24_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_24_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2478 & _GEN_2158 & _GEN_2061 & _GEN_1677 & stq_24_bits_uop_ppred_busy;
    stq_24_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h18 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h18 | (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_24_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_24_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_24_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_24_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_24_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_24_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_24_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_24_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_24_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_24_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_24_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_24_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_24_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_24_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_24_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_24_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_24_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_24_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_24_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_24_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2478 ? (_GEN_2158 ? (_GEN_2061 ? (_GEN_1677 ? stq_24_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_24_bits_addr_valid <= ~_GEN_5800 & (clear_store ? ~_GEN_5702 & _GEN_2854 : ~_GEN_5232 & _GEN_2854);
    if (_GEN_2853) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_24_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_24_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_24_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_24_bits_addr_bits <= casez_tmp_290;
        else
          stq_24_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_24_bits_addr_bits <= _GEN_280;
      stq_24_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2702) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_24_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_24_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_24_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_24_bits_addr_bits <= casez_tmp_290;
        else
          stq_24_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_24_bits_addr_bits <= _GEN_274;
      stq_24_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_24_bits_data_valid <= ~_GEN_5800 & (clear_store ? ~_GEN_5702 & _GEN_2918 : ~_GEN_5232 & _GEN_2918);
    if (_stq_bits_data_bits_T_2 & _GEN_2917)
      stq_24_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2734)
      stq_24_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_24_bits_committed <= ~_GEN_5740 & (commit_store_3 ? _GEN_5614 | _GEN_5544 | _GEN_5449 : _GEN_5544 | _GEN_5449);
    stq_24_bits_succeeded <= ~_GEN_5740 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h18 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h18 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2607)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2607)) & _GEN_2478 & _GEN_2158 & _GEN_2061 & _GEN_1677 & stq_24_bits_succeeded);
    stq_25_valid <= ~_GEN_5802 & (clear_store ? ~_GEN_5704 & _GEN_2441 : ~_GEN_5233 & _GEN_2441);
    stq_25_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_25_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_25_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_25_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_25_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_25_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_25_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_25_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_25_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_25_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_25_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_25_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_25_bits_uop_taken <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_25_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_25_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_25_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_25_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2479 & _GEN_2159 & _GEN_2062 & _GEN_1678 & stq_25_bits_uop_ppred_busy;
    stq_25_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h19 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h19 | (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_25_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_25_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_25_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_25_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_25_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_25_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_25_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_25_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_25_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_25_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_25_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_25_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_25_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_25_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_25_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_25_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_25_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_25_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_25_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_25_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2479 ? (_GEN_2159 ? (_GEN_2062 ? (_GEN_1678 ? stq_25_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_25_bits_addr_valid <= ~_GEN_5802 & (clear_store ? ~_GEN_5704 & _GEN_2856 : ~_GEN_5233 & _GEN_2856);
    if (_GEN_2855) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_25_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_25_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_25_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_25_bits_addr_bits <= casez_tmp_290;
        else
          stq_25_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_25_bits_addr_bits <= _GEN_280;
      stq_25_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2703) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_25_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_25_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_25_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_25_bits_addr_bits <= casez_tmp_290;
        else
          stq_25_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_25_bits_addr_bits <= _GEN_274;
      stq_25_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_25_bits_data_valid <= ~_GEN_5802 & (clear_store ? ~_GEN_5704 & _GEN_2920 : ~_GEN_5233 & _GEN_2920);
    if (_stq_bits_data_bits_T_2 & _GEN_2919)
      stq_25_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2735)
      stq_25_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_25_bits_committed <= ~_GEN_5741 & (commit_store_3 ? _GEN_5615 | _GEN_5546 | _GEN_5451 : _GEN_5546 | _GEN_5451);
    stq_25_bits_succeeded <= ~_GEN_5741 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h19 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h19 | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2608)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2608)) & _GEN_2479 & _GEN_2159 & _GEN_2062 & _GEN_1678 & stq_25_bits_succeeded);
    stq_26_valid <= ~_GEN_5804 & (clear_store ? ~_GEN_5706 & _GEN_2443 : ~_GEN_5234 & _GEN_2443);
    stq_26_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_26_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_26_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_26_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_26_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_26_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_26_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_26_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_26_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_26_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_26_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_26_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_26_bits_uop_taken <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_26_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_26_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_26_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_26_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2480 & _GEN_2160 & _GEN_2063 & _GEN_1679 & stq_26_bits_uop_ppred_busy;
    stq_26_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1A | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1A | (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_26_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_26_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_26_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_26_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_26_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_26_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_26_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_26_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_26_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_26_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_26_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_26_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_26_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_26_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_26_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_26_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_26_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_26_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_26_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_26_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2480 ? (_GEN_2160 ? (_GEN_2063 ? (_GEN_1679 ? stq_26_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_26_bits_addr_valid <= ~_GEN_5804 & (clear_store ? ~_GEN_5706 & _GEN_2858 : ~_GEN_5234 & _GEN_2858);
    if (_GEN_2857) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_26_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_26_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_26_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_26_bits_addr_bits <= casez_tmp_290;
        else
          stq_26_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_26_bits_addr_bits <= _GEN_280;
      stq_26_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2704) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_26_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_26_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_26_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_26_bits_addr_bits <= casez_tmp_290;
        else
          stq_26_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_26_bits_addr_bits <= _GEN_274;
      stq_26_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_26_bits_data_valid <= ~_GEN_5804 & (clear_store ? ~_GEN_5706 & _GEN_2922 : ~_GEN_5234 & _GEN_2922);
    if (_stq_bits_data_bits_T_2 & _GEN_2921)
      stq_26_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2736)
      stq_26_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_26_bits_committed <= ~_GEN_5742 & (commit_store_3 ? _GEN_5616 | _GEN_5548 | _GEN_5453 : _GEN_5548 | _GEN_5453);
    stq_26_bits_succeeded <= ~_GEN_5742 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1A | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1A | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2609)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2609)) & _GEN_2480 & _GEN_2160 & _GEN_2063 & _GEN_1679 & stq_26_bits_succeeded);
    stq_27_valid <= ~_GEN_5806 & (clear_store ? ~_GEN_5708 & _GEN_2445 : ~_GEN_5235 & _GEN_2445);
    stq_27_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_27_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_27_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_27_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_27_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_27_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_27_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_27_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_27_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_27_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_27_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_27_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_27_bits_uop_taken <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_27_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_27_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_27_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_27_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2481 & _GEN_2161 & _GEN_2064 & _GEN_1680 & stq_27_bits_uop_ppred_busy;
    stq_27_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1B | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1B | (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_27_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_27_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_27_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_27_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_27_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_27_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_27_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_27_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_27_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_27_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_27_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_27_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_27_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_27_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_27_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_27_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_27_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_27_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_27_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_27_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2481 ? (_GEN_2161 ? (_GEN_2064 ? (_GEN_1680 ? stq_27_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_27_bits_addr_valid <= ~_GEN_5806 & (clear_store ? ~_GEN_5708 & _GEN_2860 : ~_GEN_5235 & _GEN_2860);
    if (_GEN_2859) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_27_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_27_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_27_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_27_bits_addr_bits <= casez_tmp_290;
        else
          stq_27_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_27_bits_addr_bits <= _GEN_280;
      stq_27_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2705) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_27_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_27_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_27_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_27_bits_addr_bits <= casez_tmp_290;
        else
          stq_27_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_27_bits_addr_bits <= _GEN_274;
      stq_27_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_27_bits_data_valid <= ~_GEN_5806 & (clear_store ? ~_GEN_5708 & _GEN_2924 : ~_GEN_5235 & _GEN_2924);
    if (_stq_bits_data_bits_T_2 & _GEN_2923)
      stq_27_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2737)
      stq_27_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_27_bits_committed <= ~_GEN_5743 & (commit_store_3 ? _GEN_5617 | _GEN_5550 | _GEN_5455 : _GEN_5550 | _GEN_5455);
    stq_27_bits_succeeded <= ~_GEN_5743 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1B | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1B | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2610)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2610)) & _GEN_2481 & _GEN_2161 & _GEN_2064 & _GEN_1680 & stq_27_bits_succeeded);
    stq_28_valid <= ~_GEN_5808 & (clear_store ? ~_GEN_5710 & _GEN_2447 : ~_GEN_5236 & _GEN_2447);
    stq_28_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_28_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_28_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_28_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_28_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_28_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_28_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_28_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_28_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_28_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_28_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_28_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_28_bits_uop_taken <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_28_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_28_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_28_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_28_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2482 & _GEN_2162 & _GEN_2065 & _GEN_1681 & stq_28_bits_uop_ppred_busy;
    stq_28_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1C | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1C | (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_28_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_28_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_28_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_28_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_28_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_28_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_28_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_28_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_28_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_28_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_28_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_28_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_28_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_28_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_28_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_28_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_28_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_28_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_28_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_28_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2482 ? (_GEN_2162 ? (_GEN_2065 ? (_GEN_1681 ? stq_28_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_28_bits_addr_valid <= ~_GEN_5808 & (clear_store ? ~_GEN_5710 & _GEN_2862 : ~_GEN_5236 & _GEN_2862);
    if (_GEN_2861) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_28_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_28_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_28_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_28_bits_addr_bits <= casez_tmp_290;
        else
          stq_28_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_28_bits_addr_bits <= _GEN_280;
      stq_28_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2706) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_28_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_28_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_28_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_28_bits_addr_bits <= casez_tmp_290;
        else
          stq_28_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_28_bits_addr_bits <= _GEN_274;
      stq_28_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_28_bits_data_valid <= ~_GEN_5808 & (clear_store ? ~_GEN_5710 & _GEN_2926 : ~_GEN_5236 & _GEN_2926);
    if (_stq_bits_data_bits_T_2 & _GEN_2925)
      stq_28_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2738)
      stq_28_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_28_bits_committed <= ~_GEN_5744 & (commit_store_3 ? _GEN_5618 | _GEN_5552 | _GEN_5457 : _GEN_5552 | _GEN_5457);
    stq_28_bits_succeeded <= ~_GEN_5744 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1C | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1C | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2611)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2611)) & _GEN_2482 & _GEN_2162 & _GEN_2065 & _GEN_1681 & stq_28_bits_succeeded);
    stq_29_valid <= ~_GEN_5810 & (clear_store ? ~_GEN_5712 & _GEN_2449 : ~_GEN_5237 & _GEN_2449);
    stq_29_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_29_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_29_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_29_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_29_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_29_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_29_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_29_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_29_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_29_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_29_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_29_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_29_bits_uop_taken <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_29_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_29_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_29_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_29_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2483 & _GEN_2163 & _GEN_2066 & _GEN_1682 & stq_29_bits_uop_ppred_busy;
    stq_29_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1D | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1D | (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_29_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_29_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_29_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_29_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_29_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_29_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_29_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_29_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_29_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_29_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_29_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_29_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_29_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_29_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_29_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_29_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_29_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_29_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_29_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_29_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2483 ? (_GEN_2163 ? (_GEN_2066 ? (_GEN_1682 ? stq_29_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_29_bits_addr_valid <= ~_GEN_5810 & (clear_store ? ~_GEN_5712 & _GEN_2864 : ~_GEN_5237 & _GEN_2864);
    if (_GEN_2863) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_29_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_29_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_29_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_29_bits_addr_bits <= casez_tmp_290;
        else
          stq_29_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_29_bits_addr_bits <= _GEN_280;
      stq_29_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2707) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_29_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_29_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_29_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_29_bits_addr_bits <= casez_tmp_290;
        else
          stq_29_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_29_bits_addr_bits <= _GEN_274;
      stq_29_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_29_bits_data_valid <= ~_GEN_5810 & (clear_store ? ~_GEN_5712 & _GEN_2928 : ~_GEN_5237 & _GEN_2928);
    if (_stq_bits_data_bits_T_2 & _GEN_2927)
      stq_29_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2739)
      stq_29_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_29_bits_committed <= ~_GEN_5745 & (commit_store_3 ? _GEN_5619 | _GEN_5554 | _GEN_5459 : _GEN_5554 | _GEN_5459);
    stq_29_bits_succeeded <= ~_GEN_5745 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1D | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1D | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2612)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2612)) & _GEN_2483 & _GEN_2163 & _GEN_2066 & _GEN_1682 & stq_29_bits_succeeded);
    stq_30_valid <= ~_GEN_5812 & (clear_store ? ~_GEN_5714 & _GEN_2451 : ~_GEN_5238 & _GEN_2451);
    stq_30_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_30_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_30_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_30_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_30_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_30_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_30_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_30_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_30_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_30_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_30_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_30_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_30_bits_uop_taken <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_30_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_30_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_30_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_30_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2484 & _GEN_2164 & _GEN_2067 & _GEN_1683 & stq_30_bits_uop_ppred_busy;
    stq_30_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1E | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1E | (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_30_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_30_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_30_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_30_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_30_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_30_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_30_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_30_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_30_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_30_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_30_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_30_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_30_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_30_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_30_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_30_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_30_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_30_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_30_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_30_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2484 ? (_GEN_2164 ? (_GEN_2067 ? (_GEN_1683 ? stq_30_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_30_bits_addr_valid <= ~_GEN_5812 & (clear_store ? ~_GEN_5714 & _GEN_2866 : ~_GEN_5238 & _GEN_2866);
    if (_GEN_2865) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_30_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_30_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_30_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_30_bits_addr_bits <= casez_tmp_290;
        else
          stq_30_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_30_bits_addr_bits <= _GEN_280;
      stq_30_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2708) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_30_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_30_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_30_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_30_bits_addr_bits <= casez_tmp_290;
        else
          stq_30_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_30_bits_addr_bits <= _GEN_274;
      stq_30_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_30_bits_data_valid <= ~_GEN_5812 & (clear_store ? ~_GEN_5714 & _GEN_2930 : ~_GEN_5238 & _GEN_2930);
    if (_stq_bits_data_bits_T_2 & _GEN_2929)
      stq_30_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2740)
      stq_30_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_30_bits_committed <= ~_GEN_5746 & (commit_store_3 ? _GEN_5620 | _GEN_5556 | _GEN_5461 : _GEN_5556 | _GEN_5461);
    stq_30_bits_succeeded <= ~_GEN_5746 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1E | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1E | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & _GEN_2613)) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & _GEN_2613)) & _GEN_2484 & _GEN_2164 & _GEN_2067 & _GEN_1683 & stq_30_bits_succeeded);
    stq_31_valid <= ~_GEN_5814 & (clear_store ? ~_GEN_5715 & _GEN_2453 : ~_GEN_5239 & _GEN_2453);
    stq_31_bits_uop_is_rvc <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_rvc : io_core_dis_uops_0_bits_is_rvc) : io_core_dis_uops_1_bits_is_rvc) : io_core_dis_uops_2_bits_is_rvc) : io_core_dis_uops_3_bits_is_rvc);
    stq_31_bits_uop_ctrl_fcn_dw <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_ctrl_fcn_dw : io_core_dis_uops_0_bits_ctrl_fcn_dw) : io_core_dis_uops_1_bits_ctrl_fcn_dw) : io_core_dis_uops_2_bits_ctrl_fcn_dw) : io_core_dis_uops_3_bits_ctrl_fcn_dw);
    stq_31_bits_uop_ctrl_is_load <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_31_bits_uop_ctrl_is_sta <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_31_bits_uop_ctrl_is_std <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_ctrl_is_std : io_core_dis_uops_0_bits_ctrl_is_std) : io_core_dis_uops_1_bits_ctrl_is_std) : io_core_dis_uops_2_bits_ctrl_is_std) : io_core_dis_uops_3_bits_ctrl_is_std);
    stq_31_bits_uop_iw_p1_poisoned <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_iw_p1_poisoned : io_core_dis_uops_0_bits_iw_p1_poisoned) : io_core_dis_uops_1_bits_iw_p1_poisoned) : io_core_dis_uops_2_bits_iw_p1_poisoned) : io_core_dis_uops_3_bits_iw_p1_poisoned);
    stq_31_bits_uop_iw_p2_poisoned <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_iw_p2_poisoned : io_core_dis_uops_0_bits_iw_p2_poisoned) : io_core_dis_uops_1_bits_iw_p2_poisoned) : io_core_dis_uops_2_bits_iw_p2_poisoned) : io_core_dis_uops_3_bits_iw_p2_poisoned);
    stq_31_bits_uop_is_br <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_br : io_core_dis_uops_0_bits_is_br) : io_core_dis_uops_1_bits_is_br) : io_core_dis_uops_2_bits_is_br) : io_core_dis_uops_3_bits_is_br);
    stq_31_bits_uop_is_jalr <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_jalr : io_core_dis_uops_0_bits_is_jalr) : io_core_dis_uops_1_bits_is_jalr) : io_core_dis_uops_2_bits_is_jalr) : io_core_dis_uops_3_bits_is_jalr);
    stq_31_bits_uop_is_jal <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_jal : io_core_dis_uops_0_bits_is_jal) : io_core_dis_uops_1_bits_is_jal) : io_core_dis_uops_2_bits_is_jal) : io_core_dis_uops_3_bits_is_jal);
    stq_31_bits_uop_is_sfb <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_sfb : io_core_dis_uops_0_bits_is_sfb) : io_core_dis_uops_1_bits_is_sfb) : io_core_dis_uops_2_bits_is_sfb) : io_core_dis_uops_3_bits_is_sfb);
    stq_31_bits_uop_edge_inst <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_edge_inst : io_core_dis_uops_0_bits_edge_inst) : io_core_dis_uops_1_bits_edge_inst) : io_core_dis_uops_2_bits_edge_inst) : io_core_dis_uops_3_bits_edge_inst);
    stq_31_bits_uop_taken <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_taken : io_core_dis_uops_0_bits_taken) : io_core_dis_uops_1_bits_taken) : io_core_dis_uops_2_bits_taken) : io_core_dis_uops_3_bits_taken);
    stq_31_bits_uop_prs1_busy <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_prs1_busy : io_core_dis_uops_0_bits_prs1_busy) : io_core_dis_uops_1_bits_prs1_busy) : io_core_dis_uops_2_bits_prs1_busy) : io_core_dis_uops_3_bits_prs1_busy);
    stq_31_bits_uop_prs2_busy <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_prs2_busy : io_core_dis_uops_0_bits_prs2_busy) : io_core_dis_uops_1_bits_prs2_busy) : io_core_dis_uops_2_bits_prs2_busy) : io_core_dis_uops_3_bits_prs2_busy);
    stq_31_bits_uop_prs3_busy <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_prs3_busy : io_core_dis_uops_0_bits_prs3_busy) : io_core_dis_uops_1_bits_prs3_busy) : io_core_dis_uops_2_bits_prs3_busy) : io_core_dis_uops_3_bits_prs3_busy);
    stq_31_bits_uop_ppred_busy <= ~_GEN_5750 & _GEN_2485 & _GEN_2165 & _GEN_2068 & _GEN_1684 & stq_31_bits_uop_ppred_busy;
    stq_31_bits_uop_exception <= ~_GEN_5750 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & (&mem_xcpt_uops_1_stq_idx) | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & (&mem_xcpt_uops_0_stq_idx) | (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_31_bits_uop_bypassable <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_bypassable : io_core_dis_uops_0_bits_bypassable) : io_core_dis_uops_1_bits_bypassable) : io_core_dis_uops_2_bits_bypassable) : io_core_dis_uops_3_bits_bypassable);
    stq_31_bits_uop_mem_signed <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_31_bits_uop_is_fence <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_31_bits_uop_is_fencei <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_fencei : io_core_dis_uops_0_bits_is_fencei) : io_core_dis_uops_1_bits_is_fencei) : io_core_dis_uops_2_bits_is_fencei) : io_core_dis_uops_3_bits_is_fencei);
    stq_31_bits_uop_is_amo <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_31_bits_uop_uses_ldq <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_31_bits_uop_uses_stq <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_31_bits_uop_is_sys_pc2epc <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_sys_pc2epc : io_core_dis_uops_0_bits_is_sys_pc2epc) : io_core_dis_uops_1_bits_is_sys_pc2epc) : io_core_dis_uops_2_bits_is_sys_pc2epc) : io_core_dis_uops_3_bits_is_sys_pc2epc);
    stq_31_bits_uop_is_unique <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_is_unique : io_core_dis_uops_0_bits_is_unique) : io_core_dis_uops_1_bits_is_unique) : io_core_dis_uops_2_bits_is_unique) : io_core_dis_uops_3_bits_is_unique);
    stq_31_bits_uop_flush_on_commit <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_flush_on_commit : io_core_dis_uops_0_bits_flush_on_commit) : io_core_dis_uops_1_bits_flush_on_commit) : io_core_dis_uops_2_bits_flush_on_commit) : io_core_dis_uops_3_bits_flush_on_commit);
    stq_31_bits_uop_ldst_is_rs1 <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_ldst_is_rs1 : io_core_dis_uops_0_bits_ldst_is_rs1) : io_core_dis_uops_1_bits_ldst_is_rs1) : io_core_dis_uops_2_bits_ldst_is_rs1) : io_core_dis_uops_3_bits_ldst_is_rs1);
    stq_31_bits_uop_ldst_val <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_ldst_val : io_core_dis_uops_0_bits_ldst_val) : io_core_dis_uops_1_bits_ldst_val) : io_core_dis_uops_2_bits_ldst_val) : io_core_dis_uops_3_bits_ldst_val);
    stq_31_bits_uop_frs3_en <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_frs3_en : io_core_dis_uops_0_bits_frs3_en) : io_core_dis_uops_1_bits_frs3_en) : io_core_dis_uops_2_bits_frs3_en) : io_core_dis_uops_3_bits_frs3_en);
    stq_31_bits_uop_fp_val <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_fp_val : io_core_dis_uops_0_bits_fp_val) : io_core_dis_uops_1_bits_fp_val) : io_core_dis_uops_2_bits_fp_val) : io_core_dis_uops_3_bits_fp_val);
    stq_31_bits_uop_fp_single <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_fp_single : io_core_dis_uops_0_bits_fp_single) : io_core_dis_uops_1_bits_fp_single) : io_core_dis_uops_2_bits_fp_single) : io_core_dis_uops_3_bits_fp_single);
    stq_31_bits_uop_xcpt_pf_if <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_xcpt_pf_if : io_core_dis_uops_0_bits_xcpt_pf_if) : io_core_dis_uops_1_bits_xcpt_pf_if) : io_core_dis_uops_2_bits_xcpt_pf_if) : io_core_dis_uops_3_bits_xcpt_pf_if);
    stq_31_bits_uop_xcpt_ae_if <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_xcpt_ae_if : io_core_dis_uops_0_bits_xcpt_ae_if) : io_core_dis_uops_1_bits_xcpt_ae_if) : io_core_dis_uops_2_bits_xcpt_ae_if) : io_core_dis_uops_3_bits_xcpt_ae_if);
    stq_31_bits_uop_xcpt_ma_if <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_xcpt_ma_if : io_core_dis_uops_0_bits_xcpt_ma_if) : io_core_dis_uops_1_bits_xcpt_ma_if) : io_core_dis_uops_2_bits_xcpt_ma_if) : io_core_dis_uops_3_bits_xcpt_ma_if);
    stq_31_bits_uop_bp_debug_if <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_bp_debug_if : io_core_dis_uops_0_bits_bp_debug_if) : io_core_dis_uops_1_bits_bp_debug_if) : io_core_dis_uops_2_bits_bp_debug_if) : io_core_dis_uops_3_bits_bp_debug_if);
    stq_31_bits_uop_bp_xcpt_if <= ~_GEN_5750 & (_GEN_2485 ? (_GEN_2165 ? (_GEN_2068 ? (_GEN_1684 ? stq_31_bits_uop_bp_xcpt_if : io_core_dis_uops_0_bits_bp_xcpt_if) : io_core_dis_uops_1_bits_bp_xcpt_if) : io_core_dis_uops_2_bits_bp_xcpt_if) : io_core_dis_uops_3_bits_bp_xcpt_if);
    stq_31_bits_addr_valid <= ~_GEN_5814 & (clear_store ? ~_GEN_5715 & _GEN_2868 : ~_GEN_5239 & _GEN_2868);
    if (_GEN_2867) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8)
          stq_31_bits_addr_bits <= exe_req_1_bits_addr;
        else if (will_fire_sfence_1_will_fire)
          stq_31_bits_addr_bits <= _GEN_273;
        else if (will_fire_load_retry_1_will_fire)
          stq_31_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_1_will_fire)
          stq_31_bits_addr_bits <= casez_tmp_290;
        else
          stq_31_bits_addr_bits <= _exe_tlb_vaddr_T_9;
      end
      else
        stq_31_bits_addr_bits <= _GEN_280;
      stq_31_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_2709) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1)
          stq_31_bits_addr_bits <= exe_req_0_bits_addr;
        else if (will_fire_sfence_0_will_fire)
          stq_31_bits_addr_bits <= _GEN_272;
        else if (will_fire_load_retry_0_will_fire)
          stq_31_bits_addr_bits <= casez_tmp_202;
        else if (will_fire_sta_retry_0_will_fire)
          stq_31_bits_addr_bits <= casez_tmp_290;
        else
          stq_31_bits_addr_bits <= _exe_tlb_vaddr_T_2;
      end
      else
        stq_31_bits_addr_bits <= _GEN_274;
      stq_31_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_31_bits_data_valid <= ~_GEN_5814 & (clear_store ? ~_GEN_5715 & _GEN_2931 : ~_GEN_5239 & _GEN_2931);
    if (_stq_bits_data_bits_T_2 & (&sidx_1))
      stq_31_bits_data_bits <= _stq_bits_data_bits_T_3;
    else if (_GEN_2741)
      stq_31_bits_data_bits <= _stq_bits_data_bits_T_1;
    stq_31_bits_committed <= ~_GEN_5747 & (commit_store_3 ? (&idx_3) | _GEN_5557 | _GEN_5462 : _GEN_5557 | _GEN_5462);
    stq_31_bits_succeeded <= ~_GEN_5747 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & (&io_dmem_resp_1_bits_uop_stq_idx) | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & (&io_dmem_resp_0_bits_uop_stq_idx) | (_GEN_281 | ~(will_fire_store_commit_1_will_fire & (&stq_execute_head))) & (_GEN_275 | ~(will_fire_store_commit_0_will_fire & (&stq_execute_head))) & _GEN_2485 & _GEN_2165 & _GEN_2068 & _GEN_1684 & stq_31_bits_succeeded);
    if (_GEN_5749) begin
      ldq_head <= 5'h0;
      ldq_tail <= 5'h0;
      stq_tail <= reset ? 5'h0 : stq_commit_head;
    end
    else begin
      if (commit_load_3)
        ldq_head <= _GEN_1557 + 5'h1;
      else if (commit_load_2)
        ldq_head <= _GEN_1556;
      else if (commit_load_1)
        ldq_head <= _GEN_1551;
      else if (commit_load)
        ldq_head <= _GEN_1546;
      if (io_core_brupdate_b2_mispredict & ~io_core_exception) begin
        ldq_tail <= io_core_brupdate_b2_uop_ldq_idx;
        stq_tail <= io_core_brupdate_b2_uop_stq_idx;
      end
      else begin
        if (dis_ld_val_3)
          ldq_tail <= _GEN_15;
        else if (dis_ld_val_2)
          ldq_tail <= _GEN_11;
        else if (dis_ld_val_1)
          ldq_tail <= _GEN_7;
        else if (dis_ld_val)
          ldq_tail <= _GEN_3;
        if (dis_st_val_3)
          stq_tail <= _GEN_16;
        else if (dis_st_val_2)
          stq_tail <= _GEN_12;
        else if (dis_st_val_1)
          stq_tail <= _GEN_8;
        else if (dis_st_val)
          stq_tail <= _GEN_4;
      end
    end
    if (_io_hellacache_req_ready_output & _GEN_1579)
      hella_req_addr <= io_hellacache_req_bits_addr;
    if (_GEN_5748) begin
    end
    else
      hella_data_data <= 64'h0;
    if (will_fire_load_incoming_1_will_fire | will_fire_load_retry_1_will_fire | _GEN_282 | ~will_fire_hella_incoming_1_will_fire) begin
      if (will_fire_load_incoming_0_will_fire | will_fire_load_retry_0_will_fire | _GEN_276 | ~will_fire_hella_incoming_0_will_fire) begin
      end
      else
        hella_paddr <= exe_tlb_paddr_0;
    end
    else
      hella_paddr <= exe_tlb_paddr_1;
    if (_GEN_5748) begin
    end
    else begin
      hella_xcpt_ma_ld <= _dtlb_io_resp_1_ma_ld;
      hella_xcpt_ma_st <= _dtlb_io_resp_1_ma_st;
      hella_xcpt_pf_ld <= _dtlb_io_resp_1_pf_ld;
      hella_xcpt_pf_st <= _dtlb_io_resp_1_pf_st;
    end
    hella_xcpt_gf_ld <= _GEN_5748 & hella_xcpt_gf_ld;
    hella_xcpt_gf_st <= _GEN_5748 & hella_xcpt_gf_st;
    if (_GEN_5748) begin
    end
    else begin
      hella_xcpt_ae_ld <= _dtlb_io_resp_1_ae_ld;
      hella_xcpt_ae_st <= _dtlb_io_resp_1_ae_st;
    end
    if (will_fire_load_wakeup_1_will_fire) begin
      p1_block_load_mask_0 <= _GEN_145;
      p1_block_load_mask_1 <= _GEN_146;
      p1_block_load_mask_2 <= _GEN_147;
      p1_block_load_mask_3 <= _GEN_148;
      p1_block_load_mask_4 <= _GEN_149;
      p1_block_load_mask_5 <= _GEN_150;
      p1_block_load_mask_6 <= _GEN_151;
      p1_block_load_mask_7 <= _GEN_152;
      p1_block_load_mask_8 <= _GEN_153;
      p1_block_load_mask_9 <= _GEN_154;
      p1_block_load_mask_10 <= _GEN_155;
      p1_block_load_mask_11 <= _GEN_156;
      p1_block_load_mask_12 <= _GEN_157;
      p1_block_load_mask_13 <= _GEN_158;
      p1_block_load_mask_14 <= _GEN_159;
      p1_block_load_mask_15 <= _GEN_160;
      p1_block_load_mask_16 <= _GEN_161;
      p1_block_load_mask_17 <= _GEN_162;
      p1_block_load_mask_18 <= _GEN_163;
      p1_block_load_mask_19 <= _GEN_164;
      p1_block_load_mask_20 <= _GEN_165;
      p1_block_load_mask_21 <= _GEN_166;
      p1_block_load_mask_22 <= _GEN_167;
      p1_block_load_mask_23 <= _GEN_168;
      p1_block_load_mask_24 <= _GEN_169;
      p1_block_load_mask_25 <= _GEN_170;
      p1_block_load_mask_26 <= _GEN_171;
      p1_block_load_mask_27 <= _GEN_172;
      p1_block_load_mask_28 <= _GEN_173;
      p1_block_load_mask_29 <= _GEN_174;
      p1_block_load_mask_30 <= _GEN_175;
      p1_block_load_mask_31 <= _GEN_176;
    end
    else if (will_fire_load_incoming_1_will_fire) begin
      p1_block_load_mask_0 <= _GEN_178;
      p1_block_load_mask_1 <= _GEN_180;
      p1_block_load_mask_2 <= _GEN_182;
      p1_block_load_mask_3 <= _GEN_184;
      p1_block_load_mask_4 <= _GEN_186;
      p1_block_load_mask_5 <= _GEN_188;
      p1_block_load_mask_6 <= _GEN_190;
      p1_block_load_mask_7 <= _GEN_192;
      p1_block_load_mask_8 <= _GEN_194;
      p1_block_load_mask_9 <= _GEN_196;
      p1_block_load_mask_10 <= _GEN_198;
      p1_block_load_mask_11 <= _GEN_200;
      p1_block_load_mask_12 <= _GEN_202;
      p1_block_load_mask_13 <= _GEN_204;
      p1_block_load_mask_14 <= _GEN_206;
      p1_block_load_mask_15 <= _GEN_208;
      p1_block_load_mask_16 <= _GEN_210;
      p1_block_load_mask_17 <= _GEN_212;
      p1_block_load_mask_18 <= _GEN_214;
      p1_block_load_mask_19 <= _GEN_216;
      p1_block_load_mask_20 <= _GEN_218;
      p1_block_load_mask_21 <= _GEN_220;
      p1_block_load_mask_22 <= _GEN_222;
      p1_block_load_mask_23 <= _GEN_224;
      p1_block_load_mask_24 <= _GEN_226;
      p1_block_load_mask_25 <= _GEN_228;
      p1_block_load_mask_26 <= _GEN_230;
      p1_block_load_mask_27 <= _GEN_232;
      p1_block_load_mask_28 <= _GEN_234;
      p1_block_load_mask_29 <= _GEN_236;
      p1_block_load_mask_30 <= _GEN_238;
      p1_block_load_mask_31 <= _GEN_239;
    end
    else begin
      p1_block_load_mask_0 <= _GEN_240;
      p1_block_load_mask_1 <= _GEN_241;
      p1_block_load_mask_2 <= _GEN_242;
      p1_block_load_mask_3 <= _GEN_243;
      p1_block_load_mask_4 <= _GEN_244;
      p1_block_load_mask_5 <= _GEN_245;
      p1_block_load_mask_6 <= _GEN_246;
      p1_block_load_mask_7 <= _GEN_247;
      p1_block_load_mask_8 <= _GEN_248;
      p1_block_load_mask_9 <= _GEN_249;
      p1_block_load_mask_10 <= _GEN_250;
      p1_block_load_mask_11 <= _GEN_251;
      p1_block_load_mask_12 <= _GEN_252;
      p1_block_load_mask_13 <= _GEN_253;
      p1_block_load_mask_14 <= _GEN_254;
      p1_block_load_mask_15 <= _GEN_255;
      p1_block_load_mask_16 <= _GEN_256;
      p1_block_load_mask_17 <= _GEN_257;
      p1_block_load_mask_18 <= _GEN_258;
      p1_block_load_mask_19 <= _GEN_259;
      p1_block_load_mask_20 <= _GEN_260;
      p1_block_load_mask_21 <= _GEN_261;
      p1_block_load_mask_22 <= _GEN_262;
      p1_block_load_mask_23 <= _GEN_263;
      p1_block_load_mask_24 <= _GEN_264;
      p1_block_load_mask_25 <= _GEN_265;
      p1_block_load_mask_26 <= _GEN_266;
      p1_block_load_mask_27 <= _GEN_267;
      p1_block_load_mask_28 <= _GEN_268;
      p1_block_load_mask_29 <= _GEN_269;
      p1_block_load_mask_30 <= _GEN_270;
      p1_block_load_mask_31 <= _GEN_271;
    end
    p2_block_load_mask_0 <= p1_block_load_mask_0;
    p2_block_load_mask_1 <= p1_block_load_mask_1;
    p2_block_load_mask_2 <= p1_block_load_mask_2;
    p2_block_load_mask_3 <= p1_block_load_mask_3;
    p2_block_load_mask_4 <= p1_block_load_mask_4;
    p2_block_load_mask_5 <= p1_block_load_mask_5;
    p2_block_load_mask_6 <= p1_block_load_mask_6;
    p2_block_load_mask_7 <= p1_block_load_mask_7;
    p2_block_load_mask_8 <= p1_block_load_mask_8;
    p2_block_load_mask_9 <= p1_block_load_mask_9;
    p2_block_load_mask_10 <= p1_block_load_mask_10;
    p2_block_load_mask_11 <= p1_block_load_mask_11;
    p2_block_load_mask_12 <= p1_block_load_mask_12;
    p2_block_load_mask_13 <= p1_block_load_mask_13;
    p2_block_load_mask_14 <= p1_block_load_mask_14;
    p2_block_load_mask_15 <= p1_block_load_mask_15;
    p2_block_load_mask_16 <= p1_block_load_mask_16;
    p2_block_load_mask_17 <= p1_block_load_mask_17;
    p2_block_load_mask_18 <= p1_block_load_mask_18;
    p2_block_load_mask_19 <= p1_block_load_mask_19;
    p2_block_load_mask_20 <= p1_block_load_mask_20;
    p2_block_load_mask_21 <= p1_block_load_mask_21;
    p2_block_load_mask_22 <= p1_block_load_mask_22;
    p2_block_load_mask_23 <= p1_block_load_mask_23;
    p2_block_load_mask_24 <= p1_block_load_mask_24;
    p2_block_load_mask_25 <= p1_block_load_mask_25;
    p2_block_load_mask_26 <= p1_block_load_mask_26;
    p2_block_load_mask_27 <= p1_block_load_mask_27;
    p2_block_load_mask_28 <= p1_block_load_mask_28;
    p2_block_load_mask_29 <= p1_block_load_mask_29;
    p2_block_load_mask_30 <= p1_block_load_mask_30;
    p2_block_load_mask_31 <= p1_block_load_mask_31;
    ldq_retry_idx <= _ldq_retry_idx_T_2 & _temp_bits_T ? 5'h0 : _ldq_retry_idx_T_5 & _temp_bits_T_2 ? 5'h1 : _ldq_retry_idx_T_8 & _temp_bits_T_4 ? 5'h2 : _ldq_retry_idx_T_11 & _temp_bits_T_6 ? 5'h3 : _ldq_retry_idx_T_14 & _temp_bits_T_8 ? 5'h4 : _ldq_retry_idx_T_17 & _temp_bits_T_10 ? 5'h5 : _ldq_retry_idx_T_20 & _temp_bits_T_12 ? 5'h6 : _ldq_retry_idx_T_23 & _temp_bits_T_14 ? 5'h7 : _ldq_retry_idx_T_26 & _temp_bits_T_16 ? 5'h8 : _ldq_retry_idx_T_29 & _temp_bits_T_18 ? 5'h9 : _ldq_retry_idx_T_32 & _temp_bits_T_20 ? 5'hA : _ldq_retry_idx_T_35 & _temp_bits_T_22 ? 5'hB : _ldq_retry_idx_T_38 & _temp_bits_T_24 ? 5'hC : _ldq_retry_idx_T_41 & _temp_bits_T_26 ? 5'hD : _ldq_retry_idx_T_44 & _temp_bits_T_28 ? 5'hE : _ldq_retry_idx_T_47 & ~(ldq_head[4]) ? 5'hF : _ldq_retry_idx_T_50 & _temp_bits_T_32 ? 5'h10 : _ldq_retry_idx_T_53 & _temp_bits_T_34 ? 5'h11 : _ldq_retry_idx_T_56 & _temp_bits_T_36 ? 5'h12 : _ldq_retry_idx_T_59 & _temp_bits_T_38 ? 5'h13 : _ldq_retry_idx_idx_T_42[4:0];
    stq_retry_idx <= _stq_retry_idx_T & stq_commit_head == 5'h0 ? 5'h0 : _stq_retry_idx_T_1 & stq_commit_head < 5'h2 ? 5'h1 : _stq_retry_idx_T_2 & stq_commit_head < 5'h3 ? 5'h2 : _stq_retry_idx_T_3 & stq_commit_head < 5'h4 ? 5'h3 : _stq_retry_idx_T_4 & stq_commit_head < 5'h5 ? 5'h4 : _stq_retry_idx_T_5 & stq_commit_head < 5'h6 ? 5'h5 : _stq_retry_idx_T_6 & stq_commit_head < 5'h7 ? 5'h6 : _stq_retry_idx_T_7 & stq_commit_head < 5'h8 ? 5'h7 : _stq_retry_idx_T_8 & stq_commit_head < 5'h9 ? 5'h8 : _stq_retry_idx_T_9 & stq_commit_head < 5'hA ? 5'h9 : _stq_retry_idx_T_10 & stq_commit_head < 5'hB ? 5'hA : _stq_retry_idx_T_11 & stq_commit_head < 5'hC ? 5'hB : _stq_retry_idx_T_12 & stq_commit_head < 5'hD ? 5'hC : _stq_retry_idx_T_13 & stq_commit_head < 5'hE ? 5'hD : _stq_retry_idx_T_14 & stq_commit_head < 5'hF ? 5'hE : _stq_retry_idx_T_15 & ~(stq_commit_head[4]) ? 5'hF : _stq_retry_idx_T_16 & stq_commit_head < 5'h11 ? 5'h10 : _stq_retry_idx_T_17 & stq_commit_head < 5'h12 ? 5'h11 : _stq_retry_idx_T_18 & stq_commit_head < 5'h13 ? 5'h12 : _stq_retry_idx_T_19 & stq_commit_head < 5'h14 ? 5'h13 : _stq_retry_idx_idx_T_42[4:0];
    ldq_wakeup_idx <= _ldq_wakeup_idx_T_7 & _temp_bits_T ? 5'h0 : _ldq_wakeup_idx_T_15 & _temp_bits_T_2 ? 5'h1 : _ldq_wakeup_idx_T_23 & _temp_bits_T_4 ? 5'h2 : _ldq_wakeup_idx_T_31 & _temp_bits_T_6 ? 5'h3 : _ldq_wakeup_idx_T_39 & _temp_bits_T_8 ? 5'h4 : _ldq_wakeup_idx_T_47 & _temp_bits_T_10 ? 5'h5 : _ldq_wakeup_idx_T_55 & _temp_bits_T_12 ? 5'h6 : _ldq_wakeup_idx_T_63 & _temp_bits_T_14 ? 5'h7 : _ldq_wakeup_idx_T_71 & _temp_bits_T_16 ? 5'h8 : _ldq_wakeup_idx_T_79 & _temp_bits_T_18 ? 5'h9 : _ldq_wakeup_idx_T_87 & _temp_bits_T_20 ? 5'hA : _ldq_wakeup_idx_T_95 & _temp_bits_T_22 ? 5'hB : _ldq_wakeup_idx_T_103 & _temp_bits_T_24 ? 5'hC : _ldq_wakeup_idx_T_111 & _temp_bits_T_26 ? 5'hD : _ldq_wakeup_idx_T_119 & _temp_bits_T_28 ? 5'hE : _ldq_wakeup_idx_T_127 & ~(ldq_head[4]) ? 5'hF : _ldq_wakeup_idx_T_135 & _temp_bits_T_32 ? 5'h10 : _ldq_wakeup_idx_T_143 & _temp_bits_T_34 ? 5'h11 : _ldq_wakeup_idx_T_151 & _temp_bits_T_36 ? 5'h12 : _ldq_wakeup_idx_T_159 & _temp_bits_T_38 ? 5'h13 : _ldq_wakeup_idx_idx_T_42[4:0];
    can_fire_load_retry_REG_1 <= _dtlb_io_miss_rdy;
    can_fire_sta_retry_REG_1 <= _dtlb_io_miss_rdy;
    mem_xcpt_valids_0 <= (pf_ld_0 | pf_st_0 | ae_ld_0 | ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_ae_st & _mem_xcpt_uops_WIRE_0_uses_stq | ma_ld_0 | ma_st_0) & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & exe_tlb_uop_0_br_mask) == 20'h0;
    mem_xcpt_valids_1 <= (pf_ld_1 | pf_st_1 | ae_ld_1 | ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_ae_st & _mem_xcpt_uops_WIRE_1_uses_stq | ma_ld_1 | ma_st_1) & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & exe_tlb_uop_1_br_mask) == 20'h0;
    mem_xcpt_uops_0_br_mask <= exe_tlb_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask;
    mem_xcpt_uops_0_rob_idx <= _mem_xcpt_uops_WIRE_0_rob_idx;
    mem_xcpt_uops_0_ldq_idx <= _mem_xcpt_uops_WIRE_0_ldq_idx;
    mem_xcpt_uops_0_stq_idx <= _mem_xcpt_uops_WIRE_0_stq_idx;
    mem_xcpt_uops_0_uses_ldq <= _mem_xcpt_uops_WIRE_0_uses_ldq;
    mem_xcpt_uops_0_uses_stq <= _mem_xcpt_uops_WIRE_0_uses_stq;
    mem_xcpt_uops_1_br_mask <= exe_tlb_uop_1_br_mask & ~io_core_brupdate_b1_resolve_mask;
    mem_xcpt_uops_1_rob_idx <= _mem_xcpt_uops_WIRE_1_rob_idx;
    mem_xcpt_uops_1_ldq_idx <= _mem_xcpt_uops_WIRE_1_ldq_idx;
    mem_xcpt_uops_1_stq_idx <= _mem_xcpt_uops_WIRE_1_stq_idx;
    mem_xcpt_uops_1_uses_ldq <= _mem_xcpt_uops_WIRE_1_uses_ldq;
    mem_xcpt_uops_1_uses_stq <= _mem_xcpt_uops_WIRE_1_uses_stq;
    mem_xcpt_causes_0 <= ma_ld_0 ? 4'h4 : ma_st_0 ? 4'h6 : pf_ld_0 ? 4'hD : pf_st_0 ? 4'hF : {2'h1, ~ae_ld_0, 1'h1};
    mem_xcpt_causes_1 <= ma_ld_1 ? 4'h4 : ma_st_1 ? 4'h6 : pf_ld_1 ? 4'hD : pf_st_1 ? 4'hF : {2'h1, ~ae_ld_1, 1'h1};
    mem_xcpt_vaddrs_0 <= exe_tlb_vaddr_0;
    mem_xcpt_vaddrs_1 <= exe_tlb_vaddr_1;
    REG <= _GEN_18 | will_fire_load_retry_0_will_fire | will_fire_sta_retry_0_will_fire;
    REG_1 <= _GEN_144 | will_fire_load_retry_1_will_fire | will_fire_sta_retry_1_will_fire;
    fired_load_incoming_REG <= will_fire_load_incoming_0_will_fire & _fired_std_incoming_T;
    fired_load_incoming_REG_1 <= will_fire_load_incoming_1_will_fire & _fired_std_incoming_T_2;
    fired_stad_incoming_REG <= will_fire_stad_incoming_0_will_fire & _fired_std_incoming_T;
    fired_stad_incoming_REG_1 <= will_fire_stad_incoming_1_will_fire & _fired_std_incoming_T_2;
    fired_sta_incoming_REG <= will_fire_sta_incoming_0_will_fire & _fired_std_incoming_T;
    fired_sta_incoming_REG_1 <= will_fire_sta_incoming_1_will_fire & _fired_std_incoming_T_2;
    fired_std_incoming_REG <= will_fire_std_incoming_0_will_fire & _fired_std_incoming_T;
    fired_std_incoming_REG_1 <= will_fire_std_incoming_1_will_fire & _fired_std_incoming_T_2;
    fired_stdf_incoming <= fp_stdata_fire & (io_core_brupdate_b1_mispredict_mask & io_core_fp_stdata_bits_uop_br_mask) == 20'h0;
    fired_sfence_0 <= will_fire_sfence_0_will_fire;
    fired_sfence_1 <= will_fire_sfence_1_will_fire;
    fired_release_0 <= will_fire_release_0_will_fire;
    fired_release_1 <= will_fire_release_1_will_fire;
    fired_load_retry_REG <= will_fire_load_retry_0_will_fire & _mem_ldq_retry_e_out_valid_T == 20'h0;
    fired_load_retry_REG_1 <= will_fire_load_retry_1_will_fire & _mem_ldq_retry_e_out_valid_T == 20'h0;
    fired_sta_retry_REG <= will_fire_sta_retry_0_will_fire & _mem_stq_retry_e_out_valid_T == 20'h0;
    fired_sta_retry_REG_1 <= will_fire_sta_retry_1_will_fire & _mem_stq_retry_e_out_valid_T == 20'h0;
    fired_load_wakeup_REG <= will_fire_load_wakeup_0_will_fire & _mem_ldq_wakeup_e_out_valid_T == 20'h0;
    fired_load_wakeup_REG_1 <= will_fire_load_wakeup_1_will_fire & _mem_ldq_wakeup_e_out_valid_T == 20'h0;
    mem_incoming_uop_0_br_mask <= exe_req_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    mem_incoming_uop_0_rob_idx <= _mem_incoming_uop_WIRE_0_rob_idx;
    mem_incoming_uop_0_ldq_idx <= _mem_incoming_uop_WIRE_0_ldq_idx;
    mem_incoming_uop_0_stq_idx <= _mem_incoming_uop_WIRE_0_stq_idx;
    mem_incoming_uop_0_pdst <= _mem_incoming_uop_WIRE_0_pdst;
    mem_incoming_uop_0_fp_val <= _mem_incoming_uop_WIRE_0_fp_val;
    mem_incoming_uop_1_br_mask <= exe_req_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    mem_incoming_uop_1_rob_idx <= _mem_incoming_uop_WIRE_1_rob_idx;
    mem_incoming_uop_1_ldq_idx <= _mem_incoming_uop_WIRE_1_ldq_idx;
    mem_incoming_uop_1_stq_idx <= _mem_incoming_uop_WIRE_1_stq_idx;
    mem_incoming_uop_1_pdst <= _mem_incoming_uop_WIRE_1_pdst;
    mem_incoming_uop_1_fp_val <= _mem_incoming_uop_WIRE_1_fp_val;
    mem_ldq_incoming_e_0_bits_uop_br_mask <= casez_tmp_93 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_incoming_e_0_bits_uop_stq_idx <= casez_tmp_94;
    mem_ldq_incoming_e_0_bits_uop_mem_size <= casez_tmp_95;
    mem_ldq_incoming_e_0_bits_st_dep_mask <= casez_tmp_98;
    mem_ldq_incoming_e_1_bits_uop_br_mask <= casez_tmp_99 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_incoming_e_1_bits_uop_stq_idx <= casez_tmp_100;
    mem_ldq_incoming_e_1_bits_uop_mem_size <= casez_tmp_101;
    mem_ldq_incoming_e_1_bits_st_dep_mask <= casez_tmp_104;
    mem_stq_incoming_e_0_valid <= casez_tmp_105 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_106) == 20'h0;
    mem_stq_incoming_e_0_bits_uop_br_mask <= casez_tmp_106 & ~io_core_brupdate_b1_resolve_mask;
    mem_stq_incoming_e_0_bits_uop_rob_idx <= casez_tmp_107;
    mem_stq_incoming_e_0_bits_uop_stq_idx <= casez_tmp_108;
    mem_stq_incoming_e_0_bits_uop_mem_size <= casez_tmp_109;
    mem_stq_incoming_e_0_bits_uop_is_amo <= casez_tmp_110;
    mem_stq_incoming_e_0_bits_addr_valid <= casez_tmp_111;
    mem_stq_incoming_e_0_bits_addr_is_virtual <= casez_tmp_112;
    mem_stq_incoming_e_0_bits_data_valid <= casez_tmp_113;
    mem_stq_incoming_e_1_valid <= casez_tmp_114 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_115) == 20'h0;
    mem_stq_incoming_e_1_bits_uop_br_mask <= casez_tmp_115 & ~io_core_brupdate_b1_resolve_mask;
    mem_stq_incoming_e_1_bits_uop_rob_idx <= casez_tmp_116;
    mem_stq_incoming_e_1_bits_uop_stq_idx <= casez_tmp_117;
    mem_stq_incoming_e_1_bits_uop_mem_size <= casez_tmp_118;
    mem_stq_incoming_e_1_bits_uop_is_amo <= casez_tmp_119;
    mem_stq_incoming_e_1_bits_addr_valid <= casez_tmp_120;
    mem_stq_incoming_e_1_bits_addr_is_virtual <= casez_tmp_121;
    mem_stq_incoming_e_1_bits_data_valid <= casez_tmp_122;
    mem_ldq_wakeup_e_bits_uop_br_mask <= casez_tmp_318 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_wakeup_e_bits_uop_stq_idx <= casez_tmp_328;
    mem_ldq_wakeup_e_bits_uop_mem_size <= casez_tmp_342;
    mem_ldq_wakeup_e_bits_st_dep_mask <= casez_tmp_378;
    mem_ldq_retry_e_bits_uop_br_mask <= casez_tmp_148 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_retry_e_bits_uop_stq_idx <= casez_tmp_158;
    mem_ldq_retry_e_bits_uop_mem_size <= casez_tmp_172;
    mem_ldq_retry_e_bits_st_dep_mask <= casez_tmp_206;
    mem_stq_retry_e_valid <= casez_tmp_209 & _mem_stq_retry_e_out_valid_T == 20'h0;
    mem_stq_retry_e_bits_uop_br_mask <= casez_tmp_234 & ~io_core_brupdate_b1_resolve_mask;
    mem_stq_retry_e_bits_uop_rob_idx <= casez_tmp_242;
    mem_stq_retry_e_bits_uop_stq_idx <= casez_tmp_244;
    mem_stq_retry_e_bits_uop_mem_size <= casez_tmp_260;
    mem_stq_retry_e_bits_uop_is_amo <= casez_tmp_264;
    mem_stq_retry_e_bits_data_valid <= casez_tmp_292;
    mem_stdf_uop_br_mask <= io_core_fp_stdata_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    mem_stdf_uop_rob_idx <= io_core_fp_stdata_bits_uop_rob_idx;
    mem_stdf_uop_stq_idx <= io_core_fp_stdata_bits_uop_stq_idx;
    mem_tlb_miss_0 <= exe_tlb_miss_0;
    mem_tlb_miss_1 <= exe_tlb_miss_1;
    mem_tlb_uncacheable_0 <= ~_dtlb_io_resp_0_cacheable;
    mem_tlb_uncacheable_1 <= ~_dtlb_io_resp_1_cacheable;
    mem_paddr_0 <= _mem_paddr_WIRE_0;
    mem_paddr_1 <= _mem_paddr_WIRE_1;
    clr_bsy_rob_idx_0 <= fired_stad_incoming_REG | fired_sta_incoming_REG | fired_std_incoming_REG ? mem_stq_incoming_e_0_bits_uop_rob_idx : fired_sfence_0 ? mem_incoming_uop_0_rob_idx : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_rob_idx : 7'h0;
    clr_bsy_rob_idx_1 <= fired_stad_incoming_REG_1 | fired_sta_incoming_REG_1 | fired_std_incoming_REG_1 ? mem_stq_incoming_e_1_bits_uop_rob_idx : fired_sfence_1 ? mem_incoming_uop_1_rob_idx : fired_sta_retry_REG_1 ? mem_stq_retry_e_bits_uop_rob_idx : 7'h0;
    clr_bsy_brmask_0 <= fired_stad_incoming_REG ? mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_sta_incoming_REG ? mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_std_incoming_REG ? mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_sfence_0 ? mem_incoming_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : 20'h0;
    clr_bsy_brmask_1 <= fired_stad_incoming_REG_1 ? mem_stq_incoming_e_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_sta_incoming_REG_1 ? mem_stq_incoming_e_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_std_incoming_REG_1 ? mem_stq_incoming_e_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_sfence_1 ? mem_incoming_uop_1_br_mask & ~io_core_brupdate_b1_resolve_mask : fired_sta_retry_REG_1 ? mem_stq_retry_e_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : 20'h0;
    io_core_clr_bsy_0_valid_REG <= io_core_exception;
    io_core_clr_bsy_0_valid_REG_1 <= io_core_exception;
    io_core_clr_bsy_0_valid_REG_2 <= io_core_clr_bsy_0_valid_REG_1;
    io_core_clr_bsy_1_valid_REG <= io_core_exception;
    io_core_clr_bsy_1_valid_REG_1 <= io_core_exception;
    io_core_clr_bsy_1_valid_REG_2 <= io_core_clr_bsy_1_valid_REG_1;
    stdf_clr_bsy_rob_idx <= fired_stdf_incoming ? mem_stdf_uop_rob_idx : 7'h0;
    stdf_clr_bsy_brmask <= fired_stdf_incoming ? mem_stdf_uop_br_mask & ~io_core_brupdate_b1_resolve_mask : 20'h0;
    io_core_clr_bsy_2_valid_REG <= io_core_exception;
    io_core_clr_bsy_2_valid_REG_1 <= io_core_exception;
    io_core_clr_bsy_2_valid_REG_2 <= io_core_clr_bsy_2_valid_REG_1;
    lcam_addr_REG <= exe_tlb_paddr_0;
    lcam_addr_REG_1 <= io_dmem_release_bits_address;
    lcam_addr_REG_2 <= exe_tlb_paddr_1;
    lcam_addr_REG_3 <= io_dmem_release_bits_address;
    lcam_ldq_idx_REG <= ldq_wakeup_idx;
    lcam_ldq_idx_REG_1 <= ldq_retry_idx;
    lcam_ldq_idx_REG_2 <= ldq_wakeup_idx;
    lcam_ldq_idx_REG_3 <= ldq_retry_idx;
    lcam_stq_idx_REG <= stq_retry_idx;
    lcam_stq_idx_REG_1 <= stq_retry_idx;
    s1_executing_loads_0 <= will_fire_load_incoming_1_will_fire ? (_GEN_177 ? dmem_req_fire_1 : _GEN_2614) : will_fire_load_retry_1_will_fire ? (_GEN_81 ? dmem_req_fire_1 : _GEN_2614) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_19) ? _GEN_2614 : dmem_req_fire_1;
    s1_executing_loads_1 <= will_fire_load_incoming_1_will_fire ? (_GEN_179 ? dmem_req_fire_1 : _GEN_2615) : will_fire_load_retry_1_will_fire ? (_GEN_83 ? dmem_req_fire_1 : _GEN_2615) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_20) ? _GEN_2615 : dmem_req_fire_1;
    s1_executing_loads_2 <= will_fire_load_incoming_1_will_fire ? (_GEN_181 ? dmem_req_fire_1 : _GEN_2616) : will_fire_load_retry_1_will_fire ? (_GEN_85 ? dmem_req_fire_1 : _GEN_2616) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_21) ? _GEN_2616 : dmem_req_fire_1;
    s1_executing_loads_3 <= will_fire_load_incoming_1_will_fire ? (_GEN_183 ? dmem_req_fire_1 : _GEN_2617) : will_fire_load_retry_1_will_fire ? (_GEN_87 ? dmem_req_fire_1 : _GEN_2617) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_22) ? _GEN_2617 : dmem_req_fire_1;
    s1_executing_loads_4 <= will_fire_load_incoming_1_will_fire ? (_GEN_185 ? dmem_req_fire_1 : _GEN_2618) : will_fire_load_retry_1_will_fire ? (_GEN_89 ? dmem_req_fire_1 : _GEN_2618) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_23) ? _GEN_2618 : dmem_req_fire_1;
    s1_executing_loads_5 <= will_fire_load_incoming_1_will_fire ? (_GEN_187 ? dmem_req_fire_1 : _GEN_2619) : will_fire_load_retry_1_will_fire ? (_GEN_91 ? dmem_req_fire_1 : _GEN_2619) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_24) ? _GEN_2619 : dmem_req_fire_1;
    s1_executing_loads_6 <= will_fire_load_incoming_1_will_fire ? (_GEN_189 ? dmem_req_fire_1 : _GEN_2620) : will_fire_load_retry_1_will_fire ? (_GEN_93 ? dmem_req_fire_1 : _GEN_2620) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_25) ? _GEN_2620 : dmem_req_fire_1;
    s1_executing_loads_7 <= will_fire_load_incoming_1_will_fire ? (_GEN_191 ? dmem_req_fire_1 : _GEN_2621) : will_fire_load_retry_1_will_fire ? (_GEN_95 ? dmem_req_fire_1 : _GEN_2621) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_26) ? _GEN_2621 : dmem_req_fire_1;
    s1_executing_loads_8 <= will_fire_load_incoming_1_will_fire ? (_GEN_193 ? dmem_req_fire_1 : _GEN_2622) : will_fire_load_retry_1_will_fire ? (_GEN_97 ? dmem_req_fire_1 : _GEN_2622) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_27) ? _GEN_2622 : dmem_req_fire_1;
    s1_executing_loads_9 <= will_fire_load_incoming_1_will_fire ? (_GEN_195 ? dmem_req_fire_1 : _GEN_2623) : will_fire_load_retry_1_will_fire ? (_GEN_99 ? dmem_req_fire_1 : _GEN_2623) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_28) ? _GEN_2623 : dmem_req_fire_1;
    s1_executing_loads_10 <= will_fire_load_incoming_1_will_fire ? (_GEN_197 ? dmem_req_fire_1 : _GEN_2624) : will_fire_load_retry_1_will_fire ? (_GEN_101 ? dmem_req_fire_1 : _GEN_2624) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_29) ? _GEN_2624 : dmem_req_fire_1;
    s1_executing_loads_11 <= will_fire_load_incoming_1_will_fire ? (_GEN_199 ? dmem_req_fire_1 : _GEN_2625) : will_fire_load_retry_1_will_fire ? (_GEN_103 ? dmem_req_fire_1 : _GEN_2625) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_30) ? _GEN_2625 : dmem_req_fire_1;
    s1_executing_loads_12 <= will_fire_load_incoming_1_will_fire ? (_GEN_201 ? dmem_req_fire_1 : _GEN_2626) : will_fire_load_retry_1_will_fire ? (_GEN_105 ? dmem_req_fire_1 : _GEN_2626) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_31) ? _GEN_2626 : dmem_req_fire_1;
    s1_executing_loads_13 <= will_fire_load_incoming_1_will_fire ? (_GEN_203 ? dmem_req_fire_1 : _GEN_2627) : will_fire_load_retry_1_will_fire ? (_GEN_107 ? dmem_req_fire_1 : _GEN_2627) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_32) ? _GEN_2627 : dmem_req_fire_1;
    s1_executing_loads_14 <= will_fire_load_incoming_1_will_fire ? (_GEN_205 ? dmem_req_fire_1 : _GEN_2628) : will_fire_load_retry_1_will_fire ? (_GEN_109 ? dmem_req_fire_1 : _GEN_2628) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_33) ? _GEN_2628 : dmem_req_fire_1;
    s1_executing_loads_15 <= will_fire_load_incoming_1_will_fire ? (_GEN_207 ? dmem_req_fire_1 : _GEN_2629) : will_fire_load_retry_1_will_fire ? (_GEN_111 ? dmem_req_fire_1 : _GEN_2629) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_34) ? _GEN_2629 : dmem_req_fire_1;
    s1_executing_loads_16 <= will_fire_load_incoming_1_will_fire ? (_GEN_209 ? dmem_req_fire_1 : _GEN_2630) : will_fire_load_retry_1_will_fire ? (_GEN_113 ? dmem_req_fire_1 : _GEN_2630) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_35) ? _GEN_2630 : dmem_req_fire_1;
    s1_executing_loads_17 <= will_fire_load_incoming_1_will_fire ? (_GEN_211 ? dmem_req_fire_1 : _GEN_2631) : will_fire_load_retry_1_will_fire ? (_GEN_115 ? dmem_req_fire_1 : _GEN_2631) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_36) ? _GEN_2631 : dmem_req_fire_1;
    s1_executing_loads_18 <= will_fire_load_incoming_1_will_fire ? (_GEN_213 ? dmem_req_fire_1 : _GEN_2632) : will_fire_load_retry_1_will_fire ? (_GEN_117 ? dmem_req_fire_1 : _GEN_2632) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_37) ? _GEN_2632 : dmem_req_fire_1;
    s1_executing_loads_19 <= will_fire_load_incoming_1_will_fire ? (_GEN_215 ? dmem_req_fire_1 : _GEN_2633) : will_fire_load_retry_1_will_fire ? (_GEN_119 ? dmem_req_fire_1 : _GEN_2633) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_38) ? _GEN_2633 : dmem_req_fire_1;
    s1_executing_loads_20 <= will_fire_load_incoming_1_will_fire ? (_GEN_217 ? dmem_req_fire_1 : _GEN_2634) : will_fire_load_retry_1_will_fire ? (_GEN_121 ? dmem_req_fire_1 : _GEN_2634) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_39) ? _GEN_2634 : dmem_req_fire_1;
    s1_executing_loads_21 <= will_fire_load_incoming_1_will_fire ? (_GEN_219 ? dmem_req_fire_1 : _GEN_2635) : will_fire_load_retry_1_will_fire ? (_GEN_123 ? dmem_req_fire_1 : _GEN_2635) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_40) ? _GEN_2635 : dmem_req_fire_1;
    s1_executing_loads_22 <= will_fire_load_incoming_1_will_fire ? (_GEN_221 ? dmem_req_fire_1 : _GEN_2636) : will_fire_load_retry_1_will_fire ? (_GEN_125 ? dmem_req_fire_1 : _GEN_2636) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_41) ? _GEN_2636 : dmem_req_fire_1;
    s1_executing_loads_23 <= will_fire_load_incoming_1_will_fire ? (_GEN_223 ? dmem_req_fire_1 : _GEN_2637) : will_fire_load_retry_1_will_fire ? (_GEN_127 ? dmem_req_fire_1 : _GEN_2637) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_42) ? _GEN_2637 : dmem_req_fire_1;
    s1_executing_loads_24 <= will_fire_load_incoming_1_will_fire ? (_GEN_225 ? dmem_req_fire_1 : _GEN_2638) : will_fire_load_retry_1_will_fire ? (_GEN_129 ? dmem_req_fire_1 : _GEN_2638) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_43) ? _GEN_2638 : dmem_req_fire_1;
    s1_executing_loads_25 <= will_fire_load_incoming_1_will_fire ? (_GEN_227 ? dmem_req_fire_1 : _GEN_2639) : will_fire_load_retry_1_will_fire ? (_GEN_131 ? dmem_req_fire_1 : _GEN_2639) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_44) ? _GEN_2639 : dmem_req_fire_1;
    s1_executing_loads_26 <= will_fire_load_incoming_1_will_fire ? (_GEN_229 ? dmem_req_fire_1 : _GEN_2640) : will_fire_load_retry_1_will_fire ? (_GEN_133 ? dmem_req_fire_1 : _GEN_2640) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_45) ? _GEN_2640 : dmem_req_fire_1;
    s1_executing_loads_27 <= will_fire_load_incoming_1_will_fire ? (_GEN_231 ? dmem_req_fire_1 : _GEN_2641) : will_fire_load_retry_1_will_fire ? (_GEN_135 ? dmem_req_fire_1 : _GEN_2641) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_46) ? _GEN_2641 : dmem_req_fire_1;
    s1_executing_loads_28 <= will_fire_load_incoming_1_will_fire ? (_GEN_233 ? dmem_req_fire_1 : _GEN_2642) : will_fire_load_retry_1_will_fire ? (_GEN_137 ? dmem_req_fire_1 : _GEN_2642) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_47) ? _GEN_2642 : dmem_req_fire_1;
    s1_executing_loads_29 <= will_fire_load_incoming_1_will_fire ? (_GEN_235 ? dmem_req_fire_1 : _GEN_2643) : will_fire_load_retry_1_will_fire ? (_GEN_139 ? dmem_req_fire_1 : _GEN_2643) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_48) ? _GEN_2643 : dmem_req_fire_1;
    s1_executing_loads_30 <= will_fire_load_incoming_1_will_fire ? (_GEN_237 ? dmem_req_fire_1 : _GEN_2644) : will_fire_load_retry_1_will_fire ? (_GEN_141 ? dmem_req_fire_1 : _GEN_2644) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & _GEN_49) ? _GEN_2644 : dmem_req_fire_1;
    s1_executing_loads_31 <= will_fire_load_incoming_1_will_fire ? ((&_mem_incoming_uop_WIRE_1_ldq_idx) ? dmem_req_fire_1 : _GEN_2645) : will_fire_load_retry_1_will_fire ? ((&ldq_retry_idx) ? dmem_req_fire_1 : _GEN_2645) : will_fire_store_commit_1_will_fire | ~(will_fire_load_wakeup_1_will_fire & (&ldq_wakeup_idx)) ? _GEN_2645 : dmem_req_fire_1;
    wb_forward_valid_0 <= casez_tmp_455 & (io_core_brupdate_b1_mispredict_mask & (do_st_search_0 ? (_lcam_stq_idx_T ? mem_stq_incoming_e_0_bits_uop_br_mask : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_br_mask : 20'h0) : do_ld_search_0 ? (fired_load_incoming_REG ? mem_ldq_incoming_e_0_bits_uop_br_mask : fired_load_retry_REG ? mem_ldq_retry_e_bits_uop_br_mask : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_uop_br_mask : 20'h0) : 20'h0)) == 20'h0 & ~io_core_exception & ~REG_2;
    wb_forward_valid_1 <= casez_tmp_456 & (io_core_brupdate_b1_mispredict_mask & (do_st_search_1 ? (_lcam_stq_idx_T_3 ? mem_stq_incoming_e_1_bits_uop_br_mask : fired_sta_retry_REG_1 ? mem_stq_retry_e_bits_uop_br_mask : 20'h0) : do_ld_search_1 ? (fired_load_incoming_REG_1 ? mem_ldq_incoming_e_1_bits_uop_br_mask : fired_load_retry_REG_1 ? mem_ldq_retry_e_bits_uop_br_mask : fired_load_wakeup_REG_1 ? mem_ldq_wakeup_e_bits_uop_br_mask : 20'h0) : 20'h0)) == 20'h0 & ~io_core_exception & ~REG_3;
    wb_forward_ldq_idx_0 <= lcam_ldq_idx_0;
    wb_forward_ldq_idx_1 <= lcam_ldq_idx_1;
    wb_forward_ld_addr_0 <= lcam_addr_0;
    wb_forward_ld_addr_1 <= lcam_addr_1;
    wb_forward_stq_idx_0 <= _forwarding_age_logic_0_io_forwarding_idx;
    wb_forward_stq_idx_1 <= _forwarding_age_logic_1_io_forwarding_idx;
    older_nacked_REG <= nacking_loads_0;
    io_dmem_s1_kill_0_REG <= dmem_req_fire_0;
    older_nacked_REG_1 <= nacking_loads_0;
    io_dmem_s1_kill_1_REG <= dmem_req_fire_1;
    older_nacked_REG_2 <= nacking_loads_1;
    io_dmem_s1_kill_0_REG_1 <= dmem_req_fire_0;
    older_nacked_REG_3 <= nacking_loads_1;
    io_dmem_s1_kill_1_REG_1 <= dmem_req_fire_1;
    older_nacked_REG_4 <= nacking_loads_2;
    io_dmem_s1_kill_0_REG_2 <= dmem_req_fire_0;
    older_nacked_REG_5 <= nacking_loads_2;
    io_dmem_s1_kill_1_REG_2 <= dmem_req_fire_1;
    older_nacked_REG_6 <= nacking_loads_3;
    io_dmem_s1_kill_0_REG_3 <= dmem_req_fire_0;
    older_nacked_REG_7 <= nacking_loads_3;
    io_dmem_s1_kill_1_REG_3 <= dmem_req_fire_1;
    older_nacked_REG_8 <= nacking_loads_4;
    io_dmem_s1_kill_0_REG_4 <= dmem_req_fire_0;
    older_nacked_REG_9 <= nacking_loads_4;
    io_dmem_s1_kill_1_REG_4 <= dmem_req_fire_1;
    older_nacked_REG_10 <= nacking_loads_5;
    io_dmem_s1_kill_0_REG_5 <= dmem_req_fire_0;
    older_nacked_REG_11 <= nacking_loads_5;
    io_dmem_s1_kill_1_REG_5 <= dmem_req_fire_1;
    older_nacked_REG_12 <= nacking_loads_6;
    io_dmem_s1_kill_0_REG_6 <= dmem_req_fire_0;
    older_nacked_REG_13 <= nacking_loads_6;
    io_dmem_s1_kill_1_REG_6 <= dmem_req_fire_1;
    older_nacked_REG_14 <= nacking_loads_7;
    io_dmem_s1_kill_0_REG_7 <= dmem_req_fire_0;
    older_nacked_REG_15 <= nacking_loads_7;
    io_dmem_s1_kill_1_REG_7 <= dmem_req_fire_1;
    older_nacked_REG_16 <= nacking_loads_8;
    io_dmem_s1_kill_0_REG_8 <= dmem_req_fire_0;
    older_nacked_REG_17 <= nacking_loads_8;
    io_dmem_s1_kill_1_REG_8 <= dmem_req_fire_1;
    older_nacked_REG_18 <= nacking_loads_9;
    io_dmem_s1_kill_0_REG_9 <= dmem_req_fire_0;
    older_nacked_REG_19 <= nacking_loads_9;
    io_dmem_s1_kill_1_REG_9 <= dmem_req_fire_1;
    older_nacked_REG_20 <= nacking_loads_10;
    io_dmem_s1_kill_0_REG_10 <= dmem_req_fire_0;
    older_nacked_REG_21 <= nacking_loads_10;
    io_dmem_s1_kill_1_REG_10 <= dmem_req_fire_1;
    older_nacked_REG_22 <= nacking_loads_11;
    io_dmem_s1_kill_0_REG_11 <= dmem_req_fire_0;
    older_nacked_REG_23 <= nacking_loads_11;
    io_dmem_s1_kill_1_REG_11 <= dmem_req_fire_1;
    older_nacked_REG_24 <= nacking_loads_12;
    io_dmem_s1_kill_0_REG_12 <= dmem_req_fire_0;
    older_nacked_REG_25 <= nacking_loads_12;
    io_dmem_s1_kill_1_REG_12 <= dmem_req_fire_1;
    older_nacked_REG_26 <= nacking_loads_13;
    io_dmem_s1_kill_0_REG_13 <= dmem_req_fire_0;
    older_nacked_REG_27 <= nacking_loads_13;
    io_dmem_s1_kill_1_REG_13 <= dmem_req_fire_1;
    older_nacked_REG_28 <= nacking_loads_14;
    io_dmem_s1_kill_0_REG_14 <= dmem_req_fire_0;
    older_nacked_REG_29 <= nacking_loads_14;
    io_dmem_s1_kill_1_REG_14 <= dmem_req_fire_1;
    older_nacked_REG_30 <= nacking_loads_15;
    io_dmem_s1_kill_0_REG_15 <= dmem_req_fire_0;
    older_nacked_REG_31 <= nacking_loads_15;
    io_dmem_s1_kill_1_REG_15 <= dmem_req_fire_1;
    older_nacked_REG_32 <= nacking_loads_16;
    io_dmem_s1_kill_0_REG_16 <= dmem_req_fire_0;
    older_nacked_REG_33 <= nacking_loads_16;
    io_dmem_s1_kill_1_REG_16 <= dmem_req_fire_1;
    older_nacked_REG_34 <= nacking_loads_17;
    io_dmem_s1_kill_0_REG_17 <= dmem_req_fire_0;
    older_nacked_REG_35 <= nacking_loads_17;
    io_dmem_s1_kill_1_REG_17 <= dmem_req_fire_1;
    older_nacked_REG_36 <= nacking_loads_18;
    io_dmem_s1_kill_0_REG_18 <= dmem_req_fire_0;
    older_nacked_REG_37 <= nacking_loads_18;
    io_dmem_s1_kill_1_REG_18 <= dmem_req_fire_1;
    older_nacked_REG_38 <= nacking_loads_19;
    io_dmem_s1_kill_0_REG_19 <= dmem_req_fire_0;
    older_nacked_REG_39 <= nacking_loads_19;
    io_dmem_s1_kill_1_REG_19 <= dmem_req_fire_1;
    older_nacked_REG_40 <= nacking_loads_20;
    io_dmem_s1_kill_0_REG_20 <= dmem_req_fire_0;
    older_nacked_REG_41 <= nacking_loads_20;
    io_dmem_s1_kill_1_REG_20 <= dmem_req_fire_1;
    older_nacked_REG_42 <= nacking_loads_21;
    io_dmem_s1_kill_0_REG_21 <= dmem_req_fire_0;
    older_nacked_REG_43 <= nacking_loads_21;
    io_dmem_s1_kill_1_REG_21 <= dmem_req_fire_1;
    older_nacked_REG_44 <= nacking_loads_22;
    io_dmem_s1_kill_0_REG_22 <= dmem_req_fire_0;
    older_nacked_REG_45 <= nacking_loads_22;
    io_dmem_s1_kill_1_REG_22 <= dmem_req_fire_1;
    older_nacked_REG_46 <= nacking_loads_23;
    io_dmem_s1_kill_0_REG_23 <= dmem_req_fire_0;
    older_nacked_REG_47 <= nacking_loads_23;
    io_dmem_s1_kill_1_REG_23 <= dmem_req_fire_1;
    older_nacked_REG_48 <= nacking_loads_24;
    io_dmem_s1_kill_0_REG_24 <= dmem_req_fire_0;
    older_nacked_REG_49 <= nacking_loads_24;
    io_dmem_s1_kill_1_REG_24 <= dmem_req_fire_1;
    older_nacked_REG_50 <= nacking_loads_25;
    io_dmem_s1_kill_0_REG_25 <= dmem_req_fire_0;
    older_nacked_REG_51 <= nacking_loads_25;
    io_dmem_s1_kill_1_REG_25 <= dmem_req_fire_1;
    older_nacked_REG_52 <= nacking_loads_26;
    io_dmem_s1_kill_0_REG_26 <= dmem_req_fire_0;
    older_nacked_REG_53 <= nacking_loads_26;
    io_dmem_s1_kill_1_REG_26 <= dmem_req_fire_1;
    older_nacked_REG_54 <= nacking_loads_27;
    io_dmem_s1_kill_0_REG_27 <= dmem_req_fire_0;
    older_nacked_REG_55 <= nacking_loads_27;
    io_dmem_s1_kill_1_REG_27 <= dmem_req_fire_1;
    older_nacked_REG_56 <= nacking_loads_28;
    io_dmem_s1_kill_0_REG_28 <= dmem_req_fire_0;
    older_nacked_REG_57 <= nacking_loads_28;
    io_dmem_s1_kill_1_REG_28 <= dmem_req_fire_1;
    older_nacked_REG_58 <= nacking_loads_29;
    io_dmem_s1_kill_0_REG_29 <= dmem_req_fire_0;
    older_nacked_REG_59 <= nacking_loads_29;
    io_dmem_s1_kill_1_REG_29 <= dmem_req_fire_1;
    older_nacked_REG_60 <= nacking_loads_30;
    io_dmem_s1_kill_0_REG_30 <= dmem_req_fire_0;
    older_nacked_REG_61 <= nacking_loads_30;
    io_dmem_s1_kill_1_REG_30 <= dmem_req_fire_1;
    older_nacked_REG_62 <= nacking_loads_31;
    io_dmem_s1_kill_0_REG_31 <= dmem_req_fire_0;
    older_nacked_REG_63 <= nacking_loads_31;
    io_dmem_s1_kill_1_REG_31 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_32 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_33 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_34 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_32 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_33 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_34 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_35 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_36 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_37 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_35 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_36 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_37 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_38 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_39 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_40 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_38 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_39 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_40 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_41 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_42 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_43 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_41 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_42 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_43 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_44 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_45 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_46 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_44 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_45 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_46 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_47 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_48 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_49 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_47 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_48 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_49 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_50 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_51 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_52 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_50 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_51 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_52 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_53 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_54 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_55 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_53 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_54 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_55 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_56 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_57 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_58 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_56 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_57 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_58 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_59 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_60 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_61 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_59 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_60 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_61 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_62 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_63 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_64 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_62 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_63 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_64 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_65 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_66 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_67 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_65 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_66 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_67 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_68 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_69 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_70 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_68 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_69 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_70 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_71 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_72 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_73 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_71 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_72 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_73 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_74 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_75 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_76 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_74 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_75 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_76 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_77 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_78 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_79 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_77 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_78 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_79 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_80 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_81 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_82 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_80 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_81 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_82 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_83 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_84 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_85 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_83 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_84 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_85 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_86 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_87 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_88 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_86 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_87 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_88 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_89 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_90 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_91 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_89 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_90 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_91 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_92 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_93 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_94 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_92 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_93 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_94 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_95 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_96 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_97 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_95 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_96 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_97 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_98 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_99 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_100 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_98 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_99 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_100 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_101 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_102 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_103 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_101 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_102 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_103 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_104 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_105 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_106 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_104 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_105 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_106 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_107 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_108 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_109 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_107 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_108 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_109 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_110 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_111 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_112 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_110 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_111 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_112 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_113 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_114 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_115 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_113 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_114 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_115 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_116 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_117 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_118 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_116 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_117 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_118 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_119 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_120 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_121 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_119 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_120 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_121 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_122 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_123 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_124 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_122 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_123 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_124 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_125 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_126 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_127 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_125 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_126 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_127 <= dmem_req_fire_1;
    REG_2 <= io_core_exception;
    REG_3 <= io_core_exception;
    r_xcpt_uop_br_mask <= xcpt_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    r_xcpt_uop_rob_idx <= use_mem_xcpt ? mem_xcpt_uop_rob_idx : casez_tmp_458;
    r_xcpt_cause <= use_mem_xcpt ? {1'h0, _GEN_2550 ? mem_xcpt_causes_1 : mem_xcpt_causes_0} : 5'h10;
    r_xcpt_badvaddr <= _GEN_2550 ? mem_xcpt_vaddrs_1 : mem_xcpt_vaddrs_0;
    io_core_ld_miss_REG <= _io_core_spec_ld_wakeup_0_valid_output | _io_core_spec_ld_wakeup_1_valid_output;
    spec_ld_succeed_REG <= _io_core_spec_ld_wakeup_0_valid_output;
    spec_ld_succeed_REG_1 <= mem_incoming_uop_0_ldq_idx;
    spec_ld_succeed_REG_2 <= _io_core_spec_ld_wakeup_1_valid_output;
    spec_ld_succeed_REG_3 <= mem_incoming_uop_1_ldq_idx;
    if (reset) begin
      hella_state <= 3'h0;
      live_store_mask <= 32'h0;
      clr_bsy_valid_0 <= 1'h0;
      clr_bsy_valid_1 <= 1'h0;
      stdf_clr_bsy_valid <= 1'h0;
      r_xcpt_valid <= 1'h0;
    end
    else begin
      hella_state <= casez_tmp_547;
      live_store_mask <= ({32{dis_st_val_3}} & 32'h1 << _GEN_14 | _GEN_2166) & ~{stq_31_valid & (|_GEN_1542), stq_30_valid & (|_GEN_1541), stq_29_valid & (|_GEN_1540), stq_28_valid & (|_GEN_1539), stq_27_valid & (|_GEN_1538), stq_26_valid & (|_GEN_1537), stq_25_valid & (|_GEN_1536), stq_24_valid & (|_GEN_1535), stq_23_valid & (|_GEN_1534), stq_22_valid & (|_GEN_1533), stq_21_valid & (|_GEN_1532), stq_20_valid & (|_GEN_1531), stq_19_valid & (|_GEN_1530), stq_18_valid & (|_GEN_1529), stq_17_valid & (|_GEN_1528), stq_16_valid & (|_GEN_1527), stq_15_valid & (|_GEN_1526), stq_14_valid & (|_GEN_1525), stq_13_valid & (|_GEN_1524), stq_12_valid & (|_GEN_1523), stq_11_valid & (|_GEN_1522), stq_10_valid & (|_GEN_1521), stq_9_valid & (|_GEN_1520), stq_8_valid & (|_GEN_1519), stq_7_valid & (|_GEN_1518), stq_6_valid & (|_GEN_1517), stq_5_valid & (|_GEN_1516), stq_4_valid & (|_GEN_1515), stq_3_valid & (|_GEN_1514), stq_2_valid & (|_GEN_1513), stq_1_valid & (|_GEN_1512), stq_0_valid & (|_GEN_1511)} & ~{_GEN_5749 & ~reset & _GEN_5813, _GEN_5749 & ~reset & _GEN_5811, _GEN_5749 & ~reset & _GEN_5809, _GEN_5749 & ~reset & _GEN_5807, _GEN_5749 & ~reset & _GEN_5805, _GEN_5749 & ~reset & _GEN_5803, _GEN_5749 & ~reset & _GEN_5801, _GEN_5749 & ~reset & _GEN_5799, _GEN_5749 & ~reset & _GEN_5797, _GEN_5749 & ~reset & _GEN_5795, _GEN_5749 & ~reset & _GEN_5793, _GEN_5749 & ~reset & _GEN_5791, _GEN_5749 & ~reset & _GEN_5789, _GEN_5749 & ~reset & _GEN_5787, _GEN_5749 & ~reset & _GEN_5785, _GEN_5749 & ~reset & _GEN_5783, _GEN_5749 & ~reset & _GEN_5781, _GEN_5749 & ~reset & _GEN_5779, _GEN_5749 & ~reset & _GEN_5777, _GEN_5749 & ~reset & _GEN_5775, _GEN_5749 & ~reset & _GEN_5773, _GEN_5749 & ~reset & _GEN_5771, _GEN_5749 & ~reset & _GEN_5769, _GEN_5749 & ~reset & _GEN_5767, _GEN_5749 & ~reset & _GEN_5765, _GEN_5749 & ~reset & _GEN_5763, _GEN_5749 & ~reset & _GEN_5761, _GEN_5749 & ~reset & _GEN_5759, _GEN_5749 & ~reset & _GEN_5757, _GEN_5749 & ~reset & _GEN_5755, _GEN_5749 & ~reset & _GEN_5753, _GEN_5749 & ~reset & _GEN_5751};
      clr_bsy_valid_0 <= fired_stad_incoming_REG ? mem_stq_incoming_e_0_valid & ~mem_tlb_miss_0 & ~mem_stq_incoming_e_0_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_0_bits_uop_br_mask) == 20'h0 : fired_sta_incoming_REG ? mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_data_valid & ~mem_tlb_miss_0 & ~mem_stq_incoming_e_0_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_0_bits_uop_br_mask) == 20'h0 : fired_std_incoming_REG ? mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_addr_valid & ~mem_stq_incoming_e_0_bits_addr_is_virtual & ~mem_stq_incoming_e_0_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_0_bits_uop_br_mask) == 20'h0 : fired_sfence_0 | fired_sta_retry_REG & mem_stq_retry_e_valid & mem_stq_retry_e_bits_data_valid & ~mem_tlb_miss_0 & ~mem_stq_retry_e_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_retry_e_bits_uop_br_mask) == 20'h0;
      clr_bsy_valid_1 <= fired_stad_incoming_REG_1 ? mem_stq_incoming_e_1_valid & ~mem_tlb_miss_1 & ~mem_stq_incoming_e_1_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_1_bits_uop_br_mask) == 20'h0 : fired_sta_incoming_REG_1 ? mem_stq_incoming_e_1_valid & mem_stq_incoming_e_1_bits_data_valid & ~mem_tlb_miss_1 & ~mem_stq_incoming_e_1_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_1_bits_uop_br_mask) == 20'h0 : fired_std_incoming_REG_1 ? mem_stq_incoming_e_1_valid & mem_stq_incoming_e_1_bits_addr_valid & ~mem_stq_incoming_e_1_bits_addr_is_virtual & ~mem_stq_incoming_e_1_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_1_bits_uop_br_mask) == 20'h0 : ~fired_sfence_1 & fired_sta_retry_REG_1 & mem_stq_retry_e_valid & mem_stq_retry_e_bits_data_valid & ~mem_tlb_miss_1 & ~mem_stq_retry_e_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_retry_e_bits_uop_br_mask) == 20'h0;
      stdf_clr_bsy_valid <= fired_stdf_incoming & casez_tmp_383 & casez_tmp_385 & ~casez_tmp_386 & ~casez_tmp_384 & (io_core_brupdate_b1_mispredict_mask & mem_stdf_uop_br_mask) == 20'h0;
      r_xcpt_valid <= (ld_xcpt_valid | mem_xcpt_valid) & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & xcpt_uop_br_mask) == 20'h0;
    end
  end // always @(posedge)
  NBDTLB dtlb (
    .clock                        (clock),
    .reset                        (reset),
    .io_req_0_valid               (~_will_fire_store_commit_0_T_2),
    .io_req_0_bits_vaddr          (exe_tlb_vaddr_0),
    .io_req_0_bits_passthrough    (will_fire_hella_incoming_0_will_fire),
    .io_req_0_bits_size           (_exe_cmd_T | will_fire_sta_incoming_0_will_fire | will_fire_sfence_0_will_fire | will_fire_load_retry_0_will_fire | will_fire_sta_retry_0_will_fire ? exe_tlb_uop_0_mem_size : {2{will_fire_hella_incoming_0_will_fire}}),
    .io_req_0_bits_cmd            (_exe_cmd_T | will_fire_sta_incoming_0_will_fire | will_fire_sfence_0_will_fire | will_fire_load_retry_0_will_fire | will_fire_sta_retry_0_will_fire ? exe_tlb_uop_0_mem_cmd : 5'h0),
    .io_req_1_valid               (~_will_fire_store_commit_1_T_2),
    .io_req_1_bits_vaddr          (exe_tlb_vaddr_1),
    .io_req_1_bits_passthrough    (will_fire_hella_incoming_1_will_fire),
    .io_req_1_bits_size           (_exe_cmd_T_7 | will_fire_sta_incoming_1_will_fire | will_fire_sfence_1_will_fire | will_fire_load_retry_1_will_fire | will_fire_sta_retry_1_will_fire ? exe_tlb_uop_1_mem_size : {2{will_fire_hella_incoming_1_will_fire}}),
    .io_req_1_bits_cmd            (_exe_cmd_T_7 | will_fire_sta_incoming_1_will_fire | will_fire_sfence_1_will_fire | will_fire_load_retry_1_will_fire | will_fire_sta_retry_1_will_fire ? exe_tlb_uop_1_mem_cmd : 5'h0),
    .io_miss_rdy                  (_dtlb_io_miss_rdy),
    .io_resp_0_miss               (_dtlb_io_resp_0_miss),
    .io_resp_0_paddr              (_dtlb_io_resp_0_paddr),
    .io_resp_0_pf_ld              (_dtlb_io_resp_0_pf_ld),
    .io_resp_0_pf_st              (_dtlb_io_resp_0_pf_st),
    .io_resp_0_ae_ld              (_dtlb_io_resp_0_ae_ld),
    .io_resp_0_ae_st              (_dtlb_io_resp_0_ae_st),
    .io_resp_0_cacheable          (_dtlb_io_resp_0_cacheable),
    .io_resp_1_miss               (_dtlb_io_resp_1_miss),
    .io_resp_1_paddr              (_dtlb_io_resp_1_paddr),
    .io_resp_1_pf_ld              (_dtlb_io_resp_1_pf_ld),
    .io_resp_1_pf_st              (_dtlb_io_resp_1_pf_st),
    .io_resp_1_ae_ld              (_dtlb_io_resp_1_ae_ld),
    .io_resp_1_ae_st              (_dtlb_io_resp_1_ae_st),
    .io_resp_1_ma_ld              (_dtlb_io_resp_1_ma_ld),
    .io_resp_1_ma_st              (_dtlb_io_resp_1_ma_st),
    .io_resp_1_cacheable          (_dtlb_io_resp_1_cacheable),
    .io_sfence_valid              (will_fire_sfence_1_will_fire ? exe_req_1_bits_sfence_valid : will_fire_sfence_0_will_fire & exe_req_0_bits_sfence_valid),
    .io_sfence_bits_rs1           (will_fire_sfence_1_will_fire ? (_GEN_17 ? io_core_exe_1_req_bits_sfence_bits_rs1 : io_core_exe_0_req_bits_sfence_bits_rs1) : will_fire_sfence_0_will_fire & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_bits_rs1 : io_core_exe_0_req_bits_sfence_bits_rs1)),
    .io_sfence_bits_rs2           (will_fire_sfence_1_will_fire ? (_GEN_17 ? io_core_exe_1_req_bits_sfence_bits_rs2 : io_core_exe_0_req_bits_sfence_bits_rs2) : will_fire_sfence_0_will_fire & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_bits_rs2 : io_core_exe_0_req_bits_sfence_bits_rs2)),
    .io_sfence_bits_addr          (will_fire_sfence_1_will_fire ? exe_req_1_bits_sfence_bits_addr : will_fire_sfence_0_will_fire ? exe_req_0_bits_sfence_bits_addr : 39'h0),
    .io_ptw_req_ready             (io_ptw_req_ready),
    .io_ptw_req_valid             (io_ptw_req_valid),
    .io_ptw_req_bits_valid        (io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr    (io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid            (io_ptw_resp_valid),
    .io_ptw_resp_bits_ae_final    (io_ptw_resp_bits_ae_final),
    .io_ptw_resp_bits_pte_ppn     (io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d       (io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a       (io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g       (io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u       (io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x       (io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w       (io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r       (io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v       (io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level       (io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous (io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode             (io_ptw_ptbr_mode),
    .io_ptw_status_dprv           (io_ptw_status_dprv),
    .io_ptw_status_mxr            (io_ptw_status_mxr),
    .io_ptw_status_sum            (io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l           (io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a           (io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x           (io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w           (io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r           (io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr            (io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask            (io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l           (io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a           (io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x           (io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w           (io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r           (io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr            (io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask            (io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l           (io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a           (io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x           (io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w           (io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r           (io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr            (io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask            (io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l           (io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a           (io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x           (io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w           (io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r           (io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr            (io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask            (io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l           (io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a           (io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x           (io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w           (io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r           (io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr            (io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask            (io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l           (io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a           (io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x           (io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w           (io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r           (io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr            (io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask            (io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l           (io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a           (io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x           (io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w           (io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r           (io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr            (io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask            (io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l           (io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a           (io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x           (io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w           (io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r           (io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr            (io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask            (io_ptw_pmp_7_mask),
    .io_kill                      (will_fire_hella_incoming_0_will_fire & io_hellacache_s1_kill | will_fire_hella_incoming_1_will_fire & io_hellacache_s1_kill)
  );
  ForwardingAgeLogic forwarding_age_logic_0 (
    .io_addr_matches    ({_GEN_1421 & (_GEN_1423 | _GEN_1424 | _GEN_1425), _GEN_1410 & (_GEN_1412 | _GEN_1413 | _GEN_1414), _GEN_1399 & (_GEN_1401 | _GEN_1402 | _GEN_1403), _GEN_1388 & (_GEN_1390 | _GEN_1391 | _GEN_1392), _GEN_1377 & (_GEN_1379 | _GEN_1380 | _GEN_1381), _GEN_1366 & (_GEN_1368 | _GEN_1369 | _GEN_1370), _GEN_1355 & (_GEN_1357 | _GEN_1358 | _GEN_1359), _GEN_1344 & (_GEN_1346 | _GEN_1347 | _GEN_1348), _GEN_1333 & (_GEN_1335 | _GEN_1336 | _GEN_1337), _GEN_1322 & (_GEN_1324 | _GEN_1325 | _GEN_1326), _GEN_1311 & (_GEN_1313 | _GEN_1314 | _GEN_1315), _GEN_1300 & (_GEN_1302 | _GEN_1303 | _GEN_1304), _GEN_1289 & (_GEN_1291 | _GEN_1292 | _GEN_1293), _GEN_1278 & (_GEN_1280 | _GEN_1281 | _GEN_1282), _GEN_1267 & (_GEN_1269 | _GEN_1270 | _GEN_1271), _GEN_1256 & (_GEN_1258 | _GEN_1259 | _GEN_1260), _GEN_1245 & (_GEN_1247 | _GEN_1248 | _GEN_1249), _GEN_1234 & (_GEN_1236 | _GEN_1237 | _GEN_1238), _GEN_1223 & (_GEN_1225 | _GEN_1226 | _GEN_1227), _GEN_1212 & (_GEN_1214 | _GEN_1215 | _GEN_1216), _GEN_1201 & (_GEN_1203 | _GEN_1204 | _GEN_1205), _GEN_1190 & (_GEN_1192 | _GEN_1193 | _GEN_1194), _GEN_1179 & (_GEN_1181 | _GEN_1182 | _GEN_1183), _GEN_1168 & (_GEN_1170 | _GEN_1171 | _GEN_1172), _GEN_1157 & (_GEN_1159 | _GEN_1160 | _GEN_1161), _GEN_1146 & (_GEN_1148 | _GEN_1149 | _GEN_1150), _GEN_1135 & (_GEN_1137 | _GEN_1138 | _GEN_1139), _GEN_1124 & (_GEN_1126 | _GEN_1127 | _GEN_1128), _GEN_1113 & (_GEN_1115 | _GEN_1116 | _GEN_1117), _GEN_1102 & (_GEN_1104 | _GEN_1105 | _GEN_1106), _GEN_1091 & (_GEN_1093 | _GEN_1094 | _GEN_1095), _GEN_1080 & (_GEN_1082 | _GEN_1083 | _GEN_1084)}),
    .io_youngest_st_idx (do_st_search_0 ? (_lcam_stq_idx_T ? mem_stq_incoming_e_0_bits_uop_stq_idx : fired_sta_retry_REG ? mem_stq_retry_e_bits_uop_stq_idx : 5'h0) : do_ld_search_0 ? (fired_load_incoming_REG ? mem_ldq_incoming_e_0_bits_uop_stq_idx : fired_load_retry_REG ? mem_ldq_retry_e_bits_uop_stq_idx : fired_load_wakeup_REG ? mem_ldq_wakeup_e_bits_uop_stq_idx : 5'h0) : 5'h0),
    .io_forwarding_idx  (_forwarding_age_logic_0_io_forwarding_idx)
  );
  ForwardingAgeLogic forwarding_age_logic_1 (
    .io_addr_matches    ({_GEN_1426 & (_GEN_1428 | _GEN_1429 | _GEN_1425), _GEN_1416 & (_GEN_1418 | _GEN_1419 | _GEN_1414), _GEN_1405 & (_GEN_1407 | _GEN_1408 | _GEN_1403), _GEN_1394 & (_GEN_1396 | _GEN_1397 | _GEN_1392), _GEN_1383 & (_GEN_1385 | _GEN_1386 | _GEN_1381), _GEN_1372 & (_GEN_1374 | _GEN_1375 | _GEN_1370), _GEN_1361 & (_GEN_1363 | _GEN_1364 | _GEN_1359), _GEN_1350 & (_GEN_1352 | _GEN_1353 | _GEN_1348), _GEN_1339 & (_GEN_1341 | _GEN_1342 | _GEN_1337), _GEN_1328 & (_GEN_1330 | _GEN_1331 | _GEN_1326), _GEN_1317 & (_GEN_1319 | _GEN_1320 | _GEN_1315), _GEN_1306 & (_GEN_1308 | _GEN_1309 | _GEN_1304), _GEN_1295 & (_GEN_1297 | _GEN_1298 | _GEN_1293), _GEN_1284 & (_GEN_1286 | _GEN_1287 | _GEN_1282), _GEN_1273 & (_GEN_1275 | _GEN_1276 | _GEN_1271), _GEN_1262 & (_GEN_1264 | _GEN_1265 | _GEN_1260), _GEN_1251 & (_GEN_1253 | _GEN_1254 | _GEN_1249), _GEN_1240 & (_GEN_1242 | _GEN_1243 | _GEN_1238), _GEN_1229 & (_GEN_1231 | _GEN_1232 | _GEN_1227), _GEN_1218 & (_GEN_1220 | _GEN_1221 | _GEN_1216), _GEN_1207 & (_GEN_1209 | _GEN_1210 | _GEN_1205), _GEN_1196 & (_GEN_1198 | _GEN_1199 | _GEN_1194), _GEN_1185 & (_GEN_1187 | _GEN_1188 | _GEN_1183), _GEN_1174 & (_GEN_1176 | _GEN_1177 | _GEN_1172), _GEN_1163 & (_GEN_1165 | _GEN_1166 | _GEN_1161), _GEN_1152 & (_GEN_1154 | _GEN_1155 | _GEN_1150), _GEN_1141 & (_GEN_1143 | _GEN_1144 | _GEN_1139), _GEN_1130 & (_GEN_1132 | _GEN_1133 | _GEN_1128), _GEN_1119 & (_GEN_1121 | _GEN_1122 | _GEN_1117), _GEN_1108 & (_GEN_1110 | _GEN_1111 | _GEN_1106), _GEN_1097 & (_GEN_1099 | _GEN_1100 | _GEN_1095), _GEN_1086 & (_GEN_1088 | _GEN_1089 | _GEN_1084)}),
    .io_youngest_st_idx (do_st_search_1 ? (_lcam_stq_idx_T_3 ? mem_stq_incoming_e_1_bits_uop_stq_idx : fired_sta_retry_REG_1 ? mem_stq_retry_e_bits_uop_stq_idx : 5'h0) : do_ld_search_1 ? (fired_load_incoming_REG_1 ? mem_ldq_incoming_e_1_bits_uop_stq_idx : fired_load_retry_REG_1 ? mem_ldq_retry_e_bits_uop_stq_idx : fired_load_wakeup_REG_1 ? mem_ldq_wakeup_e_bits_uop_stq_idx : 5'h0) : 5'h0),
    .io_forwarding_idx  (_forwarding_age_logic_1_io_forwarding_idx)
  );
  assign io_core_exe_0_iresp_valid = _io_core_exe_0_iresp_valid_output;
  assign io_core_exe_0_iresp_bits_uop_rob_idx = _GEN_1470 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_462 : casez_tmp_471) : casez_tmp_479;
  assign io_core_exe_0_iresp_bits_uop_pdst = _GEN_1470 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_465 : casez_tmp_473) : casez_tmp_482;
  assign io_core_exe_0_iresp_bits_uop_is_amo = _GEN_1470 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_467 : casez_tmp_474) : casez_tmp_485;
  assign io_core_exe_0_iresp_bits_uop_uses_stq = _GEN_1470 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_468 : casez_tmp_475) : casez_tmp_486;
  assign io_core_exe_0_iresp_bits_uop_dst_rtype = _GEN_1470 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_469 : casez_tmp_476) : casez_tmp_487;
  assign io_core_exe_0_iresp_bits_data = _GEN_1470 ? io_dmem_resp_0_bits_data : {_ldq_bits_debug_wb_data_T_19 ? {56{casez_tmp_484 & io_core_exe_0_iresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_10 ? {48{casez_tmp_484 & io_core_exe_0_iresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_1 ? {32{casez_tmp_484 & io_core_exe_0_iresp_bits_data_zeroed[31]}} : casez_tmp_492[63:32], io_core_exe_0_iresp_bits_data_zeroed[31:16]}, io_core_exe_0_iresp_bits_data_zeroed_1[15:8]}, io_core_exe_0_iresp_bits_data_zeroed_2};
  assign io_core_exe_0_fresp_valid = _io_core_exe_0_fresp_valid_output;
  assign io_core_exe_0_fresp_bits_uop_uopc = _GEN_1470 ? casez_tmp_460 : casez_tmp_477;
  assign io_core_exe_0_fresp_bits_uop_br_mask = _GEN_1470 ? casez_tmp_461 : casez_tmp_478;
  assign io_core_exe_0_fresp_bits_uop_rob_idx = _GEN_1470 ? casez_tmp_462 : casez_tmp_479;
  assign io_core_exe_0_fresp_bits_uop_stq_idx = _GEN_1470 ? casez_tmp_464 : casez_tmp_481;
  assign io_core_exe_0_fresp_bits_uop_pdst = _GEN_1470 ? casez_tmp_465 : casez_tmp_482;
  assign io_core_exe_0_fresp_bits_uop_mem_size = _GEN_1470 ? casez_tmp_466 : casez_tmp_483;
  assign io_core_exe_0_fresp_bits_uop_is_amo = _GEN_1470 ? casez_tmp_467 : casez_tmp_485;
  assign io_core_exe_0_fresp_bits_uop_uses_stq = _GEN_1470 ? casez_tmp_468 : casez_tmp_486;
  assign io_core_exe_0_fresp_bits_uop_dst_rtype = _GEN_1470 ? casez_tmp_469 : casez_tmp_487;
  assign io_core_exe_0_fresp_bits_uop_fp_val = _GEN_1470 ? casez_tmp_470 : casez_tmp_488;
  assign io_core_exe_0_fresp_bits_data = {1'h0, _GEN_1470 ? io_dmem_resp_0_bits_data : {_ldq_bits_debug_wb_data_T_19 ? {56{casez_tmp_484 & io_core_exe_0_fresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_10 ? {48{casez_tmp_484 & io_core_exe_0_fresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_1 ? {32{casez_tmp_484 & io_core_exe_0_fresp_bits_data_zeroed[31]}} : casez_tmp_492[63:32], io_core_exe_0_fresp_bits_data_zeroed[31:16]}, io_core_exe_0_fresp_bits_data_zeroed_1[15:8]}, io_core_exe_0_fresp_bits_data_zeroed_2}};
  assign io_core_exe_1_iresp_valid = _io_core_exe_1_iresp_valid_output;
  assign io_core_exe_1_iresp_bits_uop_rob_idx = _GEN_1510 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_496 : casez_tmp_505) : casez_tmp_513;
  assign io_core_exe_1_iresp_bits_uop_pdst = _GEN_1510 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_499 : casez_tmp_507) : casez_tmp_516;
  assign io_core_exe_1_iresp_bits_uop_is_amo = _GEN_1510 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_501 : casez_tmp_508) : casez_tmp_519;
  assign io_core_exe_1_iresp_bits_uop_uses_stq = _GEN_1510 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_502 : casez_tmp_509) : casez_tmp_520;
  assign io_core_exe_1_iresp_bits_uop_dst_rtype = _GEN_1510 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_503 : casez_tmp_510) : casez_tmp_521;
  assign io_core_exe_1_iresp_bits_data = _GEN_1510 ? io_dmem_resp_1_bits_data : {_ldq_bits_debug_wb_data_T_46 ? {56{casez_tmp_518 & io_core_exe_1_iresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_37 ? {48{casez_tmp_518 & io_core_exe_1_iresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_28 ? {32{casez_tmp_518 & io_core_exe_1_iresp_bits_data_zeroed[31]}} : casez_tmp_526[63:32], io_core_exe_1_iresp_bits_data_zeroed[31:16]}, io_core_exe_1_iresp_bits_data_zeroed_1[15:8]}, io_core_exe_1_iresp_bits_data_zeroed_2};
  assign io_core_exe_1_fresp_valid = _io_core_exe_1_fresp_valid_output;
  assign io_core_exe_1_fresp_bits_uop_uopc = _GEN_1510 ? casez_tmp_494 : casez_tmp_511;
  assign io_core_exe_1_fresp_bits_uop_br_mask = _GEN_1510 ? casez_tmp_495 : casez_tmp_512;
  assign io_core_exe_1_fresp_bits_uop_rob_idx = _GEN_1510 ? casez_tmp_496 : casez_tmp_513;
  assign io_core_exe_1_fresp_bits_uop_stq_idx = _GEN_1510 ? casez_tmp_498 : casez_tmp_515;
  assign io_core_exe_1_fresp_bits_uop_pdst = _GEN_1510 ? casez_tmp_499 : casez_tmp_516;
  assign io_core_exe_1_fresp_bits_uop_mem_size = _GEN_1510 ? casez_tmp_500 : casez_tmp_517;
  assign io_core_exe_1_fresp_bits_uop_is_amo = _GEN_1510 ? casez_tmp_501 : casez_tmp_519;
  assign io_core_exe_1_fresp_bits_uop_uses_stq = _GEN_1510 ? casez_tmp_502 : casez_tmp_520;
  assign io_core_exe_1_fresp_bits_uop_dst_rtype = _GEN_1510 ? casez_tmp_503 : casez_tmp_521;
  assign io_core_exe_1_fresp_bits_uop_fp_val = _GEN_1510 ? casez_tmp_504 : casez_tmp_522;
  assign io_core_exe_1_fresp_bits_data = {1'h0, _GEN_1510 ? io_dmem_resp_1_bits_data : {_ldq_bits_debug_wb_data_T_46 ? {56{casez_tmp_518 & io_core_exe_1_fresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_37 ? {48{casez_tmp_518 & io_core_exe_1_fresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_28 ? {32{casez_tmp_518 & io_core_exe_1_fresp_bits_data_zeroed[31]}} : casez_tmp_526[63:32], io_core_exe_1_fresp_bits_data_zeroed[31:16]}, io_core_exe_1_fresp_bits_data_zeroed_1[15:8]}, io_core_exe_1_fresp_bits_data_zeroed_2}};
  assign io_core_dis_ldq_idx_0 = ldq_tail;
  assign io_core_dis_ldq_idx_1 = _GEN_5;
  assign io_core_dis_ldq_idx_2 = _GEN_9;
  assign io_core_dis_ldq_idx_3 = _GEN_13;
  assign io_core_dis_stq_idx_0 = stq_tail;
  assign io_core_dis_stq_idx_1 = _GEN_6;
  assign io_core_dis_stq_idx_2 = _GEN_10;
  assign io_core_dis_stq_idx_3 = _GEN_14;
  assign io_core_ldq_full_0 = _GEN_3 == ldq_head;
  assign io_core_ldq_full_1 = _GEN_7 == ldq_head;
  assign io_core_ldq_full_2 = _GEN_11 == ldq_head;
  assign io_core_ldq_full_3 = _GEN_15 == ldq_head;
  assign io_core_stq_full_0 = _GEN_4 == stq_head;
  assign io_core_stq_full_1 = _GEN_8 == stq_head;
  assign io_core_stq_full_2 = _GEN_12 == stq_head;
  assign io_core_stq_full_3 = _GEN_16 == stq_head;
  assign io_core_fp_stdata_ready = _io_core_fp_stdata_ready_output;
  assign io_core_clr_bsy_0_valid = clr_bsy_valid_0 & (io_core_brupdate_b1_mispredict_mask & clr_bsy_brmask_0) == 20'h0 & ~io_core_exception & ~io_core_clr_bsy_0_valid_REG & ~io_core_clr_bsy_0_valid_REG_2;
  assign io_core_clr_bsy_0_bits = clr_bsy_rob_idx_0;
  assign io_core_clr_bsy_1_valid = clr_bsy_valid_1 & (io_core_brupdate_b1_mispredict_mask & clr_bsy_brmask_1) == 20'h0 & ~io_core_exception & ~io_core_clr_bsy_1_valid_REG & ~io_core_clr_bsy_1_valid_REG_2;
  assign io_core_clr_bsy_1_bits = clr_bsy_rob_idx_1;
  assign io_core_clr_bsy_2_valid = stdf_clr_bsy_valid & (io_core_brupdate_b1_mispredict_mask & stdf_clr_bsy_brmask) == 20'h0 & ~io_core_exception & ~io_core_clr_bsy_2_valid_REG & ~io_core_clr_bsy_2_valid_REG_2;
  assign io_core_clr_bsy_2_bits = stdf_clr_bsy_rob_idx;
  assign io_core_spec_ld_wakeup_0_valid = _io_core_spec_ld_wakeup_0_valid_output;
  assign io_core_spec_ld_wakeup_0_bits = mem_incoming_uop_0_pdst;
  assign io_core_spec_ld_wakeup_1_valid = _io_core_spec_ld_wakeup_1_valid_output;
  assign io_core_spec_ld_wakeup_1_bits = mem_incoming_uop_1_pdst;
  assign io_core_ld_miss = ~((~spec_ld_succeed_REG | _io_core_exe_0_iresp_valid_output & (_GEN_1470 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_463 : casez_tmp_472) : casez_tmp_480) == spec_ld_succeed_REG_1) & (~spec_ld_succeed_REG_2 | _io_core_exe_1_iresp_valid_output & (_GEN_1510 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_497 : casez_tmp_506) : casez_tmp_514) == spec_ld_succeed_REG_3)) & io_core_ld_miss_REG;
  assign io_core_fencei_rdy = ~(stq_0_valid | stq_1_valid | stq_2_valid | stq_3_valid | stq_4_valid | stq_5_valid | stq_6_valid | stq_7_valid | stq_8_valid | stq_9_valid | stq_10_valid | stq_11_valid | stq_12_valid | stq_13_valid | stq_14_valid | stq_15_valid | stq_16_valid | stq_17_valid | stq_18_valid | stq_19_valid | stq_20_valid | stq_21_valid | stq_22_valid | stq_23_valid | stq_24_valid | stq_25_valid | stq_26_valid | stq_27_valid | stq_28_valid | stq_29_valid | stq_30_valid | stq_31_valid) & io_dmem_ordered;
  assign io_core_lxcpt_valid = r_xcpt_valid & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & r_xcpt_uop_br_mask) == 20'h0;
  assign io_core_lxcpt_bits_uop_br_mask = r_xcpt_uop_br_mask;
  assign io_core_lxcpt_bits_uop_rob_idx = r_xcpt_uop_rob_idx;
  assign io_core_lxcpt_bits_cause = r_xcpt_cause;
  assign io_core_lxcpt_bits_badvaddr = r_xcpt_badvaddr;
  assign io_dmem_req_valid = _io_dmem_req_valid_output;
  assign io_dmem_req_bits_0_valid = dmem_req_0_valid;
  assign io_dmem_req_bits_0_bits_uop_uopc = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_uopc : io_core_exe_0_req_bits_uop_uopc) : will_fire_load_retry_0_will_fire ? casez_tmp_124 : will_fire_sta_retry_0_will_fire ? casez_tmp_210 : 7'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_0 : will_fire_load_wakeup_0_will_fire ? casez_tmp_294 : 7'h0;
  assign io_dmem_req_bits_0_bits_uop_inst = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_inst : io_core_exe_0_req_bits_uop_inst) : will_fire_load_retry_0_will_fire ? casez_tmp_125 : will_fire_sta_retry_0_will_fire ? casez_tmp_211 : 32'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_1 : will_fire_load_wakeup_0_will_fire ? casez_tmp_295 : 32'h0;
  assign io_dmem_req_bits_0_bits_uop_debug_inst = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_debug_inst : io_core_exe_0_req_bits_uop_debug_inst) : will_fire_load_retry_0_will_fire ? casez_tmp_126 : will_fire_sta_retry_0_will_fire ? casez_tmp_212 : 32'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_2 : will_fire_load_wakeup_0_will_fire ? casez_tmp_296 : 32'h0;
  assign io_dmem_req_bits_0_bits_uop_is_rvc = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_rvc : io_core_exe_0_req_bits_uop_is_rvc) : will_fire_load_retry_0_will_fire ? casez_tmp_127 : will_fire_sta_retry_0_will_fire & casez_tmp_213) : will_fire_store_commit_0_will_fire ? casez_tmp_3 : will_fire_load_wakeup_0_will_fire & casez_tmp_297;
  assign io_dmem_req_bits_0_bits_uop_debug_pc = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_debug_pc : io_core_exe_0_req_bits_uop_debug_pc) : will_fire_load_retry_0_will_fire ? casez_tmp_128 : will_fire_sta_retry_0_will_fire ? casez_tmp_214 : 40'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_4 : will_fire_load_wakeup_0_will_fire ? casez_tmp_298 : 40'h0;
  assign io_dmem_req_bits_0_bits_uop_iq_type = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_iq_type : io_core_exe_0_req_bits_uop_iq_type) : will_fire_load_retry_0_will_fire ? casez_tmp_129 : will_fire_sta_retry_0_will_fire ? casez_tmp_215 : 3'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_5 : will_fire_load_wakeup_0_will_fire ? casez_tmp_299 : 3'h0;
  assign io_dmem_req_bits_0_bits_uop_fu_code = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_fu_code : io_core_exe_0_req_bits_uop_fu_code) : will_fire_load_retry_0_will_fire ? casez_tmp_130 : will_fire_sta_retry_0_will_fire ? casez_tmp_216 : 10'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_6 : will_fire_load_wakeup_0_will_fire ? casez_tmp_300 : 10'h0;
  assign io_dmem_req_bits_0_bits_uop_ctrl_br_type = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_br_type : io_core_exe_0_req_bits_uop_ctrl_br_type) : will_fire_load_retry_0_will_fire ? casez_tmp_131 : will_fire_sta_retry_0_will_fire ? casez_tmp_217 : 4'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_7 : will_fire_load_wakeup_0_will_fire ? casez_tmp_301 : 4'h0;
  assign io_dmem_req_bits_0_bits_uop_ctrl_op1_sel = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_op1_sel : io_core_exe_0_req_bits_uop_ctrl_op1_sel) : will_fire_load_retry_0_will_fire ? casez_tmp_132 : will_fire_sta_retry_0_will_fire ? casez_tmp_218 : 2'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_8 : will_fire_load_wakeup_0_will_fire ? casez_tmp_302 : 2'h0;
  assign io_dmem_req_bits_0_bits_uop_ctrl_op2_sel = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_op2_sel : io_core_exe_0_req_bits_uop_ctrl_op2_sel) : will_fire_load_retry_0_will_fire ? casez_tmp_133 : will_fire_sta_retry_0_will_fire ? casez_tmp_219 : 3'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_9 : will_fire_load_wakeup_0_will_fire ? casez_tmp_303 : 3'h0;
  assign io_dmem_req_bits_0_bits_uop_ctrl_imm_sel = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_imm_sel : io_core_exe_0_req_bits_uop_ctrl_imm_sel) : will_fire_load_retry_0_will_fire ? casez_tmp_134 : will_fire_sta_retry_0_will_fire ? casez_tmp_220 : 3'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_10 : will_fire_load_wakeup_0_will_fire ? casez_tmp_304 : 3'h0;
  assign io_dmem_req_bits_0_bits_uop_ctrl_op_fcn = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_op_fcn : io_core_exe_0_req_bits_uop_ctrl_op_fcn) : will_fire_load_retry_0_will_fire ? casez_tmp_135 : will_fire_sta_retry_0_will_fire ? casez_tmp_221 : 4'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_11 : will_fire_load_wakeup_0_will_fire ? casez_tmp_305 : 4'h0;
  assign io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_fcn_dw : io_core_exe_0_req_bits_uop_ctrl_fcn_dw) : will_fire_load_retry_0_will_fire ? casez_tmp_136 : will_fire_sta_retry_0_will_fire & casez_tmp_222) : will_fire_store_commit_0_will_fire ? casez_tmp_12 : will_fire_load_wakeup_0_will_fire & casez_tmp_306;
  assign io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_csr_cmd : io_core_exe_0_req_bits_uop_ctrl_csr_cmd) : will_fire_load_retry_0_will_fire ? casez_tmp_137 : will_fire_sta_retry_0_will_fire ? casez_tmp_223 : 3'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_13 : will_fire_load_wakeup_0_will_fire ? casez_tmp_307 : 3'h0;
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_load = _GEN_275 ? exe_tlb_uop_0_ctrl_is_load : will_fire_store_commit_0_will_fire ? casez_tmp_14 : will_fire_load_wakeup_0_will_fire & casez_tmp_308;
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_sta = _GEN_275 ? exe_tlb_uop_0_ctrl_is_sta : will_fire_store_commit_0_will_fire ? casez_tmp_15 : will_fire_load_wakeup_0_will_fire & casez_tmp_309;
  assign io_dmem_req_bits_0_bits_uop_ctrl_is_std = _GEN_275 ? (_exe_tlb_uop_T_2 ? exe_req_0_bits_uop_ctrl_is_std : will_fire_load_retry_0_will_fire ? casez_tmp_140 : will_fire_sta_retry_0_will_fire & casez_tmp_226) : will_fire_store_commit_0_will_fire ? casez_tmp_16 : will_fire_load_wakeup_0_will_fire & casez_tmp_310;
  assign io_dmem_req_bits_0_bits_uop_iw_state = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_iw_state : io_core_exe_0_req_bits_uop_iw_state) : will_fire_load_retry_0_will_fire ? casez_tmp_141 : will_fire_sta_retry_0_will_fire ? casez_tmp_227 : 2'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_17 : will_fire_load_wakeup_0_will_fire ? casez_tmp_311 : 2'h0;
  assign io_dmem_req_bits_0_bits_uop_iw_p1_poisoned = _GEN_275 ? ~_exe_tlb_uop_T_2 & (will_fire_load_retry_0_will_fire ? casez_tmp_142 : will_fire_sta_retry_0_will_fire & casez_tmp_228) : will_fire_store_commit_0_will_fire ? casez_tmp_18 : will_fire_load_wakeup_0_will_fire & casez_tmp_312;
  assign io_dmem_req_bits_0_bits_uop_iw_p2_poisoned = _GEN_275 ? ~_exe_tlb_uop_T_2 & (will_fire_load_retry_0_will_fire ? casez_tmp_143 : will_fire_sta_retry_0_will_fire & casez_tmp_229) : will_fire_store_commit_0_will_fire ? casez_tmp_19 : will_fire_load_wakeup_0_will_fire & casez_tmp_313;
  assign io_dmem_req_bits_0_bits_uop_is_br = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_br : io_core_exe_0_req_bits_uop_is_br) : will_fire_load_retry_0_will_fire ? casez_tmp_144 : will_fire_sta_retry_0_will_fire & casez_tmp_230) : will_fire_store_commit_0_will_fire ? casez_tmp_20 : will_fire_load_wakeup_0_will_fire & casez_tmp_314;
  assign io_dmem_req_bits_0_bits_uop_is_jalr = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_jalr : io_core_exe_0_req_bits_uop_is_jalr) : will_fire_load_retry_0_will_fire ? casez_tmp_145 : will_fire_sta_retry_0_will_fire & casez_tmp_231) : will_fire_store_commit_0_will_fire ? casez_tmp_21 : will_fire_load_wakeup_0_will_fire & casez_tmp_315;
  assign io_dmem_req_bits_0_bits_uop_is_jal = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_jal : io_core_exe_0_req_bits_uop_is_jal) : will_fire_load_retry_0_will_fire ? casez_tmp_146 : will_fire_sta_retry_0_will_fire & casez_tmp_232) : will_fire_store_commit_0_will_fire ? casez_tmp_22 : will_fire_load_wakeup_0_will_fire & casez_tmp_316;
  assign io_dmem_req_bits_0_bits_uop_is_sfb = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_sfb : io_core_exe_0_req_bits_uop_is_sfb) : will_fire_load_retry_0_will_fire ? casez_tmp_147 : will_fire_sta_retry_0_will_fire & casez_tmp_233) : will_fire_store_commit_0_will_fire ? casez_tmp_23 : will_fire_load_wakeup_0_will_fire & casez_tmp_317;
  assign io_dmem_req_bits_0_bits_uop_br_mask = _GEN_275 ? exe_tlb_uop_0_br_mask : will_fire_store_commit_0_will_fire ? casez_tmp_24 : will_fire_load_wakeup_0_will_fire ? casez_tmp_318 : 20'h0;
  assign io_dmem_req_bits_0_bits_uop_br_tag = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_br_tag : io_core_exe_0_req_bits_uop_br_tag) : will_fire_load_retry_0_will_fire ? casez_tmp_149 : will_fire_sta_retry_0_will_fire ? casez_tmp_235 : 5'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_25 : will_fire_load_wakeup_0_will_fire ? casez_tmp_319 : 5'h0;
  assign io_dmem_req_bits_0_bits_uop_ftq_idx = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ftq_idx : io_core_exe_0_req_bits_uop_ftq_idx) : will_fire_load_retry_0_will_fire ? casez_tmp_150 : will_fire_sta_retry_0_will_fire ? casez_tmp_236 : 6'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_26 : will_fire_load_wakeup_0_will_fire ? casez_tmp_320 : 6'h0;
  assign io_dmem_req_bits_0_bits_uop_edge_inst = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_edge_inst : io_core_exe_0_req_bits_uop_edge_inst) : will_fire_load_retry_0_will_fire ? casez_tmp_151 : will_fire_sta_retry_0_will_fire & casez_tmp_237) : will_fire_store_commit_0_will_fire ? casez_tmp_27 : will_fire_load_wakeup_0_will_fire & casez_tmp_321;
  assign io_dmem_req_bits_0_bits_uop_pc_lob = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_pc_lob : io_core_exe_0_req_bits_uop_pc_lob) : will_fire_load_retry_0_will_fire ? casez_tmp_152 : will_fire_sta_retry_0_will_fire ? casez_tmp_238 : 6'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_28 : will_fire_load_wakeup_0_will_fire ? casez_tmp_322 : 6'h0;
  assign io_dmem_req_bits_0_bits_uop_taken = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_taken : io_core_exe_0_req_bits_uop_taken) : will_fire_load_retry_0_will_fire ? casez_tmp_153 : will_fire_sta_retry_0_will_fire & casez_tmp_239) : will_fire_store_commit_0_will_fire ? casez_tmp_29 : will_fire_load_wakeup_0_will_fire & casez_tmp_323;
  assign io_dmem_req_bits_0_bits_uop_imm_packed = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_imm_packed : io_core_exe_0_req_bits_uop_imm_packed) : will_fire_load_retry_0_will_fire ? casez_tmp_154 : will_fire_sta_retry_0_will_fire ? casez_tmp_240 : 20'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_30 : will_fire_load_wakeup_0_will_fire ? casez_tmp_324 : 20'h0;
  assign io_dmem_req_bits_0_bits_uop_csr_addr = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_csr_addr : io_core_exe_0_req_bits_uop_csr_addr) : will_fire_load_retry_0_will_fire ? casez_tmp_155 : will_fire_sta_retry_0_will_fire ? casez_tmp_241 : 12'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_31 : will_fire_load_wakeup_0_will_fire ? casez_tmp_325 : 12'h0;
  assign io_dmem_req_bits_0_bits_uop_rob_idx = _GEN_275 ? _mem_xcpt_uops_WIRE_0_rob_idx : will_fire_store_commit_0_will_fire ? casez_tmp_32 : will_fire_load_wakeup_0_will_fire ? casez_tmp_326 : 7'h0;
  assign io_dmem_req_bits_0_bits_uop_ldq_idx = _GEN_275 ? _mem_xcpt_uops_WIRE_0_ldq_idx : will_fire_store_commit_0_will_fire ? casez_tmp_33 : will_fire_load_wakeup_0_will_fire ? casez_tmp_327 : 5'h0;
  assign io_dmem_req_bits_0_bits_uop_stq_idx = _GEN_275 ? _mem_xcpt_uops_WIRE_0_stq_idx : will_fire_store_commit_0_will_fire ? casez_tmp_34 : will_fire_load_wakeup_0_will_fire ? casez_tmp_328 : 5'h0;
  assign io_dmem_req_bits_0_bits_uop_rxq_idx = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_rxq_idx : io_core_exe_0_req_bits_uop_rxq_idx) : will_fire_load_retry_0_will_fire ? casez_tmp_159 : will_fire_sta_retry_0_will_fire ? casez_tmp_245 : 2'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_35 : will_fire_load_wakeup_0_will_fire ? casez_tmp_329 : 2'h0;
  assign io_dmem_req_bits_0_bits_uop_pdst = _GEN_275 ? (_exe_tlb_uop_T_2 ? _mem_incoming_uop_WIRE_0_pdst : will_fire_load_retry_0_will_fire ? casez_tmp_160 : _exe_tlb_uop_T_4_pdst) : will_fire_store_commit_0_will_fire ? casez_tmp_36 : will_fire_load_wakeup_0_will_fire ? casez_tmp_330 : 7'h0;
  assign io_dmem_req_bits_0_bits_uop_prs1 = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_prs1 : io_core_exe_0_req_bits_uop_prs1) : will_fire_load_retry_0_will_fire ? casez_tmp_161 : will_fire_sta_retry_0_will_fire ? casez_tmp_247 : 7'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_37 : will_fire_load_wakeup_0_will_fire ? casez_tmp_331 : 7'h0;
  assign io_dmem_req_bits_0_bits_uop_prs2 = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_prs2 : io_core_exe_0_req_bits_uop_prs2) : will_fire_load_retry_0_will_fire ? casez_tmp_162 : will_fire_sta_retry_0_will_fire ? casez_tmp_248 : 7'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_38 : will_fire_load_wakeup_0_will_fire ? casez_tmp_332 : 7'h0;
  assign io_dmem_req_bits_0_bits_uop_prs3 = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_prs3 : io_core_exe_0_req_bits_uop_prs3) : will_fire_load_retry_0_will_fire ? casez_tmp_163 : will_fire_sta_retry_0_will_fire ? casez_tmp_249 : 7'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_39 : will_fire_load_wakeup_0_will_fire ? casez_tmp_333 : 7'h0;
  assign io_dmem_req_bits_0_bits_uop_ppred = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ppred : io_core_exe_0_req_bits_uop_ppred) : will_fire_load_retry_0_will_fire | ~will_fire_sta_retry_0_will_fire ? 6'h0 : casez_tmp_250) : will_fire_store_commit_0_will_fire ? casez_tmp_40 : 6'h0;
  assign io_dmem_req_bits_0_bits_uop_prs1_busy = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_prs1_busy : io_core_exe_0_req_bits_uop_prs1_busy) : will_fire_load_retry_0_will_fire ? casez_tmp_164 : will_fire_sta_retry_0_will_fire & casez_tmp_251) : will_fire_store_commit_0_will_fire ? casez_tmp_41 : will_fire_load_wakeup_0_will_fire & casez_tmp_334;
  assign io_dmem_req_bits_0_bits_uop_prs2_busy = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_prs2_busy : io_core_exe_0_req_bits_uop_prs2_busy) : will_fire_load_retry_0_will_fire ? casez_tmp_165 : will_fire_sta_retry_0_will_fire & casez_tmp_252) : will_fire_store_commit_0_will_fire ? casez_tmp_42 : will_fire_load_wakeup_0_will_fire & casez_tmp_335;
  assign io_dmem_req_bits_0_bits_uop_prs3_busy = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_prs3_busy : io_core_exe_0_req_bits_uop_prs3_busy) : will_fire_load_retry_0_will_fire ? casez_tmp_166 : will_fire_sta_retry_0_will_fire & casez_tmp_253) : will_fire_store_commit_0_will_fire ? casez_tmp_43 : will_fire_load_wakeup_0_will_fire & casez_tmp_336;
  assign io_dmem_req_bits_0_bits_uop_ppred_busy = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ppred_busy : io_core_exe_0_req_bits_uop_ppred_busy) : ~will_fire_load_retry_0_will_fire & will_fire_sta_retry_0_will_fire & casez_tmp_254) : will_fire_store_commit_0_will_fire & casez_tmp_44;
  assign io_dmem_req_bits_0_bits_uop_stale_pdst = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_stale_pdst : io_core_exe_0_req_bits_uop_stale_pdst) : will_fire_load_retry_0_will_fire ? casez_tmp_167 : will_fire_sta_retry_0_will_fire ? casez_tmp_255 : 7'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_45 : will_fire_load_wakeup_0_will_fire ? casez_tmp_337 : 7'h0;
  assign io_dmem_req_bits_0_bits_uop_exception = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_exception : io_core_exe_0_req_bits_uop_exception) : will_fire_load_retry_0_will_fire ? casez_tmp_168 : will_fire_sta_retry_0_will_fire & casez_tmp_256) : will_fire_store_commit_0_will_fire ? casez_tmp_46 : will_fire_load_wakeup_0_will_fire & casez_tmp_338;
  assign io_dmem_req_bits_0_bits_uop_exc_cause = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_exc_cause : io_core_exe_0_req_bits_uop_exc_cause) : will_fire_load_retry_0_will_fire ? casez_tmp_169 : will_fire_sta_retry_0_will_fire ? casez_tmp_257 : 64'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_47 : will_fire_load_wakeup_0_will_fire ? casez_tmp_339 : 64'h0;
  assign io_dmem_req_bits_0_bits_uop_bypassable = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_bypassable : io_core_exe_0_req_bits_uop_bypassable) : will_fire_load_retry_0_will_fire ? casez_tmp_170 : will_fire_sta_retry_0_will_fire & casez_tmp_258) : will_fire_store_commit_0_will_fire ? casez_tmp_48 : will_fire_load_wakeup_0_will_fire & casez_tmp_340;
  assign io_dmem_req_bits_0_bits_uop_mem_cmd = _GEN_275 ? exe_tlb_uop_0_mem_cmd : will_fire_store_commit_0_will_fire ? casez_tmp_49 : will_fire_load_wakeup_0_will_fire ? casez_tmp_341 : 5'h0;
  assign io_dmem_req_bits_0_bits_uop_mem_size = _GEN_275 ? exe_tlb_uop_0_mem_size : will_fire_store_commit_0_will_fire ? casez_tmp_50 : will_fire_load_wakeup_0_will_fire ? casez_tmp_342 : {2{will_fire_hella_incoming_0_will_fire | will_fire_hella_wakeup_0_will_fire}};
  assign io_dmem_req_bits_0_bits_uop_mem_signed = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_mem_signed : io_core_exe_0_req_bits_uop_mem_signed) : will_fire_load_retry_0_will_fire ? casez_tmp_173 : will_fire_sta_retry_0_will_fire & casez_tmp_261) : will_fire_store_commit_0_will_fire ? casez_tmp_51 : will_fire_load_wakeup_0_will_fire & casez_tmp_343;
  assign io_dmem_req_bits_0_bits_uop_is_fence = _GEN_275 ? exe_tlb_uop_0_is_fence : will_fire_store_commit_0_will_fire ? casez_tmp_52 : will_fire_load_wakeup_0_will_fire & casez_tmp_344;
  assign io_dmem_req_bits_0_bits_uop_is_fencei = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_fencei : io_core_exe_0_req_bits_uop_is_fencei) : will_fire_load_retry_0_will_fire ? casez_tmp_175 : will_fire_sta_retry_0_will_fire & casez_tmp_263) : will_fire_store_commit_0_will_fire ? casez_tmp_53 : will_fire_load_wakeup_0_will_fire & casez_tmp_345;
  assign io_dmem_req_bits_0_bits_uop_is_amo = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_amo : io_core_exe_0_req_bits_uop_is_amo) : will_fire_load_retry_0_will_fire ? casez_tmp_176 : will_fire_sta_retry_0_will_fire & casez_tmp_264) : will_fire_store_commit_0_will_fire ? casez_tmp_54 : will_fire_load_wakeup_0_will_fire & casez_tmp_346;
  assign io_dmem_req_bits_0_bits_uop_uses_ldq = _GEN_275 ? _mem_xcpt_uops_WIRE_0_uses_ldq : will_fire_store_commit_0_will_fire ? casez_tmp_55 : will_fire_load_wakeup_0_will_fire & casez_tmp_347;
  assign io_dmem_req_bits_0_bits_uop_uses_stq = _GEN_275 ? _mem_xcpt_uops_WIRE_0_uses_stq : will_fire_store_commit_0_will_fire ? casez_tmp_56 : will_fire_load_wakeup_0_will_fire & casez_tmp_348;
  assign io_dmem_req_bits_0_bits_uop_is_sys_pc2epc = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_sys_pc2epc : io_core_exe_0_req_bits_uop_is_sys_pc2epc) : will_fire_load_retry_0_will_fire ? casez_tmp_179 : will_fire_sta_retry_0_will_fire & casez_tmp_267) : will_fire_store_commit_0_will_fire ? casez_tmp_57 : will_fire_load_wakeup_0_will_fire & casez_tmp_349;
  assign io_dmem_req_bits_0_bits_uop_is_unique = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_unique : io_core_exe_0_req_bits_uop_is_unique) : will_fire_load_retry_0_will_fire ? casez_tmp_180 : will_fire_sta_retry_0_will_fire & casez_tmp_268) : will_fire_store_commit_0_will_fire ? casez_tmp_58 : will_fire_load_wakeup_0_will_fire & casez_tmp_350;
  assign io_dmem_req_bits_0_bits_uop_flush_on_commit = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_flush_on_commit : io_core_exe_0_req_bits_uop_flush_on_commit) : will_fire_load_retry_0_will_fire ? casez_tmp_181 : will_fire_sta_retry_0_will_fire & casez_tmp_269) : will_fire_store_commit_0_will_fire ? casez_tmp_59 : will_fire_load_wakeup_0_will_fire & casez_tmp_351;
  assign io_dmem_req_bits_0_bits_uop_ldst_is_rs1 = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ldst_is_rs1 : io_core_exe_0_req_bits_uop_ldst_is_rs1) : will_fire_load_retry_0_will_fire ? casez_tmp_182 : will_fire_sta_retry_0_will_fire & casez_tmp_270) : will_fire_store_commit_0_will_fire ? casez_tmp_60 : will_fire_load_wakeup_0_will_fire & casez_tmp_352;
  assign io_dmem_req_bits_0_bits_uop_ldst = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ldst : io_core_exe_0_req_bits_uop_ldst) : will_fire_load_retry_0_will_fire ? casez_tmp_183 : will_fire_sta_retry_0_will_fire ? casez_tmp_271 : 6'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_61 : will_fire_load_wakeup_0_will_fire ? casez_tmp_353 : 6'h0;
  assign io_dmem_req_bits_0_bits_uop_lrs1 = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_lrs1 : io_core_exe_0_req_bits_uop_lrs1) : will_fire_load_retry_0_will_fire ? casez_tmp_184 : will_fire_sta_retry_0_will_fire ? casez_tmp_272 : 6'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_62 : will_fire_load_wakeup_0_will_fire ? casez_tmp_354 : 6'h0;
  assign io_dmem_req_bits_0_bits_uop_lrs2 = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_lrs2 : io_core_exe_0_req_bits_uop_lrs2) : will_fire_load_retry_0_will_fire ? casez_tmp_185 : will_fire_sta_retry_0_will_fire ? casez_tmp_273 : 6'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_63 : will_fire_load_wakeup_0_will_fire ? casez_tmp_355 : 6'h0;
  assign io_dmem_req_bits_0_bits_uop_lrs3 = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_lrs3 : io_core_exe_0_req_bits_uop_lrs3) : will_fire_load_retry_0_will_fire ? casez_tmp_186 : will_fire_sta_retry_0_will_fire ? casez_tmp_274 : 6'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_64 : will_fire_load_wakeup_0_will_fire ? casez_tmp_356 : 6'h0;
  assign io_dmem_req_bits_0_bits_uop_ldst_val = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ldst_val : io_core_exe_0_req_bits_uop_ldst_val) : will_fire_load_retry_0_will_fire ? casez_tmp_187 : will_fire_sta_retry_0_will_fire & casez_tmp_275) : will_fire_store_commit_0_will_fire ? casez_tmp_65 : will_fire_load_wakeup_0_will_fire & casez_tmp_357;
  assign io_dmem_req_bits_0_bits_uop_dst_rtype = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_dst_rtype : io_core_exe_0_req_bits_uop_dst_rtype) : will_fire_load_retry_0_will_fire ? casez_tmp_188 : will_fire_sta_retry_0_will_fire ? casez_tmp_276 : 2'h2) : will_fire_store_commit_0_will_fire ? casez_tmp_66 : will_fire_load_wakeup_0_will_fire ? casez_tmp_358 : 2'h2;
  assign io_dmem_req_bits_0_bits_uop_lrs1_rtype = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_lrs1_rtype : io_core_exe_0_req_bits_uop_lrs1_rtype) : will_fire_load_retry_0_will_fire ? casez_tmp_189 : will_fire_sta_retry_0_will_fire ? casez_tmp_277 : 2'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_67 : will_fire_load_wakeup_0_will_fire ? casez_tmp_359 : 2'h0;
  assign io_dmem_req_bits_0_bits_uop_lrs2_rtype = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_lrs2_rtype : io_core_exe_0_req_bits_uop_lrs2_rtype) : will_fire_load_retry_0_will_fire ? casez_tmp_190 : will_fire_sta_retry_0_will_fire ? casez_tmp_278 : 2'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_68 : will_fire_load_wakeup_0_will_fire ? casez_tmp_360 : 2'h0;
  assign io_dmem_req_bits_0_bits_uop_frs3_en = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_frs3_en : io_core_exe_0_req_bits_uop_frs3_en) : will_fire_load_retry_0_will_fire ? casez_tmp_191 : will_fire_sta_retry_0_will_fire & casez_tmp_279) : will_fire_store_commit_0_will_fire ? casez_tmp_69 : will_fire_load_wakeup_0_will_fire & casez_tmp_361;
  assign io_dmem_req_bits_0_bits_uop_fp_val = _GEN_275 ? (_exe_tlb_uop_T_2 ? _mem_incoming_uop_WIRE_0_fp_val : will_fire_load_retry_0_will_fire ? casez_tmp_192 : will_fire_sta_retry_0_will_fire & casez_tmp_280) : will_fire_store_commit_0_will_fire ? casez_tmp_70 : will_fire_load_wakeup_0_will_fire & casez_tmp_362;
  assign io_dmem_req_bits_0_bits_uop_fp_single = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_fp_single : io_core_exe_0_req_bits_uop_fp_single) : will_fire_load_retry_0_will_fire ? casez_tmp_193 : will_fire_sta_retry_0_will_fire & casez_tmp_281) : will_fire_store_commit_0_will_fire ? casez_tmp_71 : will_fire_load_wakeup_0_will_fire & casez_tmp_363;
  assign io_dmem_req_bits_0_bits_uop_xcpt_pf_if = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_xcpt_pf_if : io_core_exe_0_req_bits_uop_xcpt_pf_if) : will_fire_load_retry_0_will_fire ? casez_tmp_194 : will_fire_sta_retry_0_will_fire & casez_tmp_282) : will_fire_store_commit_0_will_fire ? casez_tmp_72 : will_fire_load_wakeup_0_will_fire & casez_tmp_364;
  assign io_dmem_req_bits_0_bits_uop_xcpt_ae_if = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_xcpt_ae_if : io_core_exe_0_req_bits_uop_xcpt_ae_if) : will_fire_load_retry_0_will_fire ? casez_tmp_195 : will_fire_sta_retry_0_will_fire & casez_tmp_283) : will_fire_store_commit_0_will_fire ? casez_tmp_73 : will_fire_load_wakeup_0_will_fire & casez_tmp_365;
  assign io_dmem_req_bits_0_bits_uop_xcpt_ma_if = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_xcpt_ma_if : io_core_exe_0_req_bits_uop_xcpt_ma_if) : will_fire_load_retry_0_will_fire ? casez_tmp_196 : will_fire_sta_retry_0_will_fire & casez_tmp_284) : will_fire_store_commit_0_will_fire ? casez_tmp_74 : will_fire_load_wakeup_0_will_fire & casez_tmp_366;
  assign io_dmem_req_bits_0_bits_uop_bp_debug_if = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_bp_debug_if : io_core_exe_0_req_bits_uop_bp_debug_if) : will_fire_load_retry_0_will_fire ? casez_tmp_197 : will_fire_sta_retry_0_will_fire & casez_tmp_285) : will_fire_store_commit_0_will_fire ? casez_tmp_75 : will_fire_load_wakeup_0_will_fire & casez_tmp_367;
  assign io_dmem_req_bits_0_bits_uop_bp_xcpt_if = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_bp_xcpt_if : io_core_exe_0_req_bits_uop_bp_xcpt_if) : will_fire_load_retry_0_will_fire ? casez_tmp_198 : will_fire_sta_retry_0_will_fire & casez_tmp_286) : will_fire_store_commit_0_will_fire ? casez_tmp_76 : will_fire_load_wakeup_0_will_fire & casez_tmp_368;
  assign io_dmem_req_bits_0_bits_uop_debug_fsrc = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_debug_fsrc : io_core_exe_0_req_bits_uop_debug_fsrc) : will_fire_load_retry_0_will_fire ? casez_tmp_199 : will_fire_sta_retry_0_will_fire ? casez_tmp_287 : 2'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_77 : will_fire_load_wakeup_0_will_fire ? casez_tmp_369 : 2'h0;
  assign io_dmem_req_bits_0_bits_uop_debug_tsrc = _GEN_275 ? (_exe_tlb_uop_T_2 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_debug_tsrc : io_core_exe_0_req_bits_uop_debug_tsrc) : will_fire_load_retry_0_will_fire ? casez_tmp_200 : will_fire_sta_retry_0_will_fire ? casez_tmp_288 : 2'h0) : will_fire_store_commit_0_will_fire ? casez_tmp_78 : will_fire_load_wakeup_0_will_fire ? casez_tmp_370 : 2'h0;
  assign io_dmem_req_bits_0_bits_addr = _mem_paddr_WIRE_0;
  assign io_dmem_req_bits_0_bits_data = _GEN_275 ? 64'h0 : will_fire_store_commit_0_will_fire ? ((|casez_tmp_50) ? (casez_tmp_50 == 2'h1 ? {2{{2{casez_tmp_83[15:0]}}}} : casez_tmp_50 == 2'h2 ? {2{casez_tmp_83[31:0]}} : casez_tmp_83) : {2{{2{{2{casez_tmp_83[7:0]}}}}}}) : will_fire_load_wakeup_0_will_fire | will_fire_hella_incoming_0_will_fire | ~will_fire_hella_wakeup_0_will_fire ? 64'h0 : hella_data_data;
  assign io_dmem_req_bits_0_bits_is_hella = ~(_GEN_275 | will_fire_store_commit_0_will_fire | will_fire_load_wakeup_0_will_fire) & (will_fire_hella_incoming_0_will_fire | will_fire_hella_wakeup_0_will_fire);
  assign io_dmem_req_bits_1_valid = dmem_req_1_valid;
  assign io_dmem_req_bits_1_bits_uop_uopc = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_uopc : io_core_exe_0_req_bits_uop_uopc) : will_fire_load_retry_1_will_fire ? casez_tmp_124 : will_fire_sta_retry_1_will_fire ? casez_tmp_210 : 7'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_0 : will_fire_load_wakeup_1_will_fire ? casez_tmp_294 : 7'h0;
  assign io_dmem_req_bits_1_bits_uop_inst = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_inst : io_core_exe_0_req_bits_uop_inst) : will_fire_load_retry_1_will_fire ? casez_tmp_125 : will_fire_sta_retry_1_will_fire ? casez_tmp_211 : 32'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_1 : will_fire_load_wakeup_1_will_fire ? casez_tmp_295 : 32'h0;
  assign io_dmem_req_bits_1_bits_uop_debug_inst = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_debug_inst : io_core_exe_0_req_bits_uop_debug_inst) : will_fire_load_retry_1_will_fire ? casez_tmp_126 : will_fire_sta_retry_1_will_fire ? casez_tmp_212 : 32'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_2 : will_fire_load_wakeup_1_will_fire ? casez_tmp_296 : 32'h0;
  assign io_dmem_req_bits_1_bits_uop_is_rvc = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_rvc : io_core_exe_0_req_bits_uop_is_rvc) : will_fire_load_retry_1_will_fire ? casez_tmp_127 : will_fire_sta_retry_1_will_fire & casez_tmp_213) : will_fire_store_commit_1_will_fire ? casez_tmp_3 : will_fire_load_wakeup_1_will_fire & casez_tmp_297;
  assign io_dmem_req_bits_1_bits_uop_debug_pc = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_debug_pc : io_core_exe_0_req_bits_uop_debug_pc) : will_fire_load_retry_1_will_fire ? casez_tmp_128 : will_fire_sta_retry_1_will_fire ? casez_tmp_214 : 40'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_4 : will_fire_load_wakeup_1_will_fire ? casez_tmp_298 : 40'h0;
  assign io_dmem_req_bits_1_bits_uop_iq_type = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_iq_type : io_core_exe_0_req_bits_uop_iq_type) : will_fire_load_retry_1_will_fire ? casez_tmp_129 : will_fire_sta_retry_1_will_fire ? casez_tmp_215 : 3'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_5 : will_fire_load_wakeup_1_will_fire ? casez_tmp_299 : 3'h0;
  assign io_dmem_req_bits_1_bits_uop_fu_code = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_fu_code : io_core_exe_0_req_bits_uop_fu_code) : will_fire_load_retry_1_will_fire ? casez_tmp_130 : will_fire_sta_retry_1_will_fire ? casez_tmp_216 : 10'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_6 : will_fire_load_wakeup_1_will_fire ? casez_tmp_300 : 10'h0;
  assign io_dmem_req_bits_1_bits_uop_ctrl_br_type = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_br_type : io_core_exe_0_req_bits_uop_ctrl_br_type) : will_fire_load_retry_1_will_fire ? casez_tmp_131 : will_fire_sta_retry_1_will_fire ? casez_tmp_217 : 4'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_7 : will_fire_load_wakeup_1_will_fire ? casez_tmp_301 : 4'h0;
  assign io_dmem_req_bits_1_bits_uop_ctrl_op1_sel = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_op1_sel : io_core_exe_0_req_bits_uop_ctrl_op1_sel) : will_fire_load_retry_1_will_fire ? casez_tmp_132 : will_fire_sta_retry_1_will_fire ? casez_tmp_218 : 2'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_8 : will_fire_load_wakeup_1_will_fire ? casez_tmp_302 : 2'h0;
  assign io_dmem_req_bits_1_bits_uop_ctrl_op2_sel = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_op2_sel : io_core_exe_0_req_bits_uop_ctrl_op2_sel) : will_fire_load_retry_1_will_fire ? casez_tmp_133 : will_fire_sta_retry_1_will_fire ? casez_tmp_219 : 3'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_9 : will_fire_load_wakeup_1_will_fire ? casez_tmp_303 : 3'h0;
  assign io_dmem_req_bits_1_bits_uop_ctrl_imm_sel = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_imm_sel : io_core_exe_0_req_bits_uop_ctrl_imm_sel) : will_fire_load_retry_1_will_fire ? casez_tmp_134 : will_fire_sta_retry_1_will_fire ? casez_tmp_220 : 3'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_10 : will_fire_load_wakeup_1_will_fire ? casez_tmp_304 : 3'h0;
  assign io_dmem_req_bits_1_bits_uop_ctrl_op_fcn = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_op_fcn : io_core_exe_0_req_bits_uop_ctrl_op_fcn) : will_fire_load_retry_1_will_fire ? casez_tmp_135 : will_fire_sta_retry_1_will_fire ? casez_tmp_221 : 4'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_11 : will_fire_load_wakeup_1_will_fire ? casez_tmp_305 : 4'h0;
  assign io_dmem_req_bits_1_bits_uop_ctrl_fcn_dw = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_fcn_dw : io_core_exe_0_req_bits_uop_ctrl_fcn_dw) : will_fire_load_retry_1_will_fire ? casez_tmp_136 : will_fire_sta_retry_1_will_fire & casez_tmp_222) : will_fire_store_commit_1_will_fire ? casez_tmp_12 : will_fire_load_wakeup_1_will_fire & casez_tmp_306;
  assign io_dmem_req_bits_1_bits_uop_ctrl_csr_cmd = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ctrl_csr_cmd : io_core_exe_0_req_bits_uop_ctrl_csr_cmd) : will_fire_load_retry_1_will_fire ? casez_tmp_137 : will_fire_sta_retry_1_will_fire ? casez_tmp_223 : 3'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_13 : will_fire_load_wakeup_1_will_fire ? casez_tmp_307 : 3'h0;
  assign io_dmem_req_bits_1_bits_uop_ctrl_is_load = _GEN_281 ? exe_tlb_uop_1_ctrl_is_load : will_fire_store_commit_1_will_fire ? casez_tmp_14 : will_fire_load_wakeup_1_will_fire & casez_tmp_308;
  assign io_dmem_req_bits_1_bits_uop_ctrl_is_sta = _GEN_281 ? exe_tlb_uop_1_ctrl_is_sta : will_fire_store_commit_1_will_fire ? casez_tmp_15 : will_fire_load_wakeup_1_will_fire & casez_tmp_309;
  assign io_dmem_req_bits_1_bits_uop_ctrl_is_std = _GEN_281 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_ctrl_is_std : will_fire_load_retry_1_will_fire ? casez_tmp_140 : will_fire_sta_retry_1_will_fire & casez_tmp_226) : will_fire_store_commit_1_will_fire ? casez_tmp_16 : will_fire_load_wakeup_1_will_fire & casez_tmp_310;
  assign io_dmem_req_bits_1_bits_uop_iw_state = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_iw_state : io_core_exe_0_req_bits_uop_iw_state) : will_fire_load_retry_1_will_fire ? casez_tmp_141 : will_fire_sta_retry_1_will_fire ? casez_tmp_227 : 2'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_17 : will_fire_load_wakeup_1_will_fire ? casez_tmp_311 : 2'h0;
  assign io_dmem_req_bits_1_bits_uop_iw_p1_poisoned = _GEN_281 ? ~_exe_tlb_uop_T_9 & (will_fire_load_retry_1_will_fire ? casez_tmp_142 : will_fire_sta_retry_1_will_fire & casez_tmp_228) : will_fire_store_commit_1_will_fire ? casez_tmp_18 : will_fire_load_wakeup_1_will_fire & casez_tmp_312;
  assign io_dmem_req_bits_1_bits_uop_iw_p2_poisoned = _GEN_281 ? ~_exe_tlb_uop_T_9 & (will_fire_load_retry_1_will_fire ? casez_tmp_143 : will_fire_sta_retry_1_will_fire & casez_tmp_229) : will_fire_store_commit_1_will_fire ? casez_tmp_19 : will_fire_load_wakeup_1_will_fire & casez_tmp_313;
  assign io_dmem_req_bits_1_bits_uop_is_br = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_br : io_core_exe_0_req_bits_uop_is_br) : will_fire_load_retry_1_will_fire ? casez_tmp_144 : will_fire_sta_retry_1_will_fire & casez_tmp_230) : will_fire_store_commit_1_will_fire ? casez_tmp_20 : will_fire_load_wakeup_1_will_fire & casez_tmp_314;
  assign io_dmem_req_bits_1_bits_uop_is_jalr = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_jalr : io_core_exe_0_req_bits_uop_is_jalr) : will_fire_load_retry_1_will_fire ? casez_tmp_145 : will_fire_sta_retry_1_will_fire & casez_tmp_231) : will_fire_store_commit_1_will_fire ? casez_tmp_21 : will_fire_load_wakeup_1_will_fire & casez_tmp_315;
  assign io_dmem_req_bits_1_bits_uop_is_jal = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_jal : io_core_exe_0_req_bits_uop_is_jal) : will_fire_load_retry_1_will_fire ? casez_tmp_146 : will_fire_sta_retry_1_will_fire & casez_tmp_232) : will_fire_store_commit_1_will_fire ? casez_tmp_22 : will_fire_load_wakeup_1_will_fire & casez_tmp_316;
  assign io_dmem_req_bits_1_bits_uop_is_sfb = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_sfb : io_core_exe_0_req_bits_uop_is_sfb) : will_fire_load_retry_1_will_fire ? casez_tmp_147 : will_fire_sta_retry_1_will_fire & casez_tmp_233) : will_fire_store_commit_1_will_fire ? casez_tmp_23 : will_fire_load_wakeup_1_will_fire & casez_tmp_317;
  assign io_dmem_req_bits_1_bits_uop_br_mask = _GEN_281 ? exe_tlb_uop_1_br_mask : will_fire_store_commit_1_will_fire ? casez_tmp_24 : will_fire_load_wakeup_1_will_fire ? casez_tmp_318 : 20'h0;
  assign io_dmem_req_bits_1_bits_uop_br_tag = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_br_tag : io_core_exe_0_req_bits_uop_br_tag) : will_fire_load_retry_1_will_fire ? casez_tmp_149 : will_fire_sta_retry_1_will_fire ? casez_tmp_235 : 5'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_25 : will_fire_load_wakeup_1_will_fire ? casez_tmp_319 : 5'h0;
  assign io_dmem_req_bits_1_bits_uop_ftq_idx = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ftq_idx : io_core_exe_0_req_bits_uop_ftq_idx) : will_fire_load_retry_1_will_fire ? casez_tmp_150 : will_fire_sta_retry_1_will_fire ? casez_tmp_236 : 6'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_26 : will_fire_load_wakeup_1_will_fire ? casez_tmp_320 : 6'h0;
  assign io_dmem_req_bits_1_bits_uop_edge_inst = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_edge_inst : io_core_exe_0_req_bits_uop_edge_inst) : will_fire_load_retry_1_will_fire ? casez_tmp_151 : will_fire_sta_retry_1_will_fire & casez_tmp_237) : will_fire_store_commit_1_will_fire ? casez_tmp_27 : will_fire_load_wakeup_1_will_fire & casez_tmp_321;
  assign io_dmem_req_bits_1_bits_uop_pc_lob = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_pc_lob : io_core_exe_0_req_bits_uop_pc_lob) : will_fire_load_retry_1_will_fire ? casez_tmp_152 : will_fire_sta_retry_1_will_fire ? casez_tmp_238 : 6'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_28 : will_fire_load_wakeup_1_will_fire ? casez_tmp_322 : 6'h0;
  assign io_dmem_req_bits_1_bits_uop_taken = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_taken : io_core_exe_0_req_bits_uop_taken) : will_fire_load_retry_1_will_fire ? casez_tmp_153 : will_fire_sta_retry_1_will_fire & casez_tmp_239) : will_fire_store_commit_1_will_fire ? casez_tmp_29 : will_fire_load_wakeup_1_will_fire & casez_tmp_323;
  assign io_dmem_req_bits_1_bits_uop_imm_packed = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_imm_packed : io_core_exe_0_req_bits_uop_imm_packed) : will_fire_load_retry_1_will_fire ? casez_tmp_154 : will_fire_sta_retry_1_will_fire ? casez_tmp_240 : 20'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_30 : will_fire_load_wakeup_1_will_fire ? casez_tmp_324 : 20'h0;
  assign io_dmem_req_bits_1_bits_uop_csr_addr = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_csr_addr : io_core_exe_0_req_bits_uop_csr_addr) : will_fire_load_retry_1_will_fire ? casez_tmp_155 : will_fire_sta_retry_1_will_fire ? casez_tmp_241 : 12'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_31 : will_fire_load_wakeup_1_will_fire ? casez_tmp_325 : 12'h0;
  assign io_dmem_req_bits_1_bits_uop_rob_idx = _GEN_281 ? _mem_xcpt_uops_WIRE_1_rob_idx : will_fire_store_commit_1_will_fire ? casez_tmp_32 : will_fire_load_wakeup_1_will_fire ? casez_tmp_326 : 7'h0;
  assign io_dmem_req_bits_1_bits_uop_ldq_idx = _GEN_281 ? _mem_xcpt_uops_WIRE_1_ldq_idx : will_fire_store_commit_1_will_fire ? casez_tmp_33 : will_fire_load_wakeup_1_will_fire ? casez_tmp_327 : 5'h0;
  assign io_dmem_req_bits_1_bits_uop_stq_idx = _GEN_281 ? _mem_xcpt_uops_WIRE_1_stq_idx : will_fire_store_commit_1_will_fire ? casez_tmp_34 : will_fire_load_wakeup_1_will_fire ? casez_tmp_328 : 5'h0;
  assign io_dmem_req_bits_1_bits_uop_rxq_idx = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_rxq_idx : io_core_exe_0_req_bits_uop_rxq_idx) : will_fire_load_retry_1_will_fire ? casez_tmp_159 : will_fire_sta_retry_1_will_fire ? casez_tmp_245 : 2'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_35 : will_fire_load_wakeup_1_will_fire ? casez_tmp_329 : 2'h0;
  assign io_dmem_req_bits_1_bits_uop_pdst = _GEN_281 ? (_exe_tlb_uop_T_9 ? _mem_incoming_uop_WIRE_1_pdst : will_fire_load_retry_1_will_fire ? casez_tmp_160 : _exe_tlb_uop_T_11_pdst) : will_fire_store_commit_1_will_fire ? casez_tmp_36 : will_fire_load_wakeup_1_will_fire ? casez_tmp_330 : 7'h0;
  assign io_dmem_req_bits_1_bits_uop_prs1 = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_prs1 : io_core_exe_0_req_bits_uop_prs1) : will_fire_load_retry_1_will_fire ? casez_tmp_161 : will_fire_sta_retry_1_will_fire ? casez_tmp_247 : 7'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_37 : will_fire_load_wakeup_1_will_fire ? casez_tmp_331 : 7'h0;
  assign io_dmem_req_bits_1_bits_uop_prs2 = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_prs2 : io_core_exe_0_req_bits_uop_prs2) : will_fire_load_retry_1_will_fire ? casez_tmp_162 : will_fire_sta_retry_1_will_fire ? casez_tmp_248 : 7'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_38 : will_fire_load_wakeup_1_will_fire ? casez_tmp_332 : 7'h0;
  assign io_dmem_req_bits_1_bits_uop_prs3 = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_prs3 : io_core_exe_0_req_bits_uop_prs3) : will_fire_load_retry_1_will_fire ? casez_tmp_163 : will_fire_sta_retry_1_will_fire ? casez_tmp_249 : 7'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_39 : will_fire_load_wakeup_1_will_fire ? casez_tmp_333 : 7'h0;
  assign io_dmem_req_bits_1_bits_uop_ppred = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ppred : io_core_exe_0_req_bits_uop_ppred) : will_fire_load_retry_1_will_fire | ~will_fire_sta_retry_1_will_fire ? 6'h0 : casez_tmp_250) : will_fire_store_commit_1_will_fire ? casez_tmp_40 : 6'h0;
  assign io_dmem_req_bits_1_bits_uop_prs1_busy = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_prs1_busy : io_core_exe_0_req_bits_uop_prs1_busy) : will_fire_load_retry_1_will_fire ? casez_tmp_164 : will_fire_sta_retry_1_will_fire & casez_tmp_251) : will_fire_store_commit_1_will_fire ? casez_tmp_41 : will_fire_load_wakeup_1_will_fire & casez_tmp_334;
  assign io_dmem_req_bits_1_bits_uop_prs2_busy = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_prs2_busy : io_core_exe_0_req_bits_uop_prs2_busy) : will_fire_load_retry_1_will_fire ? casez_tmp_165 : will_fire_sta_retry_1_will_fire & casez_tmp_252) : will_fire_store_commit_1_will_fire ? casez_tmp_42 : will_fire_load_wakeup_1_will_fire & casez_tmp_335;
  assign io_dmem_req_bits_1_bits_uop_prs3_busy = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_prs3_busy : io_core_exe_0_req_bits_uop_prs3_busy) : will_fire_load_retry_1_will_fire ? casez_tmp_166 : will_fire_sta_retry_1_will_fire & casez_tmp_253) : will_fire_store_commit_1_will_fire ? casez_tmp_43 : will_fire_load_wakeup_1_will_fire & casez_tmp_336;
  assign io_dmem_req_bits_1_bits_uop_ppred_busy = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ppred_busy : io_core_exe_0_req_bits_uop_ppred_busy) : ~will_fire_load_retry_1_will_fire & will_fire_sta_retry_1_will_fire & casez_tmp_254) : will_fire_store_commit_1_will_fire & casez_tmp_44;
  assign io_dmem_req_bits_1_bits_uop_stale_pdst = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_stale_pdst : io_core_exe_0_req_bits_uop_stale_pdst) : will_fire_load_retry_1_will_fire ? casez_tmp_167 : will_fire_sta_retry_1_will_fire ? casez_tmp_255 : 7'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_45 : will_fire_load_wakeup_1_will_fire ? casez_tmp_337 : 7'h0;
  assign io_dmem_req_bits_1_bits_uop_exception = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_exception : io_core_exe_0_req_bits_uop_exception) : will_fire_load_retry_1_will_fire ? casez_tmp_168 : will_fire_sta_retry_1_will_fire & casez_tmp_256) : will_fire_store_commit_1_will_fire ? casez_tmp_46 : will_fire_load_wakeup_1_will_fire & casez_tmp_338;
  assign io_dmem_req_bits_1_bits_uop_exc_cause = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_exc_cause : io_core_exe_0_req_bits_uop_exc_cause) : will_fire_load_retry_1_will_fire ? casez_tmp_169 : will_fire_sta_retry_1_will_fire ? casez_tmp_257 : 64'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_47 : will_fire_load_wakeup_1_will_fire ? casez_tmp_339 : 64'h0;
  assign io_dmem_req_bits_1_bits_uop_bypassable = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_bypassable : io_core_exe_0_req_bits_uop_bypassable) : will_fire_load_retry_1_will_fire ? casez_tmp_170 : will_fire_sta_retry_1_will_fire & casez_tmp_258) : will_fire_store_commit_1_will_fire ? casez_tmp_48 : will_fire_load_wakeup_1_will_fire & casez_tmp_340;
  assign io_dmem_req_bits_1_bits_uop_mem_cmd = _GEN_281 ? exe_tlb_uop_1_mem_cmd : will_fire_store_commit_1_will_fire ? casez_tmp_49 : will_fire_load_wakeup_1_will_fire ? casez_tmp_341 : 5'h0;
  assign io_dmem_req_bits_1_bits_uop_mem_size = _GEN_281 ? exe_tlb_uop_1_mem_size : will_fire_store_commit_1_will_fire ? casez_tmp_50 : will_fire_load_wakeup_1_will_fire ? casez_tmp_342 : {2{will_fire_hella_incoming_1_will_fire | will_fire_hella_wakeup_1_will_fire}};
  assign io_dmem_req_bits_1_bits_uop_mem_signed = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_mem_signed : io_core_exe_0_req_bits_uop_mem_signed) : will_fire_load_retry_1_will_fire ? casez_tmp_173 : will_fire_sta_retry_1_will_fire & casez_tmp_261) : will_fire_store_commit_1_will_fire ? casez_tmp_51 : will_fire_load_wakeup_1_will_fire & casez_tmp_343;
  assign io_dmem_req_bits_1_bits_uop_is_fence = _GEN_281 ? exe_tlb_uop_1_is_fence : will_fire_store_commit_1_will_fire ? casez_tmp_52 : will_fire_load_wakeup_1_will_fire & casez_tmp_344;
  assign io_dmem_req_bits_1_bits_uop_is_fencei = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_fencei : io_core_exe_0_req_bits_uop_is_fencei) : will_fire_load_retry_1_will_fire ? casez_tmp_175 : will_fire_sta_retry_1_will_fire & casez_tmp_263) : will_fire_store_commit_1_will_fire ? casez_tmp_53 : will_fire_load_wakeup_1_will_fire & casez_tmp_345;
  assign io_dmem_req_bits_1_bits_uop_is_amo = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_amo : io_core_exe_0_req_bits_uop_is_amo) : will_fire_load_retry_1_will_fire ? casez_tmp_176 : will_fire_sta_retry_1_will_fire & casez_tmp_264) : will_fire_store_commit_1_will_fire ? casez_tmp_54 : will_fire_load_wakeup_1_will_fire & casez_tmp_346;
  assign io_dmem_req_bits_1_bits_uop_uses_ldq = _GEN_281 ? _mem_xcpt_uops_WIRE_1_uses_ldq : will_fire_store_commit_1_will_fire ? casez_tmp_55 : will_fire_load_wakeup_1_will_fire & casez_tmp_347;
  assign io_dmem_req_bits_1_bits_uop_uses_stq = _GEN_281 ? _mem_xcpt_uops_WIRE_1_uses_stq : will_fire_store_commit_1_will_fire ? casez_tmp_56 : will_fire_load_wakeup_1_will_fire & casez_tmp_348;
  assign io_dmem_req_bits_1_bits_uop_is_sys_pc2epc = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_sys_pc2epc : io_core_exe_0_req_bits_uop_is_sys_pc2epc) : will_fire_load_retry_1_will_fire ? casez_tmp_179 : will_fire_sta_retry_1_will_fire & casez_tmp_267) : will_fire_store_commit_1_will_fire ? casez_tmp_57 : will_fire_load_wakeup_1_will_fire & casez_tmp_349;
  assign io_dmem_req_bits_1_bits_uop_is_unique = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_is_unique : io_core_exe_0_req_bits_uop_is_unique) : will_fire_load_retry_1_will_fire ? casez_tmp_180 : will_fire_sta_retry_1_will_fire & casez_tmp_268) : will_fire_store_commit_1_will_fire ? casez_tmp_58 : will_fire_load_wakeup_1_will_fire & casez_tmp_350;
  assign io_dmem_req_bits_1_bits_uop_flush_on_commit = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_flush_on_commit : io_core_exe_0_req_bits_uop_flush_on_commit) : will_fire_load_retry_1_will_fire ? casez_tmp_181 : will_fire_sta_retry_1_will_fire & casez_tmp_269) : will_fire_store_commit_1_will_fire ? casez_tmp_59 : will_fire_load_wakeup_1_will_fire & casez_tmp_351;
  assign io_dmem_req_bits_1_bits_uop_ldst_is_rs1 = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ldst_is_rs1 : io_core_exe_0_req_bits_uop_ldst_is_rs1) : will_fire_load_retry_1_will_fire ? casez_tmp_182 : will_fire_sta_retry_1_will_fire & casez_tmp_270) : will_fire_store_commit_1_will_fire ? casez_tmp_60 : will_fire_load_wakeup_1_will_fire & casez_tmp_352;
  assign io_dmem_req_bits_1_bits_uop_ldst = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ldst : io_core_exe_0_req_bits_uop_ldst) : will_fire_load_retry_1_will_fire ? casez_tmp_183 : will_fire_sta_retry_1_will_fire ? casez_tmp_271 : 6'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_61 : will_fire_load_wakeup_1_will_fire ? casez_tmp_353 : 6'h0;
  assign io_dmem_req_bits_1_bits_uop_lrs1 = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_lrs1 : io_core_exe_0_req_bits_uop_lrs1) : will_fire_load_retry_1_will_fire ? casez_tmp_184 : will_fire_sta_retry_1_will_fire ? casez_tmp_272 : 6'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_62 : will_fire_load_wakeup_1_will_fire ? casez_tmp_354 : 6'h0;
  assign io_dmem_req_bits_1_bits_uop_lrs2 = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_lrs2 : io_core_exe_0_req_bits_uop_lrs2) : will_fire_load_retry_1_will_fire ? casez_tmp_185 : will_fire_sta_retry_1_will_fire ? casez_tmp_273 : 6'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_63 : will_fire_load_wakeup_1_will_fire ? casez_tmp_355 : 6'h0;
  assign io_dmem_req_bits_1_bits_uop_lrs3 = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_lrs3 : io_core_exe_0_req_bits_uop_lrs3) : will_fire_load_retry_1_will_fire ? casez_tmp_186 : will_fire_sta_retry_1_will_fire ? casez_tmp_274 : 6'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_64 : will_fire_load_wakeup_1_will_fire ? casez_tmp_356 : 6'h0;
  assign io_dmem_req_bits_1_bits_uop_ldst_val = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_ldst_val : io_core_exe_0_req_bits_uop_ldst_val) : will_fire_load_retry_1_will_fire ? casez_tmp_187 : will_fire_sta_retry_1_will_fire & casez_tmp_275) : will_fire_store_commit_1_will_fire ? casez_tmp_65 : will_fire_load_wakeup_1_will_fire & casez_tmp_357;
  assign io_dmem_req_bits_1_bits_uop_dst_rtype = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_dst_rtype : io_core_exe_0_req_bits_uop_dst_rtype) : will_fire_load_retry_1_will_fire ? casez_tmp_188 : will_fire_sta_retry_1_will_fire ? casez_tmp_276 : 2'h2) : will_fire_store_commit_1_will_fire ? casez_tmp_66 : will_fire_load_wakeup_1_will_fire ? casez_tmp_358 : 2'h2;
  assign io_dmem_req_bits_1_bits_uop_lrs1_rtype = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_lrs1_rtype : io_core_exe_0_req_bits_uop_lrs1_rtype) : will_fire_load_retry_1_will_fire ? casez_tmp_189 : will_fire_sta_retry_1_will_fire ? casez_tmp_277 : 2'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_67 : will_fire_load_wakeup_1_will_fire ? casez_tmp_359 : 2'h0;
  assign io_dmem_req_bits_1_bits_uop_lrs2_rtype = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_lrs2_rtype : io_core_exe_0_req_bits_uop_lrs2_rtype) : will_fire_load_retry_1_will_fire ? casez_tmp_190 : will_fire_sta_retry_1_will_fire ? casez_tmp_278 : 2'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_68 : will_fire_load_wakeup_1_will_fire ? casez_tmp_360 : 2'h0;
  assign io_dmem_req_bits_1_bits_uop_frs3_en = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_frs3_en : io_core_exe_0_req_bits_uop_frs3_en) : will_fire_load_retry_1_will_fire ? casez_tmp_191 : will_fire_sta_retry_1_will_fire & casez_tmp_279) : will_fire_store_commit_1_will_fire ? casez_tmp_69 : will_fire_load_wakeup_1_will_fire & casez_tmp_361;
  assign io_dmem_req_bits_1_bits_uop_fp_val = _GEN_281 ? (_exe_tlb_uop_T_9 ? _mem_incoming_uop_WIRE_1_fp_val : will_fire_load_retry_1_will_fire ? casez_tmp_192 : will_fire_sta_retry_1_will_fire & casez_tmp_280) : will_fire_store_commit_1_will_fire ? casez_tmp_70 : will_fire_load_wakeup_1_will_fire & casez_tmp_362;
  assign io_dmem_req_bits_1_bits_uop_fp_single = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_fp_single : io_core_exe_0_req_bits_uop_fp_single) : will_fire_load_retry_1_will_fire ? casez_tmp_193 : will_fire_sta_retry_1_will_fire & casez_tmp_281) : will_fire_store_commit_1_will_fire ? casez_tmp_71 : will_fire_load_wakeup_1_will_fire & casez_tmp_363;
  assign io_dmem_req_bits_1_bits_uop_xcpt_pf_if = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_xcpt_pf_if : io_core_exe_0_req_bits_uop_xcpt_pf_if) : will_fire_load_retry_1_will_fire ? casez_tmp_194 : will_fire_sta_retry_1_will_fire & casez_tmp_282) : will_fire_store_commit_1_will_fire ? casez_tmp_72 : will_fire_load_wakeup_1_will_fire & casez_tmp_364;
  assign io_dmem_req_bits_1_bits_uop_xcpt_ae_if = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_xcpt_ae_if : io_core_exe_0_req_bits_uop_xcpt_ae_if) : will_fire_load_retry_1_will_fire ? casez_tmp_195 : will_fire_sta_retry_1_will_fire & casez_tmp_283) : will_fire_store_commit_1_will_fire ? casez_tmp_73 : will_fire_load_wakeup_1_will_fire & casez_tmp_365;
  assign io_dmem_req_bits_1_bits_uop_xcpt_ma_if = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_xcpt_ma_if : io_core_exe_0_req_bits_uop_xcpt_ma_if) : will_fire_load_retry_1_will_fire ? casez_tmp_196 : will_fire_sta_retry_1_will_fire & casez_tmp_284) : will_fire_store_commit_1_will_fire ? casez_tmp_74 : will_fire_load_wakeup_1_will_fire & casez_tmp_366;
  assign io_dmem_req_bits_1_bits_uop_bp_debug_if = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_bp_debug_if : io_core_exe_0_req_bits_uop_bp_debug_if) : will_fire_load_retry_1_will_fire ? casez_tmp_197 : will_fire_sta_retry_1_will_fire & casez_tmp_285) : will_fire_store_commit_1_will_fire ? casez_tmp_75 : will_fire_load_wakeup_1_will_fire & casez_tmp_367;
  assign io_dmem_req_bits_1_bits_uop_bp_xcpt_if = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_bp_xcpt_if : io_core_exe_0_req_bits_uop_bp_xcpt_if) : will_fire_load_retry_1_will_fire ? casez_tmp_198 : will_fire_sta_retry_1_will_fire & casez_tmp_286) : will_fire_store_commit_1_will_fire ? casez_tmp_76 : will_fire_load_wakeup_1_will_fire & casez_tmp_368;
  assign io_dmem_req_bits_1_bits_uop_debug_fsrc = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_debug_fsrc : io_core_exe_0_req_bits_uop_debug_fsrc) : will_fire_load_retry_1_will_fire ? casez_tmp_199 : will_fire_sta_retry_1_will_fire ? casez_tmp_287 : 2'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_77 : will_fire_load_wakeup_1_will_fire ? casez_tmp_369 : 2'h0;
  assign io_dmem_req_bits_1_bits_uop_debug_tsrc = _GEN_281 ? (_exe_tlb_uop_T_9 ? (_GEN_17 ? io_core_exe_1_req_bits_uop_debug_tsrc : io_core_exe_0_req_bits_uop_debug_tsrc) : will_fire_load_retry_1_will_fire ? casez_tmp_200 : will_fire_sta_retry_1_will_fire ? casez_tmp_288 : 2'h0) : will_fire_store_commit_1_will_fire ? casez_tmp_78 : will_fire_load_wakeup_1_will_fire ? casez_tmp_370 : 2'h0;
  assign io_dmem_req_bits_1_bits_addr = _mem_paddr_WIRE_1;
  assign io_dmem_req_bits_1_bits_data = _GEN_281 ? 64'h0 : will_fire_store_commit_1_will_fire ? ((|casez_tmp_50) ? (casez_tmp_50 == 2'h1 ? {2{{2{casez_tmp_83[15:0]}}}} : casez_tmp_50 == 2'h2 ? {2{casez_tmp_83[31:0]}} : casez_tmp_83) : {2{{2{{2{casez_tmp_83[7:0]}}}}}}) : will_fire_load_wakeup_1_will_fire | will_fire_hella_incoming_1_will_fire | ~will_fire_hella_wakeup_1_will_fire ? 64'h0 : hella_data_data;
  assign io_dmem_req_bits_1_bits_is_hella = ~(_GEN_281 | will_fire_store_commit_1_will_fire | will_fire_load_wakeup_1_will_fire) & (will_fire_hella_incoming_1_will_fire | will_fire_hella_wakeup_1_will_fire);
  assign io_dmem_s1_kill_0 = _GEN_1421 ? (_GEN_1423 ? io_dmem_s1_kill_0_REG_125 : _GEN_1424 ? io_dmem_s1_kill_0_REG_126 : _GEN_1425 ? io_dmem_s1_kill_0_REG_127 : _GEN_1415) : _GEN_1415;
  assign io_dmem_s1_kill_1 = _GEN_1426 ? (_GEN_1428 ? io_dmem_s1_kill_1_REG_125 : _GEN_1429 ? io_dmem_s1_kill_1_REG_126 : _GEN_1425 ? io_dmem_s1_kill_1_REG_127 : _GEN_1420) : _GEN_1420;
  assign io_dmem_brupdate_b1_resolve_mask = io_core_brupdate_b1_resolve_mask;
  assign io_dmem_brupdate_b1_mispredict_mask = io_core_brupdate_b1_mispredict_mask;
  assign io_dmem_exception = io_core_exception;
  assign io_dmem_release_ready = will_fire_release_0_will_fire | will_fire_release_1_will_fire;
  assign io_dmem_force_order = _GEN_1577 & _GEN_1578 | io_core_fence_dmem;
  assign io_hellacache_req_ready = _io_hellacache_req_ready_output;
  assign io_hellacache_s2_nack = ~_GEN_1581 & _GEN_1580;
  assign io_hellacache_resp_valid = ~(_GEN_1581 | _GEN_1580 | _GEN_1582) & _GEN_1431 & (_GEN_1584 | _GEN_1583);
  assign io_hellacache_resp_bits_data = _GEN_1584 ? io_dmem_resp_1_bits_data : io_dmem_resp_0_bits_data;
  assign io_hellacache_s2_xcpt_ae_ld = ~(_io_hellacache_req_ready_output | _GEN_2 | _GEN_1580) & _GEN_1582 & hella_xcpt_ae_ld;
endmodule

