// Standard header to adapt well known macros for prints and assertions.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module Queue_24(
  input        clock,
               reset,
  output       io_enq_ready,
  input        io_enq_valid,
               io_enq_bits_noop,
  input  [2:0] io_enq_bits_way,
  input  [9:0] io_enq_bits_set,
  input  [2:0] io_enq_bits_beat,
  input        io_deq_ready,
  output       io_deq_valid,
               io_deq_bits_noop,
  output [2:0] io_deq_bits_way,
  output [9:0] io_deq_bits_set,
  output [2:0] io_deq_bits_beat,
  output       io_deq_bits_mask
);

  reg  [17:0] ram;
  reg         full;
  wire        _io_enq_ready_output = io_deq_ready | ~full;
  wire        do_enq = _io_enq_ready_output & io_enq_valid;
  always @(posedge clock) begin
    if (do_enq)
      ram <= {1'h1, io_enq_bits_beat, io_enq_bits_set, io_enq_bits_way, io_enq_bits_noop};
    if (reset)
      full <= 1'h0;
    else if (~(do_enq == (io_deq_ready & full)))
      full <= do_enq;
  end // always @(posedge)
  assign io_enq_ready = _io_enq_ready_output;
  assign io_deq_valid = full;
  assign io_deq_bits_noop = ram[0];
  assign io_deq_bits_way = ram[3:1];
  assign io_deq_bits_set = ram[13:4];
  assign io_deq_bits_beat = ram[16:14];
  assign io_deq_bits_mask = ram[17];
endmodule

